module testbench_specparam_declaration;
    specparam_declaration0 specparam_declaration_instance0();
    specparam_declaration1 specparam_declaration_instance1();
    specparam_declaration2 specparam_declaration_instance2();
    specparam_declaration3 specparam_declaration_instance3();
    specparam_declaration4 specparam_declaration_instance4();
    specparam_declaration5 specparam_declaration_instance5();
    specparam_declaration6 specparam_declaration_instance6();
    specparam_declaration7 specparam_declaration_instance7();
    specparam_declaration8 specparam_declaration_instance8();
    specparam_declaration9 specparam_declaration_instance9();
    specparam_declaration10 specparam_declaration_instance10();
    specparam_declaration11 specparam_declaration_instance11();
    specparam_declaration12 specparam_declaration_instance12();
    specparam_declaration13 specparam_declaration_instance13();
    specparam_declaration14 specparam_declaration_instance14();
    specparam_declaration15 specparam_declaration_instance15();
    specparam_declaration16 specparam_declaration_instance16();
    specparam_declaration17 specparam_declaration_instance17();
    specparam_declaration18 specparam_declaration_instance18();
    specparam_declaration19 specparam_declaration_instance19();
    specparam_declaration20 specparam_declaration_instance20();
    specparam_declaration21 specparam_declaration_instance21();
    specparam_declaration22 specparam_declaration_instance22();
    specparam_declaration23 specparam_declaration_instance23();
    specparam_declaration24 specparam_declaration_instance24();
    specparam_declaration25 specparam_declaration_instance25();
    specparam_declaration26 specparam_declaration_instance26();
    specparam_declaration27 specparam_declaration_instance27();
    specparam_declaration28 specparam_declaration_instance28();
    specparam_declaration29 specparam_declaration_instance29();
    specparam_declaration30 specparam_declaration_instance30();
    specparam_declaration31 specparam_declaration_instance31();
    specparam_declaration32 specparam_declaration_instance32();
    specparam_declaration33 specparam_declaration_instance33();
    specparam_declaration34 specparam_declaration_instance34();
    specparam_declaration35 specparam_declaration_instance35();
    specparam_declaration36 specparam_declaration_instance36();
    specparam_declaration37 specparam_declaration_instance37();
    specparam_declaration38 specparam_declaration_instance38();
    specparam_declaration39 specparam_declaration_instance39();
    specparam_declaration40 specparam_declaration_instance40();
    specparam_declaration41 specparam_declaration_instance41();
    specparam_declaration42 specparam_declaration_instance42();
    specparam_declaration43 specparam_declaration_instance43();
    specparam_declaration44 specparam_declaration_instance44();
    specparam_declaration45 specparam_declaration_instance45();
    specparam_declaration46 specparam_declaration_instance46();
    specparam_declaration47 specparam_declaration_instance47();
    specparam_declaration48 specparam_declaration_instance48();
    specparam_declaration49 specparam_declaration_instance49();
    specparam_declaration50 specparam_declaration_instance50();
    specparam_declaration51 specparam_declaration_instance51();
    specparam_declaration52 specparam_declaration_instance52();
    specparam_declaration53 specparam_declaration_instance53();
    specparam_declaration54 specparam_declaration_instance54();
    specparam_declaration55 specparam_declaration_instance55();
    specparam_declaration56 specparam_declaration_instance56();
    specparam_declaration57 specparam_declaration_instance57();
    specparam_declaration58 specparam_declaration_instance58();
    specparam_declaration59 specparam_declaration_instance59();
    specparam_declaration60 specparam_declaration_instance60();
    specparam_declaration61 specparam_declaration_instance61();
    specparam_declaration62 specparam_declaration_instance62();
    specparam_declaration63 specparam_declaration_instance63();
    specparam_declaration64 specparam_declaration_instance64();
    specparam_declaration65 specparam_declaration_instance65();
    specparam_declaration66 specparam_declaration_instance66();
    specparam_declaration67 specparam_declaration_instance67();
    specparam_declaration68 specparam_declaration_instance68();
    specparam_declaration69 specparam_declaration_instance69();
    specparam_declaration70 specparam_declaration_instance70();
    specparam_declaration71 specparam_declaration_instance71();
    specparam_declaration72 specparam_declaration_instance72();
    specparam_declaration73 specparam_declaration_instance73();
    specparam_declaration74 specparam_declaration_instance74();
    specparam_declaration75 specparam_declaration_instance75();
    specparam_declaration76 specparam_declaration_instance76();
    specparam_declaration77 specparam_declaration_instance77();
    specparam_declaration78 specparam_declaration_instance78();
    specparam_declaration79 specparam_declaration_instance79();
    specparam_declaration80 specparam_declaration_instance80();
    specparam_declaration81 specparam_declaration_instance81();
    specparam_declaration82 specparam_declaration_instance82();
    specparam_declaration83 specparam_declaration_instance83();
    specparam_declaration84 specparam_declaration_instance84();
    specparam_declaration85 specparam_declaration_instance85();
    specparam_declaration86 specparam_declaration_instance86();
    specparam_declaration87 specparam_declaration_instance87();
    specparam_declaration88 specparam_declaration_instance88();
    specparam_declaration89 specparam_declaration_instance89();
    specparam_declaration90 specparam_declaration_instance90();
    specparam_declaration91 specparam_declaration_instance91();
    specparam_declaration92 specparam_declaration_instance92();
    specparam_declaration93 specparam_declaration_instance93();
    specparam_declaration94 specparam_declaration_instance94();
    specparam_declaration95 specparam_declaration_instance95();
    specparam_declaration96 specparam_declaration_instance96();
    specparam_declaration97 specparam_declaration_instance97();
    specparam_declaration98 specparam_declaration_instance98();
    specparam_declaration99 specparam_declaration_instance99();
    specparam_declaration100 specparam_declaration_instance100();
    specparam_declaration101 specparam_declaration_instance101();
    specparam_declaration102 specparam_declaration_instance102();
    specparam_declaration103 specparam_declaration_instance103();
    specparam_declaration104 specparam_declaration_instance104();
    specparam_declaration105 specparam_declaration_instance105();
    specparam_declaration106 specparam_declaration_instance106();
    specparam_declaration107 specparam_declaration_instance107();
    specparam_declaration108 specparam_declaration_instance108();
    specparam_declaration109 specparam_declaration_instance109();
    specparam_declaration110 specparam_declaration_instance110();
    specparam_declaration111 specparam_declaration_instance111();
    specparam_declaration112 specparam_declaration_instance112();
    specparam_declaration113 specparam_declaration_instance113();
    specparam_declaration114 specparam_declaration_instance114();
    specparam_declaration115 specparam_declaration_instance115();
    specparam_declaration116 specparam_declaration_instance116();
    specparam_declaration117 specparam_declaration_instance117();
    specparam_declaration118 specparam_declaration_instance118();
    specparam_declaration119 specparam_declaration_instance119();
    specparam_declaration120 specparam_declaration_instance120();
    specparam_declaration121 specparam_declaration_instance121();
    specparam_declaration122 specparam_declaration_instance122();
    specparam_declaration123 specparam_declaration_instance123();
    specparam_declaration124 specparam_declaration_instance124();
    specparam_declaration125 specparam_declaration_instance125();
    specparam_declaration126 specparam_declaration_instance126();
    specparam_declaration127 specparam_declaration_instance127();
    specparam_declaration128 specparam_declaration_instance128();
    specparam_declaration129 specparam_declaration_instance129();
    specparam_declaration130 specparam_declaration_instance130();
    specparam_declaration131 specparam_declaration_instance131();
    specparam_declaration132 specparam_declaration_instance132();
    specparam_declaration133 specparam_declaration_instance133();
    specparam_declaration134 specparam_declaration_instance134();
    specparam_declaration135 specparam_declaration_instance135();
    specparam_declaration136 specparam_declaration_instance136();
    specparam_declaration137 specparam_declaration_instance137();
    specparam_declaration138 specparam_declaration_instance138();
    specparam_declaration139 specparam_declaration_instance139();
    specparam_declaration140 specparam_declaration_instance140();
    specparam_declaration141 specparam_declaration_instance141();
    specparam_declaration142 specparam_declaration_instance142();
    specparam_declaration143 specparam_declaration_instance143();
    specparam_declaration144 specparam_declaration_instance144();
    specparam_declaration145 specparam_declaration_instance145();
    specparam_declaration146 specparam_declaration_instance146();
    specparam_declaration147 specparam_declaration_instance147();
    specparam_declaration148 specparam_declaration_instance148();
    specparam_declaration149 specparam_declaration_instance149();
    specparam_declaration150 specparam_declaration_instance150();
    specparam_declaration151 specparam_declaration_instance151();
    specparam_declaration152 specparam_declaration_instance152();
    specparam_declaration153 specparam_declaration_instance153();
    specparam_declaration154 specparam_declaration_instance154();
    specparam_declaration155 specparam_declaration_instance155();
    specparam_declaration156 specparam_declaration_instance156();
    specparam_declaration157 specparam_declaration_instance157();
    specparam_declaration158 specparam_declaration_instance158();
    specparam_declaration159 specparam_declaration_instance159();
    specparam_declaration160 specparam_declaration_instance160();
    specparam_declaration161 specparam_declaration_instance161();
    specparam_declaration162 specparam_declaration_instance162();
    specparam_declaration163 specparam_declaration_instance163();
    specparam_declaration164 specparam_declaration_instance164();
    specparam_declaration165 specparam_declaration_instance165();
    specparam_declaration166 specparam_declaration_instance166();
    specparam_declaration167 specparam_declaration_instance167();
    specparam_declaration168 specparam_declaration_instance168();
    specparam_declaration169 specparam_declaration_instance169();
    specparam_declaration170 specparam_declaration_instance170();
    specparam_declaration171 specparam_declaration_instance171();
    specparam_declaration172 specparam_declaration_instance172();
    specparam_declaration173 specparam_declaration_instance173();
    specparam_declaration174 specparam_declaration_instance174();
    specparam_declaration175 specparam_declaration_instance175();
    specparam_declaration176 specparam_declaration_instance176();
    specparam_declaration177 specparam_declaration_instance177();
    specparam_declaration178 specparam_declaration_instance178();
    specparam_declaration179 specparam_declaration_instance179();
    specparam_declaration180 specparam_declaration_instance180();
    specparam_declaration181 specparam_declaration_instance181();
    specparam_declaration182 specparam_declaration_instance182();
    specparam_declaration183 specparam_declaration_instance183();
    specparam_declaration184 specparam_declaration_instance184();
    specparam_declaration185 specparam_declaration_instance185();
    specparam_declaration186 specparam_declaration_instance186();
    specparam_declaration187 specparam_declaration_instance187();
    specparam_declaration188 specparam_declaration_instance188();
    specparam_declaration189 specparam_declaration_instance189();
    specparam_declaration190 specparam_declaration_instance190();
    specparam_declaration191 specparam_declaration_instance191();
    specparam_declaration192 specparam_declaration_instance192();
    specparam_declaration193 specparam_declaration_instance193();
    specparam_declaration194 specparam_declaration_instance194();
    specparam_declaration195 specparam_declaration_instance195();
    specparam_declaration196 specparam_declaration_instance196();
    specparam_declaration197 specparam_declaration_instance197();
    specparam_declaration198 specparam_declaration_instance198();
    specparam_declaration199 specparam_declaration_instance199();
    specparam_declaration200 specparam_declaration_instance200();
    specparam_declaration201 specparam_declaration_instance201();
    specparam_declaration202 specparam_declaration_instance202();
    specparam_declaration203 specparam_declaration_instance203();
    specparam_declaration204 specparam_declaration_instance204();
    specparam_declaration205 specparam_declaration_instance205();
    specparam_declaration206 specparam_declaration_instance206();
    specparam_declaration207 specparam_declaration_instance207();
    specparam_declaration208 specparam_declaration_instance208();
    specparam_declaration209 specparam_declaration_instance209();
    specparam_declaration210 specparam_declaration_instance210();
    specparam_declaration211 specparam_declaration_instance211();
    specparam_declaration212 specparam_declaration_instance212();
    specparam_declaration213 specparam_declaration_instance213();
    specparam_declaration214 specparam_declaration_instance214();
    specparam_declaration215 specparam_declaration_instance215();
    specparam_declaration216 specparam_declaration_instance216();
    specparam_declaration217 specparam_declaration_instance217();
    specparam_declaration218 specparam_declaration_instance218();
    specparam_declaration219 specparam_declaration_instance219();
    specparam_declaration220 specparam_declaration_instance220();
    specparam_declaration221 specparam_declaration_instance221();
    specparam_declaration222 specparam_declaration_instance222();
    specparam_declaration223 specparam_declaration_instance223();
    specparam_declaration224 specparam_declaration_instance224();
    specparam_declaration225 specparam_declaration_instance225();
    specparam_declaration226 specparam_declaration_instance226();
    specparam_declaration227 specparam_declaration_instance227();
    specparam_declaration228 specparam_declaration_instance228();
    specparam_declaration229 specparam_declaration_instance229();
    specparam_declaration230 specparam_declaration_instance230();
    specparam_declaration231 specparam_declaration_instance231();
    specparam_declaration232 specparam_declaration_instance232();
    specparam_declaration233 specparam_declaration_instance233();
    specparam_declaration234 specparam_declaration_instance234();
    specparam_declaration235 specparam_declaration_instance235();
    specparam_declaration236 specparam_declaration_instance236();
    specparam_declaration237 specparam_declaration_instance237();
    specparam_declaration238 specparam_declaration_instance238();
    specparam_declaration239 specparam_declaration_instance239();
    specparam_declaration240 specparam_declaration_instance240();
    specparam_declaration241 specparam_declaration_instance241();
    specparam_declaration242 specparam_declaration_instance242();
    specparam_declaration243 specparam_declaration_instance243();
    specparam_declaration244 specparam_declaration_instance244();
    specparam_declaration245 specparam_declaration_instance245();
    specparam_declaration246 specparam_declaration_instance246();
    specparam_declaration247 specparam_declaration_instance247();
    specparam_declaration248 specparam_declaration_instance248();
    specparam_declaration249 specparam_declaration_instance249();
    specparam_declaration250 specparam_declaration_instance250();
    specparam_declaration251 specparam_declaration_instance251();
    specparam_declaration252 specparam_declaration_instance252();
    specparam_declaration253 specparam_declaration_instance253();
    specparam_declaration254 specparam_declaration_instance254();
    specparam_declaration255 specparam_declaration_instance255();
    specparam_declaration256 specparam_declaration_instance256();
    specparam_declaration257 specparam_declaration_instance257();
    specparam_declaration258 specparam_declaration_instance258();
    specparam_declaration259 specparam_declaration_instance259();
    specparam_declaration260 specparam_declaration_instance260();
    specparam_declaration261 specparam_declaration_instance261();
    specparam_declaration262 specparam_declaration_instance262();
    specparam_declaration263 specparam_declaration_instance263();
    specparam_declaration264 specparam_declaration_instance264();
    specparam_declaration265 specparam_declaration_instance265();
    specparam_declaration266 specparam_declaration_instance266();
    specparam_declaration267 specparam_declaration_instance267();
    specparam_declaration268 specparam_declaration_instance268();
    specparam_declaration269 specparam_declaration_instance269();
    specparam_declaration270 specparam_declaration_instance270();
    specparam_declaration271 specparam_declaration_instance271();
    specparam_declaration272 specparam_declaration_instance272();
    specparam_declaration273 specparam_declaration_instance273();
    specparam_declaration274 specparam_declaration_instance274();
    specparam_declaration275 specparam_declaration_instance275();
    specparam_declaration276 specparam_declaration_instance276();
    specparam_declaration277 specparam_declaration_instance277();
    specparam_declaration278 specparam_declaration_instance278();
    specparam_declaration279 specparam_declaration_instance279();
    specparam_declaration280 specparam_declaration_instance280();
    specparam_declaration281 specparam_declaration_instance281();
    specparam_declaration282 specparam_declaration_instance282();
    specparam_declaration283 specparam_declaration_instance283();
    specparam_declaration284 specparam_declaration_instance284();
    specparam_declaration285 specparam_declaration_instance285();
    specparam_declaration286 specparam_declaration_instance286();
    specparam_declaration287 specparam_declaration_instance287();
    specparam_declaration288 specparam_declaration_instance288();
    specparam_declaration289 specparam_declaration_instance289();
    specparam_declaration290 specparam_declaration_instance290();
    specparam_declaration291 specparam_declaration_instance291();
    specparam_declaration292 specparam_declaration_instance292();
    specparam_declaration293 specparam_declaration_instance293();
    specparam_declaration294 specparam_declaration_instance294();
    specparam_declaration295 specparam_declaration_instance295();
    specparam_declaration296 specparam_declaration_instance296();
    specparam_declaration297 specparam_declaration_instance297();
    specparam_declaration298 specparam_declaration_instance298();
    specparam_declaration299 specparam_declaration_instance299();
    specparam_declaration300 specparam_declaration_instance300();
    specparam_declaration301 specparam_declaration_instance301();
    specparam_declaration302 specparam_declaration_instance302();
    specparam_declaration303 specparam_declaration_instance303();
    specparam_declaration304 specparam_declaration_instance304();
    specparam_declaration305 specparam_declaration_instance305();
    specparam_declaration306 specparam_declaration_instance306();
    specparam_declaration307 specparam_declaration_instance307();
    specparam_declaration308 specparam_declaration_instance308();
    specparam_declaration309 specparam_declaration_instance309();
    specparam_declaration310 specparam_declaration_instance310();
    specparam_declaration311 specparam_declaration_instance311();
    specparam_declaration312 specparam_declaration_instance312();
    specparam_declaration313 specparam_declaration_instance313();
    specparam_declaration314 specparam_declaration_instance314();
    specparam_declaration315 specparam_declaration_instance315();
    specparam_declaration316 specparam_declaration_instance316();
    specparam_declaration317 specparam_declaration_instance317();
    specparam_declaration318 specparam_declaration_instance318();
    specparam_declaration319 specparam_declaration_instance319();
    specparam_declaration320 specparam_declaration_instance320();
    specparam_declaration321 specparam_declaration_instance321();
    specparam_declaration322 specparam_declaration_instance322();
    specparam_declaration323 specparam_declaration_instance323();
    specparam_declaration324 specparam_declaration_instance324();
    specparam_declaration325 specparam_declaration_instance325();
    specparam_declaration326 specparam_declaration_instance326();
    specparam_declaration327 specparam_declaration_instance327();
    specparam_declaration328 specparam_declaration_instance328();
    specparam_declaration329 specparam_declaration_instance329();
    specparam_declaration330 specparam_declaration_instance330();
    specparam_declaration331 specparam_declaration_instance331();
    specparam_declaration332 specparam_declaration_instance332();
    specparam_declaration333 specparam_declaration_instance333();
    specparam_declaration334 specparam_declaration_instance334();
    specparam_declaration335 specparam_declaration_instance335();
    specparam_declaration336 specparam_declaration_instance336();
    specparam_declaration337 specparam_declaration_instance337();
    specparam_declaration338 specparam_declaration_instance338();
    specparam_declaration339 specparam_declaration_instance339();
    specparam_declaration340 specparam_declaration_instance340();
    specparam_declaration341 specparam_declaration_instance341();
    specparam_declaration342 specparam_declaration_instance342();
    specparam_declaration343 specparam_declaration_instance343();
    specparam_declaration344 specparam_declaration_instance344();
    specparam_declaration345 specparam_declaration_instance345();
    specparam_declaration346 specparam_declaration_instance346();
    specparam_declaration347 specparam_declaration_instance347();
    specparam_declaration348 specparam_declaration_instance348();
    specparam_declaration349 specparam_declaration_instance349();
    specparam_declaration350 specparam_declaration_instance350();
    specparam_declaration351 specparam_declaration_instance351();
    specparam_declaration352 specparam_declaration_instance352();
    specparam_declaration353 specparam_declaration_instance353();
    specparam_declaration354 specparam_declaration_instance354();
    specparam_declaration355 specparam_declaration_instance355();
    specparam_declaration356 specparam_declaration_instance356();
    specparam_declaration357 specparam_declaration_instance357();
    specparam_declaration358 specparam_declaration_instance358();
    specparam_declaration359 specparam_declaration_instance359();
    specparam_declaration360 specparam_declaration_instance360();
    specparam_declaration361 specparam_declaration_instance361();
    specparam_declaration362 specparam_declaration_instance362();
    specparam_declaration363 specparam_declaration_instance363();
    specparam_declaration364 specparam_declaration_instance364();
    specparam_declaration365 specparam_declaration_instance365();
    specparam_declaration366 specparam_declaration_instance366();
    specparam_declaration367 specparam_declaration_instance367();
    specparam_declaration368 specparam_declaration_instance368();
    specparam_declaration369 specparam_declaration_instance369();
    specparam_declaration370 specparam_declaration_instance370();
    specparam_declaration371 specparam_declaration_instance371();
    specparam_declaration372 specparam_declaration_instance372();
    specparam_declaration373 specparam_declaration_instance373();
    specparam_declaration374 specparam_declaration_instance374();
    specparam_declaration375 specparam_declaration_instance375();
    specparam_declaration376 specparam_declaration_instance376();
    specparam_declaration377 specparam_declaration_instance377();
    specparam_declaration378 specparam_declaration_instance378();
    specparam_declaration379 specparam_declaration_instance379();
    specparam_declaration380 specparam_declaration_instance380();
    specparam_declaration381 specparam_declaration_instance381();
    specparam_declaration382 specparam_declaration_instance382();
    specparam_declaration383 specparam_declaration_instance383();
    specparam_declaration384 specparam_declaration_instance384();
    specparam_declaration385 specparam_declaration_instance385();
    specparam_declaration386 specparam_declaration_instance386();
    specparam_declaration387 specparam_declaration_instance387();
    specparam_declaration388 specparam_declaration_instance388();
    specparam_declaration389 specparam_declaration_instance389();
    specparam_declaration390 specparam_declaration_instance390();
    specparam_declaration391 specparam_declaration_instance391();
    specparam_declaration392 specparam_declaration_instance392();
    specparam_declaration393 specparam_declaration_instance393();
    specparam_declaration394 specparam_declaration_instance394();
    specparam_declaration395 specparam_declaration_instance395();
    specparam_declaration396 specparam_declaration_instance396();
    specparam_declaration397 specparam_declaration_instance397();
    specparam_declaration398 specparam_declaration_instance398();
    specparam_declaration399 specparam_declaration_instance399();
    specparam_declaration400 specparam_declaration_instance400();
    specparam_declaration401 specparam_declaration_instance401();
    specparam_declaration402 specparam_declaration_instance402();
    specparam_declaration403 specparam_declaration_instance403();
    specparam_declaration404 specparam_declaration_instance404();
    specparam_declaration405 specparam_declaration_instance405();
    specparam_declaration406 specparam_declaration_instance406();
    specparam_declaration407 specparam_declaration_instance407();
    specparam_declaration408 specparam_declaration_instance408();
    specparam_declaration409 specparam_declaration_instance409();
    specparam_declaration410 specparam_declaration_instance410();
    specparam_declaration411 specparam_declaration_instance411();
    specparam_declaration412 specparam_declaration_instance412();
    specparam_declaration413 specparam_declaration_instance413();
    specparam_declaration414 specparam_declaration_instance414();
    specparam_declaration415 specparam_declaration_instance415();
    specparam_declaration416 specparam_declaration_instance416();
    specparam_declaration417 specparam_declaration_instance417();
    specparam_declaration418 specparam_declaration_instance418();
    specparam_declaration419 specparam_declaration_instance419();
    specparam_declaration420 specparam_declaration_instance420();
    specparam_declaration421 specparam_declaration_instance421();
    specparam_declaration422 specparam_declaration_instance422();
    specparam_declaration423 specparam_declaration_instance423();
    specparam_declaration424 specparam_declaration_instance424();
    specparam_declaration425 specparam_declaration_instance425();
    specparam_declaration426 specparam_declaration_instance426();
    specparam_declaration427 specparam_declaration_instance427();
    specparam_declaration428 specparam_declaration_instance428();
    specparam_declaration429 specparam_declaration_instance429();
    specparam_declaration430 specparam_declaration_instance430();
    specparam_declaration431 specparam_declaration_instance431();
    specparam_declaration432 specparam_declaration_instance432();
    specparam_declaration433 specparam_declaration_instance433();
    specparam_declaration434 specparam_declaration_instance434();
    specparam_declaration435 specparam_declaration_instance435();
    specparam_declaration436 specparam_declaration_instance436();
    specparam_declaration437 specparam_declaration_instance437();
    specparam_declaration438 specparam_declaration_instance438();
    specparam_declaration439 specparam_declaration_instance439();
    specparam_declaration440 specparam_declaration_instance440();
    specparam_declaration441 specparam_declaration_instance441();
    specparam_declaration442 specparam_declaration_instance442();
    specparam_declaration443 specparam_declaration_instance443();
    specparam_declaration444 specparam_declaration_instance444();
    specparam_declaration445 specparam_declaration_instance445();
    specparam_declaration446 specparam_declaration_instance446();
    specparam_declaration447 specparam_declaration_instance447();
    specparam_declaration448 specparam_declaration_instance448();
    specparam_declaration449 specparam_declaration_instance449();
    specparam_declaration450 specparam_declaration_instance450();
    specparam_declaration451 specparam_declaration_instance451();
    specparam_declaration452 specparam_declaration_instance452();
    specparam_declaration453 specparam_declaration_instance453();
    specparam_declaration454 specparam_declaration_instance454();
    specparam_declaration455 specparam_declaration_instance455();
    specparam_declaration456 specparam_declaration_instance456();
    specparam_declaration457 specparam_declaration_instance457();
    specparam_declaration458 specparam_declaration_instance458();
    specparam_declaration459 specparam_declaration_instance459();
    specparam_declaration460 specparam_declaration_instance460();
    specparam_declaration461 specparam_declaration_instance461();
    specparam_declaration462 specparam_declaration_instance462();
    specparam_declaration463 specparam_declaration_instance463();
    specparam_declaration464 specparam_declaration_instance464();
    specparam_declaration465 specparam_declaration_instance465();
    specparam_declaration466 specparam_declaration_instance466();
    specparam_declaration467 specparam_declaration_instance467();
    specparam_declaration468 specparam_declaration_instance468();
    specparam_declaration469 specparam_declaration_instance469();
    specparam_declaration470 specparam_declaration_instance470();
    specparam_declaration471 specparam_declaration_instance471();
    specparam_declaration472 specparam_declaration_instance472();
    specparam_declaration473 specparam_declaration_instance473();
    specparam_declaration474 specparam_declaration_instance474();
    specparam_declaration475 specparam_declaration_instance475();
    specparam_declaration476 specparam_declaration_instance476();
    specparam_declaration477 specparam_declaration_instance477();
    specparam_declaration478 specparam_declaration_instance478();
    specparam_declaration479 specparam_declaration_instance479();
    specparam_declaration480 specparam_declaration_instance480();
    specparam_declaration481 specparam_declaration_instance481();
    specparam_declaration482 specparam_declaration_instance482();
    specparam_declaration483 specparam_declaration_instance483();
    specparam_declaration484 specparam_declaration_instance484();
    specparam_declaration485 specparam_declaration_instance485();
    specparam_declaration486 specparam_declaration_instance486();
    specparam_declaration487 specparam_declaration_instance487();
    specparam_declaration488 specparam_declaration_instance488();
    specparam_declaration489 specparam_declaration_instance489();
    specparam_declaration490 specparam_declaration_instance490();
    specparam_declaration491 specparam_declaration_instance491();
    specparam_declaration492 specparam_declaration_instance492();
    specparam_declaration493 specparam_declaration_instance493();
    specparam_declaration494 specparam_declaration_instance494();
    specparam_declaration495 specparam_declaration_instance495();
    specparam_declaration496 specparam_declaration_instance496();
    specparam_declaration497 specparam_declaration_instance497();
    specparam_declaration498 specparam_declaration_instance498();
    specparam_declaration499 specparam_declaration_instance499();
    specparam_declaration500 specparam_declaration_instance500();
    specparam_declaration501 specparam_declaration_instance501();
    specparam_declaration502 specparam_declaration_instance502();
    specparam_declaration503 specparam_declaration_instance503();
    specparam_declaration504 specparam_declaration_instance504();
    specparam_declaration505 specparam_declaration_instance505();
    specparam_declaration506 specparam_declaration_instance506();
    specparam_declaration507 specparam_declaration_instance507();
    specparam_declaration508 specparam_declaration_instance508();
    specparam_declaration509 specparam_declaration_instance509();
    specparam_declaration510 specparam_declaration_instance510();
    specparam_declaration511 specparam_declaration_instance511();
    specparam_declaration512 specparam_declaration_instance512();
    specparam_declaration513 specparam_declaration_instance513();
    specparam_declaration514 specparam_declaration_instance514();
    specparam_declaration515 specparam_declaration_instance515();
    specparam_declaration516 specparam_declaration_instance516();
    specparam_declaration517 specparam_declaration_instance517();
    specparam_declaration518 specparam_declaration_instance518();
    specparam_declaration519 specparam_declaration_instance519();
    specparam_declaration520 specparam_declaration_instance520();
    specparam_declaration521 specparam_declaration_instance521();
    specparam_declaration522 specparam_declaration_instance522();
    specparam_declaration523 specparam_declaration_instance523();
    specparam_declaration524 specparam_declaration_instance524();
    specparam_declaration525 specparam_declaration_instance525();
    specparam_declaration526 specparam_declaration_instance526();
    specparam_declaration527 specparam_declaration_instance527();
    specparam_declaration528 specparam_declaration_instance528();
    specparam_declaration529 specparam_declaration_instance529();
    specparam_declaration530 specparam_declaration_instance530();
    specparam_declaration531 specparam_declaration_instance531();
    specparam_declaration532 specparam_declaration_instance532();
    specparam_declaration533 specparam_declaration_instance533();
    specparam_declaration534 specparam_declaration_instance534();
    specparam_declaration535 specparam_declaration_instance535();
    specparam_declaration536 specparam_declaration_instance536();
    specparam_declaration537 specparam_declaration_instance537();
    specparam_declaration538 specparam_declaration_instance538();
    specparam_declaration539 specparam_declaration_instance539();
    specparam_declaration540 specparam_declaration_instance540();
    specparam_declaration541 specparam_declaration_instance541();
    specparam_declaration542 specparam_declaration_instance542();
    specparam_declaration543 specparam_declaration_instance543();
    specparam_declaration544 specparam_declaration_instance544();
    specparam_declaration545 specparam_declaration_instance545();
    specparam_declaration546 specparam_declaration_instance546();
    specparam_declaration547 specparam_declaration_instance547();
    specparam_declaration548 specparam_declaration_instance548();
    specparam_declaration549 specparam_declaration_instance549();
    specparam_declaration550 specparam_declaration_instance550();
    specparam_declaration551 specparam_declaration_instance551();
    specparam_declaration552 specparam_declaration_instance552();
    specparam_declaration553 specparam_declaration_instance553();
    specparam_declaration554 specparam_declaration_instance554();
    specparam_declaration555 specparam_declaration_instance555();
    specparam_declaration556 specparam_declaration_instance556();
    specparam_declaration557 specparam_declaration_instance557();
    specparam_declaration558 specparam_declaration_instance558();
    specparam_declaration559 specparam_declaration_instance559();
    specparam_declaration560 specparam_declaration_instance560();
    specparam_declaration561 specparam_declaration_instance561();
    specparam_declaration562 specparam_declaration_instance562();
    specparam_declaration563 specparam_declaration_instance563();
    specparam_declaration564 specparam_declaration_instance564();
    specparam_declaration565 specparam_declaration_instance565();
    specparam_declaration566 specparam_declaration_instance566();
    specparam_declaration567 specparam_declaration_instance567();
    specparam_declaration568 specparam_declaration_instance568();
    specparam_declaration569 specparam_declaration_instance569();
    specparam_declaration570 specparam_declaration_instance570();
    specparam_declaration571 specparam_declaration_instance571();
    specparam_declaration572 specparam_declaration_instance572();
    specparam_declaration573 specparam_declaration_instance573();
    specparam_declaration574 specparam_declaration_instance574();
    specparam_declaration575 specparam_declaration_instance575();
    specparam_declaration576 specparam_declaration_instance576();
    specparam_declaration577 specparam_declaration_instance577();
    specparam_declaration578 specparam_declaration_instance578();
    specparam_declaration579 specparam_declaration_instance579();
    specparam_declaration580 specparam_declaration_instance580();
    specparam_declaration581 specparam_declaration_instance581();
    specparam_declaration582 specparam_declaration_instance582();
    specparam_declaration583 specparam_declaration_instance583();
    specparam_declaration584 specparam_declaration_instance584();
    specparam_declaration585 specparam_declaration_instance585();
    specparam_declaration586 specparam_declaration_instance586();
    specparam_declaration587 specparam_declaration_instance587();
    specparam_declaration588 specparam_declaration_instance588();
    specparam_declaration589 specparam_declaration_instance589();
    specparam_declaration590 specparam_declaration_instance590();
    specparam_declaration591 specparam_declaration_instance591();
    specparam_declaration592 specparam_declaration_instance592();
    specparam_declaration593 specparam_declaration_instance593();
    specparam_declaration594 specparam_declaration_instance594();
    specparam_declaration595 specparam_declaration_instance595();
    specparam_declaration596 specparam_declaration_instance596();
    specparam_declaration597 specparam_declaration_instance597();
    specparam_declaration598 specparam_declaration_instance598();
    specparam_declaration599 specparam_declaration_instance599();
    specparam_declaration600 specparam_declaration_instance600();
    specparam_declaration601 specparam_declaration_instance601();
    specparam_declaration602 specparam_declaration_instance602();
    specparam_declaration603 specparam_declaration_instance603();
    specparam_declaration604 specparam_declaration_instance604();
    specparam_declaration605 specparam_declaration_instance605();
    specparam_declaration606 specparam_declaration_instance606();
    specparam_declaration607 specparam_declaration_instance607();
    specparam_declaration608 specparam_declaration_instance608();
    specparam_declaration609 specparam_declaration_instance609();
    specparam_declaration610 specparam_declaration_instance610();
    specparam_declaration611 specparam_declaration_instance611();
    specparam_declaration612 specparam_declaration_instance612();
    specparam_declaration613 specparam_declaration_instance613();
    specparam_declaration614 specparam_declaration_instance614();
    specparam_declaration615 specparam_declaration_instance615();
    specparam_declaration616 specparam_declaration_instance616();
    specparam_declaration617 specparam_declaration_instance617();
    specparam_declaration618 specparam_declaration_instance618();
    specparam_declaration619 specparam_declaration_instance619();
    specparam_declaration620 specparam_declaration_instance620();
    specparam_declaration621 specparam_declaration_instance621();
    specparam_declaration622 specparam_declaration_instance622();
    specparam_declaration623 specparam_declaration_instance623();
    specparam_declaration624 specparam_declaration_instance624();
    specparam_declaration625 specparam_declaration_instance625();
    specparam_declaration626 specparam_declaration_instance626();
    specparam_declaration627 specparam_declaration_instance627();
    specparam_declaration628 specparam_declaration_instance628();
    specparam_declaration629 specparam_declaration_instance629();
    specparam_declaration630 specparam_declaration_instance630();
    specparam_declaration631 specparam_declaration_instance631();
    specparam_declaration632 specparam_declaration_instance632();
    specparam_declaration633 specparam_declaration_instance633();
    specparam_declaration634 specparam_declaration_instance634();
    specparam_declaration635 specparam_declaration_instance635();
    specparam_declaration636 specparam_declaration_instance636();
    specparam_declaration637 specparam_declaration_instance637();
    specparam_declaration638 specparam_declaration_instance638();
    specparam_declaration639 specparam_declaration_instance639();
    specparam_declaration640 specparam_declaration_instance640();
    specparam_declaration641 specparam_declaration_instance641();
    specparam_declaration642 specparam_declaration_instance642();
    specparam_declaration643 specparam_declaration_instance643();
    specparam_declaration644 specparam_declaration_instance644();
    specparam_declaration645 specparam_declaration_instance645();
    specparam_declaration646 specparam_declaration_instance646();
    specparam_declaration647 specparam_declaration_instance647();
    specparam_declaration648 specparam_declaration_instance648();
    specparam_declaration649 specparam_declaration_instance649();
    specparam_declaration650 specparam_declaration_instance650();
    specparam_declaration651 specparam_declaration_instance651();
    specparam_declaration652 specparam_declaration_instance652();
    specparam_declaration653 specparam_declaration_instance653();
    specparam_declaration654 specparam_declaration_instance654();
    specparam_declaration655 specparam_declaration_instance655();
    specparam_declaration656 specparam_declaration_instance656();
    specparam_declaration657 specparam_declaration_instance657();
    specparam_declaration658 specparam_declaration_instance658();
    specparam_declaration659 specparam_declaration_instance659();
    specparam_declaration660 specparam_declaration_instance660();
    specparam_declaration661 specparam_declaration_instance661();
    specparam_declaration662 specparam_declaration_instance662();
    specparam_declaration663 specparam_declaration_instance663();
    specparam_declaration664 specparam_declaration_instance664();
    specparam_declaration665 specparam_declaration_instance665();
    specparam_declaration666 specparam_declaration_instance666();
    specparam_declaration667 specparam_declaration_instance667();
    specparam_declaration668 specparam_declaration_instance668();
    specparam_declaration669 specparam_declaration_instance669();
    specparam_declaration670 specparam_declaration_instance670();
    specparam_declaration671 specparam_declaration_instance671();
    specparam_declaration672 specparam_declaration_instance672();
    specparam_declaration673 specparam_declaration_instance673();
    specparam_declaration674 specparam_declaration_instance674();
    specparam_declaration675 specparam_declaration_instance675();
    specparam_declaration676 specparam_declaration_instance676();
    specparam_declaration677 specparam_declaration_instance677();
    specparam_declaration678 specparam_declaration_instance678();
    specparam_declaration679 specparam_declaration_instance679();
    specparam_declaration680 specparam_declaration_instance680();
    specparam_declaration681 specparam_declaration_instance681();
    specparam_declaration682 specparam_declaration_instance682();
    specparam_declaration683 specparam_declaration_instance683();
    specparam_declaration684 specparam_declaration_instance684();
    specparam_declaration685 specparam_declaration_instance685();
    specparam_declaration686 specparam_declaration_instance686();
    specparam_declaration687 specparam_declaration_instance687();
    specparam_declaration688 specparam_declaration_instance688();
    specparam_declaration689 specparam_declaration_instance689();
    specparam_declaration690 specparam_declaration_instance690();
    specparam_declaration691 specparam_declaration_instance691();
    specparam_declaration692 specparam_declaration_instance692();
    specparam_declaration693 specparam_declaration_instance693();
    specparam_declaration694 specparam_declaration_instance694();
    specparam_declaration695 specparam_declaration_instance695();
    specparam_declaration696 specparam_declaration_instance696();
    specparam_declaration697 specparam_declaration_instance697();
    specparam_declaration698 specparam_declaration_instance698();
    specparam_declaration699 specparam_declaration_instance699();
    specparam_declaration700 specparam_declaration_instance700();
    specparam_declaration701 specparam_declaration_instance701();
    specparam_declaration702 specparam_declaration_instance702();
    specparam_declaration703 specparam_declaration_instance703();
    specparam_declaration704 specparam_declaration_instance704();
    specparam_declaration705 specparam_declaration_instance705();
    specparam_declaration706 specparam_declaration_instance706();
    specparam_declaration707 specparam_declaration_instance707();
    specparam_declaration708 specparam_declaration_instance708();
    specparam_declaration709 specparam_declaration_instance709();
    specparam_declaration710 specparam_declaration_instance710();
    specparam_declaration711 specparam_declaration_instance711();
    specparam_declaration712 specparam_declaration_instance712();
    specparam_declaration713 specparam_declaration_instance713();
    specparam_declaration714 specparam_declaration_instance714();
    specparam_declaration715 specparam_declaration_instance715();
    specparam_declaration716 specparam_declaration_instance716();
    specparam_declaration717 specparam_declaration_instance717();
    specparam_declaration718 specparam_declaration_instance718();
    specparam_declaration719 specparam_declaration_instance719();
    specparam_declaration720 specparam_declaration_instance720();
    specparam_declaration721 specparam_declaration_instance721();
    specparam_declaration722 specparam_declaration_instance722();
    specparam_declaration723 specparam_declaration_instance723();
    specparam_declaration724 specparam_declaration_instance724();
    specparam_declaration725 specparam_declaration_instance725();
    specparam_declaration726 specparam_declaration_instance726();
    specparam_declaration727 specparam_declaration_instance727();
    specparam_declaration728 specparam_declaration_instance728();
    specparam_declaration729 specparam_declaration_instance729();
    specparam_declaration730 specparam_declaration_instance730();
    specparam_declaration731 specparam_declaration_instance731();
    specparam_declaration732 specparam_declaration_instance732();
    specparam_declaration733 specparam_declaration_instance733();
    specparam_declaration734 specparam_declaration_instance734();
    specparam_declaration735 specparam_declaration_instance735();
    specparam_declaration736 specparam_declaration_instance736();
    specparam_declaration737 specparam_declaration_instance737();
    specparam_declaration738 specparam_declaration_instance738();
    specparam_declaration739 specparam_declaration_instance739();
    specparam_declaration740 specparam_declaration_instance740();
    specparam_declaration741 specparam_declaration_instance741();
    specparam_declaration742 specparam_declaration_instance742();
    specparam_declaration743 specparam_declaration_instance743();
    specparam_declaration744 specparam_declaration_instance744();
    specparam_declaration745 specparam_declaration_instance745();
    specparam_declaration746 specparam_declaration_instance746();
    specparam_declaration747 specparam_declaration_instance747();
    specparam_declaration748 specparam_declaration_instance748();
    specparam_declaration749 specparam_declaration_instance749();
    specparam_declaration750 specparam_declaration_instance750();
    specparam_declaration751 specparam_declaration_instance751();
    specparam_declaration752 specparam_declaration_instance752();
    specparam_declaration753 specparam_declaration_instance753();
    specparam_declaration754 specparam_declaration_instance754();
    specparam_declaration755 specparam_declaration_instance755();
    specparam_declaration756 specparam_declaration_instance756();
    specparam_declaration757 specparam_declaration_instance757();
    specparam_declaration758 specparam_declaration_instance758();
    specparam_declaration759 specparam_declaration_instance759();
    specparam_declaration760 specparam_declaration_instance760();
    specparam_declaration761 specparam_declaration_instance761();
    specparam_declaration762 specparam_declaration_instance762();
    specparam_declaration763 specparam_declaration_instance763();
    specparam_declaration764 specparam_declaration_instance764();
    specparam_declaration765 specparam_declaration_instance765();
    specparam_declaration766 specparam_declaration_instance766();
    specparam_declaration767 specparam_declaration_instance767();
    specparam_declaration768 specparam_declaration_instance768();
    specparam_declaration769 specparam_declaration_instance769();
    specparam_declaration770 specparam_declaration_instance770();
    specparam_declaration771 specparam_declaration_instance771();
    specparam_declaration772 specparam_declaration_instance772();
    specparam_declaration773 specparam_declaration_instance773();
    specparam_declaration774 specparam_declaration_instance774();
    specparam_declaration775 specparam_declaration_instance775();
    specparam_declaration776 specparam_declaration_instance776();
    specparam_declaration777 specparam_declaration_instance777();
    specparam_declaration778 specparam_declaration_instance778();
    specparam_declaration779 specparam_declaration_instance779();
    specparam_declaration780 specparam_declaration_instance780();
    specparam_declaration781 specparam_declaration_instance781();
    specparam_declaration782 specparam_declaration_instance782();
    specparam_declaration783 specparam_declaration_instance783();
    specparam_declaration784 specparam_declaration_instance784();
    specparam_declaration785 specparam_declaration_instance785();
    specparam_declaration786 specparam_declaration_instance786();
    specparam_declaration787 specparam_declaration_instance787();
    specparam_declaration788 specparam_declaration_instance788();
    specparam_declaration789 specparam_declaration_instance789();
    specparam_declaration790 specparam_declaration_instance790();
    specparam_declaration791 specparam_declaration_instance791();
    specparam_declaration792 specparam_declaration_instance792();
    specparam_declaration793 specparam_declaration_instance793();
    specparam_declaration794 specparam_declaration_instance794();
    specparam_declaration795 specparam_declaration_instance795();
    specparam_declaration796 specparam_declaration_instance796();
    specparam_declaration797 specparam_declaration_instance797();
    specparam_declaration798 specparam_declaration_instance798();
    specparam_declaration799 specparam_declaration_instance799();
    specparam_declaration800 specparam_declaration_instance800();
    specparam_declaration801 specparam_declaration_instance801();
    specparam_declaration802 specparam_declaration_instance802();
    specparam_declaration803 specparam_declaration_instance803();
    specparam_declaration804 specparam_declaration_instance804();
    specparam_declaration805 specparam_declaration_instance805();
    specparam_declaration806 specparam_declaration_instance806();
    specparam_declaration807 specparam_declaration_instance807();
    specparam_declaration808 specparam_declaration_instance808();
    specparam_declaration809 specparam_declaration_instance809();
    specparam_declaration810 specparam_declaration_instance810();
    specparam_declaration811 specparam_declaration_instance811();
    specparam_declaration812 specparam_declaration_instance812();
    specparam_declaration813 specparam_declaration_instance813();
    specparam_declaration814 specparam_declaration_instance814();
    specparam_declaration815 specparam_declaration_instance815();
    specparam_declaration816 specparam_declaration_instance816();
    specparam_declaration817 specparam_declaration_instance817();
    specparam_declaration818 specparam_declaration_instance818();
    specparam_declaration819 specparam_declaration_instance819();
    specparam_declaration820 specparam_declaration_instance820();
    specparam_declaration821 specparam_declaration_instance821();
    specparam_declaration822 specparam_declaration_instance822();
    specparam_declaration823 specparam_declaration_instance823();
    specparam_declaration824 specparam_declaration_instance824();
    specparam_declaration825 specparam_declaration_instance825();
    specparam_declaration826 specparam_declaration_instance826();
    specparam_declaration827 specparam_declaration_instance827();
    specparam_declaration828 specparam_declaration_instance828();
    specparam_declaration829 specparam_declaration_instance829();
    specparam_declaration830 specparam_declaration_instance830();
    specparam_declaration831 specparam_declaration_instance831();
    specparam_declaration832 specparam_declaration_instance832();
    specparam_declaration833 specparam_declaration_instance833();
    specparam_declaration834 specparam_declaration_instance834();
    specparam_declaration835 specparam_declaration_instance835();
    specparam_declaration836 specparam_declaration_instance836();
    specparam_declaration837 specparam_declaration_instance837();
    specparam_declaration838 specparam_declaration_instance838();
    specparam_declaration839 specparam_declaration_instance839();
    specparam_declaration840 specparam_declaration_instance840();
    specparam_declaration841 specparam_declaration_instance841();
    specparam_declaration842 specparam_declaration_instance842();
    specparam_declaration843 specparam_declaration_instance843();
    specparam_declaration844 specparam_declaration_instance844();
    specparam_declaration845 specparam_declaration_instance845();
    specparam_declaration846 specparam_declaration_instance846();
    specparam_declaration847 specparam_declaration_instance847();
    specparam_declaration848 specparam_declaration_instance848();
    specparam_declaration849 specparam_declaration_instance849();
    specparam_declaration850 specparam_declaration_instance850();
    specparam_declaration851 specparam_declaration_instance851();
    specparam_declaration852 specparam_declaration_instance852();
    specparam_declaration853 specparam_declaration_instance853();
    specparam_declaration854 specparam_declaration_instance854();
    specparam_declaration855 specparam_declaration_instance855();
    specparam_declaration856 specparam_declaration_instance856();
    specparam_declaration857 specparam_declaration_instance857();
    specparam_declaration858 specparam_declaration_instance858();
    specparam_declaration859 specparam_declaration_instance859();
    specparam_declaration860 specparam_declaration_instance860();
    specparam_declaration861 specparam_declaration_instance861();
    specparam_declaration862 specparam_declaration_instance862();
    specparam_declaration863 specparam_declaration_instance863();
    specparam_declaration864 specparam_declaration_instance864();
    specparam_declaration865 specparam_declaration_instance865();
    specparam_declaration866 specparam_declaration_instance866();
    specparam_declaration867 specparam_declaration_instance867();
    specparam_declaration868 specparam_declaration_instance868();
    specparam_declaration869 specparam_declaration_instance869();
    specparam_declaration870 specparam_declaration_instance870();
    specparam_declaration871 specparam_declaration_instance871();
    specparam_declaration872 specparam_declaration_instance872();
    specparam_declaration873 specparam_declaration_instance873();
    specparam_declaration874 specparam_declaration_instance874();
    specparam_declaration875 specparam_declaration_instance875();
    specparam_declaration876 specparam_declaration_instance876();
    specparam_declaration877 specparam_declaration_instance877();
    specparam_declaration878 specparam_declaration_instance878();
    specparam_declaration879 specparam_declaration_instance879();
    specparam_declaration880 specparam_declaration_instance880();
    specparam_declaration881 specparam_declaration_instance881();
    specparam_declaration882 specparam_declaration_instance882();
    specparam_declaration883 specparam_declaration_instance883();
    specparam_declaration884 specparam_declaration_instance884();
    specparam_declaration885 specparam_declaration_instance885();
    specparam_declaration886 specparam_declaration_instance886();
    specparam_declaration887 specparam_declaration_instance887();
    specparam_declaration888 specparam_declaration_instance888();
    specparam_declaration889 specparam_declaration_instance889();
    specparam_declaration890 specparam_declaration_instance890();
    specparam_declaration891 specparam_declaration_instance891();
    specparam_declaration892 specparam_declaration_instance892();
    specparam_declaration893 specparam_declaration_instance893();
    specparam_declaration894 specparam_declaration_instance894();
    specparam_declaration895 specparam_declaration_instance895();
    specparam_declaration896 specparam_declaration_instance896();
    specparam_declaration897 specparam_declaration_instance897();
    specparam_declaration898 specparam_declaration_instance898();
    specparam_declaration899 specparam_declaration_instance899();
    specparam_declaration900 specparam_declaration_instance900();
    specparam_declaration901 specparam_declaration_instance901();
    specparam_declaration902 specparam_declaration_instance902();
    specparam_declaration903 specparam_declaration_instance903();
    specparam_declaration904 specparam_declaration_instance904();
    specparam_declaration905 specparam_declaration_instance905();
    specparam_declaration906 specparam_declaration_instance906();
    specparam_declaration907 specparam_declaration_instance907();
    specparam_declaration908 specparam_declaration_instance908();
    specparam_declaration909 specparam_declaration_instance909();
    specparam_declaration910 specparam_declaration_instance910();
    specparam_declaration911 specparam_declaration_instance911();
    specparam_declaration912 specparam_declaration_instance912();
    specparam_declaration913 specparam_declaration_instance913();
    specparam_declaration914 specparam_declaration_instance914();
    specparam_declaration915 specparam_declaration_instance915();
    specparam_declaration916 specparam_declaration_instance916();
    specparam_declaration917 specparam_declaration_instance917();
    specparam_declaration918 specparam_declaration_instance918();
    specparam_declaration919 specparam_declaration_instance919();
    specparam_declaration920 specparam_declaration_instance920();
    specparam_declaration921 specparam_declaration_instance921();
    specparam_declaration922 specparam_declaration_instance922();
    specparam_declaration923 specparam_declaration_instance923();
    specparam_declaration924 specparam_declaration_instance924();
    specparam_declaration925 specparam_declaration_instance925();
    specparam_declaration926 specparam_declaration_instance926();
    specparam_declaration927 specparam_declaration_instance927();
    specparam_declaration928 specparam_declaration_instance928();
    specparam_declaration929 specparam_declaration_instance929();
    specparam_declaration930 specparam_declaration_instance930();
    specparam_declaration931 specparam_declaration_instance931();
    specparam_declaration932 specparam_declaration_instance932();
    specparam_declaration933 specparam_declaration_instance933();
    specparam_declaration934 specparam_declaration_instance934();
    specparam_declaration935 specparam_declaration_instance935();
    specparam_declaration936 specparam_declaration_instance936();
    specparam_declaration937 specparam_declaration_instance937();
    specparam_declaration938 specparam_declaration_instance938();
    specparam_declaration939 specparam_declaration_instance939();
    specparam_declaration940 specparam_declaration_instance940();
    specparam_declaration941 specparam_declaration_instance941();
    specparam_declaration942 specparam_declaration_instance942();
    specparam_declaration943 specparam_declaration_instance943();
    specparam_declaration944 specparam_declaration_instance944();
    specparam_declaration945 specparam_declaration_instance945();
    specparam_declaration946 specparam_declaration_instance946();
    specparam_declaration947 specparam_declaration_instance947();
    specparam_declaration948 specparam_declaration_instance948();
    specparam_declaration949 specparam_declaration_instance949();
    specparam_declaration950 specparam_declaration_instance950();
    specparam_declaration951 specparam_declaration_instance951();
    specparam_declaration952 specparam_declaration_instance952();
    specparam_declaration953 specparam_declaration_instance953();
    specparam_declaration954 specparam_declaration_instance954();
    specparam_declaration955 specparam_declaration_instance955();
    specparam_declaration956 specparam_declaration_instance956();
    specparam_declaration957 specparam_declaration_instance957();
    specparam_declaration958 specparam_declaration_instance958();
    specparam_declaration959 specparam_declaration_instance959();
    specparam_declaration960 specparam_declaration_instance960();
    specparam_declaration961 specparam_declaration_instance961();
    specparam_declaration962 specparam_declaration_instance962();
    specparam_declaration963 specparam_declaration_instance963();
    specparam_declaration964 specparam_declaration_instance964();
    specparam_declaration965 specparam_declaration_instance965();
    specparam_declaration966 specparam_declaration_instance966();
    specparam_declaration967 specparam_declaration_instance967();
    specparam_declaration968 specparam_declaration_instance968();
    specparam_declaration969 specparam_declaration_instance969();
    specparam_declaration970 specparam_declaration_instance970();
    specparam_declaration971 specparam_declaration_instance971();
    specparam_declaration972 specparam_declaration_instance972();
    specparam_declaration973 specparam_declaration_instance973();
    specparam_declaration974 specparam_declaration_instance974();
    specparam_declaration975 specparam_declaration_instance975();
    specparam_declaration976 specparam_declaration_instance976();
    specparam_declaration977 specparam_declaration_instance977();
    specparam_declaration978 specparam_declaration_instance978();
    specparam_declaration979 specparam_declaration_instance979();
    specparam_declaration980 specparam_declaration_instance980();
    specparam_declaration981 specparam_declaration_instance981();
    specparam_declaration982 specparam_declaration_instance982();
    specparam_declaration983 specparam_declaration_instance983();
    specparam_declaration984 specparam_declaration_instance984();
    specparam_declaration985 specparam_declaration_instance985();
    specparam_declaration986 specparam_declaration_instance986();
    specparam_declaration987 specparam_declaration_instance987();
    specparam_declaration988 specparam_declaration_instance988();
    specparam_declaration989 specparam_declaration_instance989();
    specparam_declaration990 specparam_declaration_instance990();
    specparam_declaration991 specparam_declaration_instance991();
    specparam_declaration992 specparam_declaration_instance992();
    specparam_declaration993 specparam_declaration_instance993();
    specparam_declaration994 specparam_declaration_instance994();
    specparam_declaration995 specparam_declaration_instance995();
    specparam_declaration996 specparam_declaration_instance996();
    specparam_declaration997 specparam_declaration_instance997();
    specparam_declaration998 specparam_declaration_instance998();
    specparam_declaration999 specparam_declaration_instance999();
    specparam_declaration1000 specparam_declaration_instance1000();
    specparam_declaration1001 specparam_declaration_instance1001();
    specparam_declaration1002 specparam_declaration_instance1002();
    specparam_declaration1003 specparam_declaration_instance1003();
    specparam_declaration1004 specparam_declaration_instance1004();
    specparam_declaration1005 specparam_declaration_instance1005();
    specparam_declaration1006 specparam_declaration_instance1006();
    specparam_declaration1007 specparam_declaration_instance1007();
    specparam_declaration1008 specparam_declaration_instance1008();
    specparam_declaration1009 specparam_declaration_instance1009();
    specparam_declaration1010 specparam_declaration_instance1010();
    specparam_declaration1011 specparam_declaration_instance1011();
    specparam_declaration1012 specparam_declaration_instance1012();
    specparam_declaration1013 specparam_declaration_instance1013();
    specparam_declaration1014 specparam_declaration_instance1014();
    specparam_declaration1015 specparam_declaration_instance1015();
    specparam_declaration1016 specparam_declaration_instance1016();
    specparam_declaration1017 specparam_declaration_instance1017();
    specparam_declaration1018 specparam_declaration_instance1018();
    specparam_declaration1019 specparam_declaration_instance1019();
    specparam_declaration1020 specparam_declaration_instance1020();
    specparam_declaration1021 specparam_declaration_instance1021();
    specparam_declaration1022 specparam_declaration_instance1022();
    specparam_declaration1023 specparam_declaration_instance1023();
    specparam_declaration1024 specparam_declaration_instance1024();
    specparam_declaration1025 specparam_declaration_instance1025();
    specparam_declaration1026 specparam_declaration_instance1026();
    specparam_declaration1027 specparam_declaration_instance1027();
    specparam_declaration1028 specparam_declaration_instance1028();
    specparam_declaration1029 specparam_declaration_instance1029();
    specparam_declaration1030 specparam_declaration_instance1030();
    specparam_declaration1031 specparam_declaration_instance1031();
    specparam_declaration1032 specparam_declaration_instance1032();
    specparam_declaration1033 specparam_declaration_instance1033();
    specparam_declaration1034 specparam_declaration_instance1034();
    specparam_declaration1035 specparam_declaration_instance1035();
    specparam_declaration1036 specparam_declaration_instance1036();
    specparam_declaration1037 specparam_declaration_instance1037();
    specparam_declaration1038 specparam_declaration_instance1038();
    specparam_declaration1039 specparam_declaration_instance1039();
    specparam_declaration1040 specparam_declaration_instance1040();
    specparam_declaration1041 specparam_declaration_instance1041();
    specparam_declaration1042 specparam_declaration_instance1042();
    specparam_declaration1043 specparam_declaration_instance1043();
    specparam_declaration1044 specparam_declaration_instance1044();
    specparam_declaration1045 specparam_declaration_instance1045();
    specparam_declaration1046 specparam_declaration_instance1046();
    specparam_declaration1047 specparam_declaration_instance1047();
    specparam_declaration1048 specparam_declaration_instance1048();
    specparam_declaration1049 specparam_declaration_instance1049();
    specparam_declaration1050 specparam_declaration_instance1050();
    specparam_declaration1051 specparam_declaration_instance1051();
    specparam_declaration1052 specparam_declaration_instance1052();
    specparam_declaration1053 specparam_declaration_instance1053();
    specparam_declaration1054 specparam_declaration_instance1054();
    specparam_declaration1055 specparam_declaration_instance1055();
    specparam_declaration1056 specparam_declaration_instance1056();
    specparam_declaration1057 specparam_declaration_instance1057();
    specparam_declaration1058 specparam_declaration_instance1058();
    specparam_declaration1059 specparam_declaration_instance1059();
    specparam_declaration1060 specparam_declaration_instance1060();
    specparam_declaration1061 specparam_declaration_instance1061();
    specparam_declaration1062 specparam_declaration_instance1062();
    specparam_declaration1063 specparam_declaration_instance1063();
    specparam_declaration1064 specparam_declaration_instance1064();
    specparam_declaration1065 specparam_declaration_instance1065();
    specparam_declaration1066 specparam_declaration_instance1066();
    specparam_declaration1067 specparam_declaration_instance1067();
    specparam_declaration1068 specparam_declaration_instance1068();
    specparam_declaration1069 specparam_declaration_instance1069();
    specparam_declaration1070 specparam_declaration_instance1070();
    specparam_declaration1071 specparam_declaration_instance1071();
    specparam_declaration1072 specparam_declaration_instance1072();
    specparam_declaration1073 specparam_declaration_instance1073();
    specparam_declaration1074 specparam_declaration_instance1074();
    specparam_declaration1075 specparam_declaration_instance1075();
    specparam_declaration1076 specparam_declaration_instance1076();
    specparam_declaration1077 specparam_declaration_instance1077();
    specparam_declaration1078 specparam_declaration_instance1078();
    specparam_declaration1079 specparam_declaration_instance1079();
    specparam_declaration1080 specparam_declaration_instance1080();
    specparam_declaration1081 specparam_declaration_instance1081();
    specparam_declaration1082 specparam_declaration_instance1082();
    specparam_declaration1083 specparam_declaration_instance1083();
    specparam_declaration1084 specparam_declaration_instance1084();
    specparam_declaration1085 specparam_declaration_instance1085();
    specparam_declaration1086 specparam_declaration_instance1086();
    specparam_declaration1087 specparam_declaration_instance1087();
    specparam_declaration1088 specparam_declaration_instance1088();
    specparam_declaration1089 specparam_declaration_instance1089();
    specparam_declaration1090 specparam_declaration_instance1090();
    specparam_declaration1091 specparam_declaration_instance1091();
    specparam_declaration1092 specparam_declaration_instance1092();
    specparam_declaration1093 specparam_declaration_instance1093();
    specparam_declaration1094 specparam_declaration_instance1094();
    specparam_declaration1095 specparam_declaration_instance1095();
    specparam_declaration1096 specparam_declaration_instance1096();
    specparam_declaration1097 specparam_declaration_instance1097();
    specparam_declaration1098 specparam_declaration_instance1098();
    specparam_declaration1099 specparam_declaration_instance1099();
    specparam_declaration1100 specparam_declaration_instance1100();
    specparam_declaration1101 specparam_declaration_instance1101();
    specparam_declaration1102 specparam_declaration_instance1102();
    specparam_declaration1103 specparam_declaration_instance1103();
    specparam_declaration1104 specparam_declaration_instance1104();
    specparam_declaration1105 specparam_declaration_instance1105();
    specparam_declaration1106 specparam_declaration_instance1106();
    specparam_declaration1107 specparam_declaration_instance1107();
    specparam_declaration1108 specparam_declaration_instance1108();
    specparam_declaration1109 specparam_declaration_instance1109();
    specparam_declaration1110 specparam_declaration_instance1110();
    specparam_declaration1111 specparam_declaration_instance1111();
    specparam_declaration1112 specparam_declaration_instance1112();
    specparam_declaration1113 specparam_declaration_instance1113();
    specparam_declaration1114 specparam_declaration_instance1114();
    specparam_declaration1115 specparam_declaration_instance1115();
    specparam_declaration1116 specparam_declaration_instance1116();
    specparam_declaration1117 specparam_declaration_instance1117();
    specparam_declaration1118 specparam_declaration_instance1118();
    specparam_declaration1119 specparam_declaration_instance1119();
    specparam_declaration1120 specparam_declaration_instance1120();
    specparam_declaration1121 specparam_declaration_instance1121();
    specparam_declaration1122 specparam_declaration_instance1122();
    specparam_declaration1123 specparam_declaration_instance1123();
    specparam_declaration1124 specparam_declaration_instance1124();
    specparam_declaration1125 specparam_declaration_instance1125();
    specparam_declaration1126 specparam_declaration_instance1126();
    specparam_declaration1127 specparam_declaration_instance1127();
    specparam_declaration1128 specparam_declaration_instance1128();
    specparam_declaration1129 specparam_declaration_instance1129();
    specparam_declaration1130 specparam_declaration_instance1130();
    specparam_declaration1131 specparam_declaration_instance1131();
    specparam_declaration1132 specparam_declaration_instance1132();
    specparam_declaration1133 specparam_declaration_instance1133();
    specparam_declaration1134 specparam_declaration_instance1134();
    specparam_declaration1135 specparam_declaration_instance1135();
    specparam_declaration1136 specparam_declaration_instance1136();
    specparam_declaration1137 specparam_declaration_instance1137();
    specparam_declaration1138 specparam_declaration_instance1138();
    specparam_declaration1139 specparam_declaration_instance1139();
    specparam_declaration1140 specparam_declaration_instance1140();
    specparam_declaration1141 specparam_declaration_instance1141();
    specparam_declaration1142 specparam_declaration_instance1142();
    specparam_declaration1143 specparam_declaration_instance1143();
    specparam_declaration1144 specparam_declaration_instance1144();
    specparam_declaration1145 specparam_declaration_instance1145();
    specparam_declaration1146 specparam_declaration_instance1146();
    specparam_declaration1147 specparam_declaration_instance1147();
    specparam_declaration1148 specparam_declaration_instance1148();
    specparam_declaration1149 specparam_declaration_instance1149();
    specparam_declaration1150 specparam_declaration_instance1150();
    specparam_declaration1151 specparam_declaration_instance1151();
    specparam_declaration1152 specparam_declaration_instance1152();
    specparam_declaration1153 specparam_declaration_instance1153();
    specparam_declaration1154 specparam_declaration_instance1154();
    specparam_declaration1155 specparam_declaration_instance1155();
    specparam_declaration1156 specparam_declaration_instance1156();
    specparam_declaration1157 specparam_declaration_instance1157();
    specparam_declaration1158 specparam_declaration_instance1158();
    specparam_declaration1159 specparam_declaration_instance1159();
    specparam_declaration1160 specparam_declaration_instance1160();
    specparam_declaration1161 specparam_declaration_instance1161();
    specparam_declaration1162 specparam_declaration_instance1162();
    specparam_declaration1163 specparam_declaration_instance1163();
    specparam_declaration1164 specparam_declaration_instance1164();
    specparam_declaration1165 specparam_declaration_instance1165();
    specparam_declaration1166 specparam_declaration_instance1166();
    specparam_declaration1167 specparam_declaration_instance1167();
    specparam_declaration1168 specparam_declaration_instance1168();
    specparam_declaration1169 specparam_declaration_instance1169();
    specparam_declaration1170 specparam_declaration_instance1170();
    specparam_declaration1171 specparam_declaration_instance1171();
    specparam_declaration1172 specparam_declaration_instance1172();
    specparam_declaration1173 specparam_declaration_instance1173();
    specparam_declaration1174 specparam_declaration_instance1174();
    specparam_declaration1175 specparam_declaration_instance1175();
    specparam_declaration1176 specparam_declaration_instance1176();
    specparam_declaration1177 specparam_declaration_instance1177();
    specparam_declaration1178 specparam_declaration_instance1178();
    specparam_declaration1179 specparam_declaration_instance1179();
    specparam_declaration1180 specparam_declaration_instance1180();
    specparam_declaration1181 specparam_declaration_instance1181();
    specparam_declaration1182 specparam_declaration_instance1182();
    specparam_declaration1183 specparam_declaration_instance1183();
    specparam_declaration1184 specparam_declaration_instance1184();
    specparam_declaration1185 specparam_declaration_instance1185();
    specparam_declaration1186 specparam_declaration_instance1186();
    specparam_declaration1187 specparam_declaration_instance1187();
    specparam_declaration1188 specparam_declaration_instance1188();
    specparam_declaration1189 specparam_declaration_instance1189();
    specparam_declaration1190 specparam_declaration_instance1190();
    specparam_declaration1191 specparam_declaration_instance1191();
    specparam_declaration1192 specparam_declaration_instance1192();
    specparam_declaration1193 specparam_declaration_instance1193();
    specparam_declaration1194 specparam_declaration_instance1194();
    specparam_declaration1195 specparam_declaration_instance1195();
    specparam_declaration1196 specparam_declaration_instance1196();
    specparam_declaration1197 specparam_declaration_instance1197();
    specparam_declaration1198 specparam_declaration_instance1198();
    specparam_declaration1199 specparam_declaration_instance1199();
    specparam_declaration1200 specparam_declaration_instance1200();
    specparam_declaration1201 specparam_declaration_instance1201();
    specparam_declaration1202 specparam_declaration_instance1202();
    specparam_declaration1203 specparam_declaration_instance1203();
    specparam_declaration1204 specparam_declaration_instance1204();
    specparam_declaration1205 specparam_declaration_instance1205();
    specparam_declaration1206 specparam_declaration_instance1206();
    specparam_declaration1207 specparam_declaration_instance1207();
    specparam_declaration1208 specparam_declaration_instance1208();
    specparam_declaration1209 specparam_declaration_instance1209();
    specparam_declaration1210 specparam_declaration_instance1210();
    specparam_declaration1211 specparam_declaration_instance1211();
    specparam_declaration1212 specparam_declaration_instance1212();
    specparam_declaration1213 specparam_declaration_instance1213();
    specparam_declaration1214 specparam_declaration_instance1214();
    specparam_declaration1215 specparam_declaration_instance1215();
    specparam_declaration1216 specparam_declaration_instance1216();
    specparam_declaration1217 specparam_declaration_instance1217();
    specparam_declaration1218 specparam_declaration_instance1218();
    specparam_declaration1219 specparam_declaration_instance1219();
    specparam_declaration1220 specparam_declaration_instance1220();
    specparam_declaration1221 specparam_declaration_instance1221();
    specparam_declaration1222 specparam_declaration_instance1222();
    specparam_declaration1223 specparam_declaration_instance1223();
    specparam_declaration1224 specparam_declaration_instance1224();
    specparam_declaration1225 specparam_declaration_instance1225();
    specparam_declaration1226 specparam_declaration_instance1226();
    specparam_declaration1227 specparam_declaration_instance1227();
    specparam_declaration1228 specparam_declaration_instance1228();
    specparam_declaration1229 specparam_declaration_instance1229();
    specparam_declaration1230 specparam_declaration_instance1230();
    specparam_declaration1231 specparam_declaration_instance1231();
    specparam_declaration1232 specparam_declaration_instance1232();
    specparam_declaration1233 specparam_declaration_instance1233();
    specparam_declaration1234 specparam_declaration_instance1234();
    specparam_declaration1235 specparam_declaration_instance1235();
    specparam_declaration1236 specparam_declaration_instance1236();
    specparam_declaration1237 specparam_declaration_instance1237();
    specparam_declaration1238 specparam_declaration_instance1238();
    specparam_declaration1239 specparam_declaration_instance1239();
    specparam_declaration1240 specparam_declaration_instance1240();
    specparam_declaration1241 specparam_declaration_instance1241();
    specparam_declaration1242 specparam_declaration_instance1242();
    specparam_declaration1243 specparam_declaration_instance1243();
    specparam_declaration1244 specparam_declaration_instance1244();
    specparam_declaration1245 specparam_declaration_instance1245();
    specparam_declaration1246 specparam_declaration_instance1246();
    specparam_declaration1247 specparam_declaration_instance1247();
    specparam_declaration1248 specparam_declaration_instance1248();
    specparam_declaration1249 specparam_declaration_instance1249();
    specparam_declaration1250 specparam_declaration_instance1250();
    specparam_declaration1251 specparam_declaration_instance1251();
    specparam_declaration1252 specparam_declaration_instance1252();
    specparam_declaration1253 specparam_declaration_instance1253();
    specparam_declaration1254 specparam_declaration_instance1254();
    specparam_declaration1255 specparam_declaration_instance1255();
    specparam_declaration1256 specparam_declaration_instance1256();
    specparam_declaration1257 specparam_declaration_instance1257();
    specparam_declaration1258 specparam_declaration_instance1258();
    specparam_declaration1259 specparam_declaration_instance1259();
    specparam_declaration1260 specparam_declaration_instance1260();
    specparam_declaration1261 specparam_declaration_instance1261();
    specparam_declaration1262 specparam_declaration_instance1262();
    specparam_declaration1263 specparam_declaration_instance1263();
    specparam_declaration1264 specparam_declaration_instance1264();
    specparam_declaration1265 specparam_declaration_instance1265();
    specparam_declaration1266 specparam_declaration_instance1266();
    specparam_declaration1267 specparam_declaration_instance1267();
    specparam_declaration1268 specparam_declaration_instance1268();
    specparam_declaration1269 specparam_declaration_instance1269();
    specparam_declaration1270 specparam_declaration_instance1270();
    specparam_declaration1271 specparam_declaration_instance1271();
    specparam_declaration1272 specparam_declaration_instance1272();
    specparam_declaration1273 specparam_declaration_instance1273();
    specparam_declaration1274 specparam_declaration_instance1274();
    specparam_declaration1275 specparam_declaration_instance1275();
    specparam_declaration1276 specparam_declaration_instance1276();
    specparam_declaration1277 specparam_declaration_instance1277();
    specparam_declaration1278 specparam_declaration_instance1278();
    specparam_declaration1279 specparam_declaration_instance1279();
    specparam_declaration1280 specparam_declaration_instance1280();
    specparam_declaration1281 specparam_declaration_instance1281();
    specparam_declaration1282 specparam_declaration_instance1282();
    specparam_declaration1283 specparam_declaration_instance1283();
    specparam_declaration1284 specparam_declaration_instance1284();
    specparam_declaration1285 specparam_declaration_instance1285();
    specparam_declaration1286 specparam_declaration_instance1286();
    specparam_declaration1287 specparam_declaration_instance1287();
    specparam_declaration1288 specparam_declaration_instance1288();
    specparam_declaration1289 specparam_declaration_instance1289();
    specparam_declaration1290 specparam_declaration_instance1290();
    specparam_declaration1291 specparam_declaration_instance1291();
    specparam_declaration1292 specparam_declaration_instance1292();
    specparam_declaration1293 specparam_declaration_instance1293();
    specparam_declaration1294 specparam_declaration_instance1294();
    specparam_declaration1295 specparam_declaration_instance1295();
    specparam_declaration1296 specparam_declaration_instance1296();
    specparam_declaration1297 specparam_declaration_instance1297();
    specparam_declaration1298 specparam_declaration_instance1298();
    specparam_declaration1299 specparam_declaration_instance1299();
    specparam_declaration1300 specparam_declaration_instance1300();
    specparam_declaration1301 specparam_declaration_instance1301();
    specparam_declaration1302 specparam_declaration_instance1302();
    specparam_declaration1303 specparam_declaration_instance1303();
    specparam_declaration1304 specparam_declaration_instance1304();
    specparam_declaration1305 specparam_declaration_instance1305();
    specparam_declaration1306 specparam_declaration_instance1306();
    specparam_declaration1307 specparam_declaration_instance1307();
    specparam_declaration1308 specparam_declaration_instance1308();
    specparam_declaration1309 specparam_declaration_instance1309();
    specparam_declaration1310 specparam_declaration_instance1310();
    specparam_declaration1311 specparam_declaration_instance1311();
    specparam_declaration1312 specparam_declaration_instance1312();
    specparam_declaration1313 specparam_declaration_instance1313();
    specparam_declaration1314 specparam_declaration_instance1314();
    specparam_declaration1315 specparam_declaration_instance1315();
    specparam_declaration1316 specparam_declaration_instance1316();
    specparam_declaration1317 specparam_declaration_instance1317();
    specparam_declaration1318 specparam_declaration_instance1318();
    specparam_declaration1319 specparam_declaration_instance1319();
    specparam_declaration1320 specparam_declaration_instance1320();
    specparam_declaration1321 specparam_declaration_instance1321();
    specparam_declaration1322 specparam_declaration_instance1322();
    specparam_declaration1323 specparam_declaration_instance1323();
    specparam_declaration1324 specparam_declaration_instance1324();
    specparam_declaration1325 specparam_declaration_instance1325();
    specparam_declaration1326 specparam_declaration_instance1326();
    specparam_declaration1327 specparam_declaration_instance1327();
    specparam_declaration1328 specparam_declaration_instance1328();
    specparam_declaration1329 specparam_declaration_instance1329();
    specparam_declaration1330 specparam_declaration_instance1330();
    specparam_declaration1331 specparam_declaration_instance1331();
    specparam_declaration1332 specparam_declaration_instance1332();
    specparam_declaration1333 specparam_declaration_instance1333();
    specparam_declaration1334 specparam_declaration_instance1334();
    specparam_declaration1335 specparam_declaration_instance1335();
    specparam_declaration1336 specparam_declaration_instance1336();
    specparam_declaration1337 specparam_declaration_instance1337();
    specparam_declaration1338 specparam_declaration_instance1338();
    specparam_declaration1339 specparam_declaration_instance1339();
    specparam_declaration1340 specparam_declaration_instance1340();
    specparam_declaration1341 specparam_declaration_instance1341();
    specparam_declaration1342 specparam_declaration_instance1342();
    specparam_declaration1343 specparam_declaration_instance1343();
    specparam_declaration1344 specparam_declaration_instance1344();
    specparam_declaration1345 specparam_declaration_instance1345();
    specparam_declaration1346 specparam_declaration_instance1346();
    specparam_declaration1347 specparam_declaration_instance1347();
    specparam_declaration1348 specparam_declaration_instance1348();
    specparam_declaration1349 specparam_declaration_instance1349();
    specparam_declaration1350 specparam_declaration_instance1350();
    specparam_declaration1351 specparam_declaration_instance1351();
    specparam_declaration1352 specparam_declaration_instance1352();
    specparam_declaration1353 specparam_declaration_instance1353();
    specparam_declaration1354 specparam_declaration_instance1354();
    specparam_declaration1355 specparam_declaration_instance1355();
    specparam_declaration1356 specparam_declaration_instance1356();
    specparam_declaration1357 specparam_declaration_instance1357();
    specparam_declaration1358 specparam_declaration_instance1358();
    specparam_declaration1359 specparam_declaration_instance1359();
    specparam_declaration1360 specparam_declaration_instance1360();
    specparam_declaration1361 specparam_declaration_instance1361();
    specparam_declaration1362 specparam_declaration_instance1362();
    specparam_declaration1363 specparam_declaration_instance1363();
    specparam_declaration1364 specparam_declaration_instance1364();
    specparam_declaration1365 specparam_declaration_instance1365();
    specparam_declaration1366 specparam_declaration_instance1366();
    specparam_declaration1367 specparam_declaration_instance1367();
    specparam_declaration1368 specparam_declaration_instance1368();
    specparam_declaration1369 specparam_declaration_instance1369();
    specparam_declaration1370 specparam_declaration_instance1370();
    specparam_declaration1371 specparam_declaration_instance1371();
    specparam_declaration1372 specparam_declaration_instance1372();
    specparam_declaration1373 specparam_declaration_instance1373();
    specparam_declaration1374 specparam_declaration_instance1374();
    specparam_declaration1375 specparam_declaration_instance1375();
    specparam_declaration1376 specparam_declaration_instance1376();
    specparam_declaration1377 specparam_declaration_instance1377();
    specparam_declaration1378 specparam_declaration_instance1378();
    specparam_declaration1379 specparam_declaration_instance1379();
    specparam_declaration1380 specparam_declaration_instance1380();
    specparam_declaration1381 specparam_declaration_instance1381();
    specparam_declaration1382 specparam_declaration_instance1382();
    specparam_declaration1383 specparam_declaration_instance1383();
    specparam_declaration1384 specparam_declaration_instance1384();
    specparam_declaration1385 specparam_declaration_instance1385();
    specparam_declaration1386 specparam_declaration_instance1386();
    specparam_declaration1387 specparam_declaration_instance1387();
    specparam_declaration1388 specparam_declaration_instance1388();
    specparam_declaration1389 specparam_declaration_instance1389();
    specparam_declaration1390 specparam_declaration_instance1390();
    specparam_declaration1391 specparam_declaration_instance1391();
    specparam_declaration1392 specparam_declaration_instance1392();
    specparam_declaration1393 specparam_declaration_instance1393();
    specparam_declaration1394 specparam_declaration_instance1394();
    specparam_declaration1395 specparam_declaration_instance1395();
    specparam_declaration1396 specparam_declaration_instance1396();
    specparam_declaration1397 specparam_declaration_instance1397();
    specparam_declaration1398 specparam_declaration_instance1398();
    specparam_declaration1399 specparam_declaration_instance1399();
    specparam_declaration1400 specparam_declaration_instance1400();
    specparam_declaration1401 specparam_declaration_instance1401();
    specparam_declaration1402 specparam_declaration_instance1402();
    specparam_declaration1403 specparam_declaration_instance1403();
    specparam_declaration1404 specparam_declaration_instance1404();
    specparam_declaration1405 specparam_declaration_instance1405();
    specparam_declaration1406 specparam_declaration_instance1406();
    specparam_declaration1407 specparam_declaration_instance1407();
    specparam_declaration1408 specparam_declaration_instance1408();
    specparam_declaration1409 specparam_declaration_instance1409();
    specparam_declaration1410 specparam_declaration_instance1410();
    specparam_declaration1411 specparam_declaration_instance1411();
    specparam_declaration1412 specparam_declaration_instance1412();
    specparam_declaration1413 specparam_declaration_instance1413();
    specparam_declaration1414 specparam_declaration_instance1414();
    specparam_declaration1415 specparam_declaration_instance1415();
    specparam_declaration1416 specparam_declaration_instance1416();
    specparam_declaration1417 specparam_declaration_instance1417();
    specparam_declaration1418 specparam_declaration_instance1418();
    specparam_declaration1419 specparam_declaration_instance1419();
    specparam_declaration1420 specparam_declaration_instance1420();
    specparam_declaration1421 specparam_declaration_instance1421();
    specparam_declaration1422 specparam_declaration_instance1422();
    specparam_declaration1423 specparam_declaration_instance1423();
    specparam_declaration1424 specparam_declaration_instance1424();
    specparam_declaration1425 specparam_declaration_instance1425();
    specparam_declaration1426 specparam_declaration_instance1426();
    specparam_declaration1427 specparam_declaration_instance1427();
    specparam_declaration1428 specparam_declaration_instance1428();
    specparam_declaration1429 specparam_declaration_instance1429();
    specparam_declaration1430 specparam_declaration_instance1430();
    specparam_declaration1431 specparam_declaration_instance1431();
    specparam_declaration1432 specparam_declaration_instance1432();
    specparam_declaration1433 specparam_declaration_instance1433();
    specparam_declaration1434 specparam_declaration_instance1434();
    specparam_declaration1435 specparam_declaration_instance1435();
    specparam_declaration1436 specparam_declaration_instance1436();
    specparam_declaration1437 specparam_declaration_instance1437();
    specparam_declaration1438 specparam_declaration_instance1438();
    specparam_declaration1439 specparam_declaration_instance1439();
    specparam_declaration1440 specparam_declaration_instance1440();
    specparam_declaration1441 specparam_declaration_instance1441();
    specparam_declaration1442 specparam_declaration_instance1442();
    specparam_declaration1443 specparam_declaration_instance1443();
    specparam_declaration1444 specparam_declaration_instance1444();
    specparam_declaration1445 specparam_declaration_instance1445();
    specparam_declaration1446 specparam_declaration_instance1446();
    specparam_declaration1447 specparam_declaration_instance1447();
    specparam_declaration1448 specparam_declaration_instance1448();
    specparam_declaration1449 specparam_declaration_instance1449();
    specparam_declaration1450 specparam_declaration_instance1450();
    specparam_declaration1451 specparam_declaration_instance1451();
    specparam_declaration1452 specparam_declaration_instance1452();
    specparam_declaration1453 specparam_declaration_instance1453();
    specparam_declaration1454 specparam_declaration_instance1454();
    specparam_declaration1455 specparam_declaration_instance1455();
    specparam_declaration1456 specparam_declaration_instance1456();
    specparam_declaration1457 specparam_declaration_instance1457();
    specparam_declaration1458 specparam_declaration_instance1458();
    specparam_declaration1459 specparam_declaration_instance1459();
    specparam_declaration1460 specparam_declaration_instance1460();
    specparam_declaration1461 specparam_declaration_instance1461();
    specparam_declaration1462 specparam_declaration_instance1462();
    specparam_declaration1463 specparam_declaration_instance1463();
    specparam_declaration1464 specparam_declaration_instance1464();
    specparam_declaration1465 specparam_declaration_instance1465();
    specparam_declaration1466 specparam_declaration_instance1466();
    specparam_declaration1467 specparam_declaration_instance1467();
    specparam_declaration1468 specparam_declaration_instance1468();
    specparam_declaration1469 specparam_declaration_instance1469();
    specparam_declaration1470 specparam_declaration_instance1470();
    specparam_declaration1471 specparam_declaration_instance1471();
    specparam_declaration1472 specparam_declaration_instance1472();
    specparam_declaration1473 specparam_declaration_instance1473();
    specparam_declaration1474 specparam_declaration_instance1474();
    specparam_declaration1475 specparam_declaration_instance1475();
    specparam_declaration1476 specparam_declaration_instance1476();
    specparam_declaration1477 specparam_declaration_instance1477();
    specparam_declaration1478 specparam_declaration_instance1478();
    specparam_declaration1479 specparam_declaration_instance1479();
    specparam_declaration1480 specparam_declaration_instance1480();
    specparam_declaration1481 specparam_declaration_instance1481();
    specparam_declaration1482 specparam_declaration_instance1482();
    specparam_declaration1483 specparam_declaration_instance1483();
    specparam_declaration1484 specparam_declaration_instance1484();
    specparam_declaration1485 specparam_declaration_instance1485();
    specparam_declaration1486 specparam_declaration_instance1486();
    specparam_declaration1487 specparam_declaration_instance1487();
    specparam_declaration1488 specparam_declaration_instance1488();
    specparam_declaration1489 specparam_declaration_instance1489();
    specparam_declaration1490 specparam_declaration_instance1490();
    specparam_declaration1491 specparam_declaration_instance1491();
    specparam_declaration1492 specparam_declaration_instance1492();
    specparam_declaration1493 specparam_declaration_instance1493();
    specparam_declaration1494 specparam_declaration_instance1494();
    specparam_declaration1495 specparam_declaration_instance1495();
    specparam_declaration1496 specparam_declaration_instance1496();
    specparam_declaration1497 specparam_declaration_instance1497();
    specparam_declaration1498 specparam_declaration_instance1498();
    specparam_declaration1499 specparam_declaration_instance1499();
    specparam_declaration1500 specparam_declaration_instance1500();
    specparam_declaration1501 specparam_declaration_instance1501();
    specparam_declaration1502 specparam_declaration_instance1502();
    specparam_declaration1503 specparam_declaration_instance1503();
    specparam_declaration1504 specparam_declaration_instance1504();
    specparam_declaration1505 specparam_declaration_instance1505();
    specparam_declaration1506 specparam_declaration_instance1506();
    specparam_declaration1507 specparam_declaration_instance1507();
    specparam_declaration1508 specparam_declaration_instance1508();
    specparam_declaration1509 specparam_declaration_instance1509();
    specparam_declaration1510 specparam_declaration_instance1510();
    specparam_declaration1511 specparam_declaration_instance1511();
    specparam_declaration1512 specparam_declaration_instance1512();
    specparam_declaration1513 specparam_declaration_instance1513();
    specparam_declaration1514 specparam_declaration_instance1514();
    specparam_declaration1515 specparam_declaration_instance1515();
    specparam_declaration1516 specparam_declaration_instance1516();
    specparam_declaration1517 specparam_declaration_instance1517();
    specparam_declaration1518 specparam_declaration_instance1518();
    specparam_declaration1519 specparam_declaration_instance1519();
    specparam_declaration1520 specparam_declaration_instance1520();
    specparam_declaration1521 specparam_declaration_instance1521();
    specparam_declaration1522 specparam_declaration_instance1522();
    specparam_declaration1523 specparam_declaration_instance1523();
    specparam_declaration1524 specparam_declaration_instance1524();
    specparam_declaration1525 specparam_declaration_instance1525();
    specparam_declaration1526 specparam_declaration_instance1526();
    specparam_declaration1527 specparam_declaration_instance1527();
    specparam_declaration1528 specparam_declaration_instance1528();
    specparam_declaration1529 specparam_declaration_instance1529();
    specparam_declaration1530 specparam_declaration_instance1530();
    specparam_declaration1531 specparam_declaration_instance1531();
    specparam_declaration1532 specparam_declaration_instance1532();
    specparam_declaration1533 specparam_declaration_instance1533();
    specparam_declaration1534 specparam_declaration_instance1534();
    specparam_declaration1535 specparam_declaration_instance1535();
    specparam_declaration1536 specparam_declaration_instance1536();
    specparam_declaration1537 specparam_declaration_instance1537();
    specparam_declaration1538 specparam_declaration_instance1538();
    specparam_declaration1539 specparam_declaration_instance1539();
    specparam_declaration1540 specparam_declaration_instance1540();
    specparam_declaration1541 specparam_declaration_instance1541();
    specparam_declaration1542 specparam_declaration_instance1542();
    specparam_declaration1543 specparam_declaration_instance1543();
    specparam_declaration1544 specparam_declaration_instance1544();
    specparam_declaration1545 specparam_declaration_instance1545();
    specparam_declaration1546 specparam_declaration_instance1546();
    specparam_declaration1547 specparam_declaration_instance1547();
    specparam_declaration1548 specparam_declaration_instance1548();
    specparam_declaration1549 specparam_declaration_instance1549();
    specparam_declaration1550 specparam_declaration_instance1550();
    specparam_declaration1551 specparam_declaration_instance1551();
    specparam_declaration1552 specparam_declaration_instance1552();
    specparam_declaration1553 specparam_declaration_instance1553();
    specparam_declaration1554 specparam_declaration_instance1554();
    specparam_declaration1555 specparam_declaration_instance1555();
    specparam_declaration1556 specparam_declaration_instance1556();
    specparam_declaration1557 specparam_declaration_instance1557();
    specparam_declaration1558 specparam_declaration_instance1558();
    specparam_declaration1559 specparam_declaration_instance1559();
    specparam_declaration1560 specparam_declaration_instance1560();
    specparam_declaration1561 specparam_declaration_instance1561();
    specparam_declaration1562 specparam_declaration_instance1562();
    specparam_declaration1563 specparam_declaration_instance1563();
    specparam_declaration1564 specparam_declaration_instance1564();
    specparam_declaration1565 specparam_declaration_instance1565();
    specparam_declaration1566 specparam_declaration_instance1566();
    specparam_declaration1567 specparam_declaration_instance1567();
    specparam_declaration1568 specparam_declaration_instance1568();
    specparam_declaration1569 specparam_declaration_instance1569();
    specparam_declaration1570 specparam_declaration_instance1570();
    specparam_declaration1571 specparam_declaration_instance1571();
    specparam_declaration1572 specparam_declaration_instance1572();
    specparam_declaration1573 specparam_declaration_instance1573();
    specparam_declaration1574 specparam_declaration_instance1574();
    specparam_declaration1575 specparam_declaration_instance1575();
    specparam_declaration1576 specparam_declaration_instance1576();
    specparam_declaration1577 specparam_declaration_instance1577();
    specparam_declaration1578 specparam_declaration_instance1578();
    specparam_declaration1579 specparam_declaration_instance1579();
    specparam_declaration1580 specparam_declaration_instance1580();
    specparam_declaration1581 specparam_declaration_instance1581();
    specparam_declaration1582 specparam_declaration_instance1582();
    specparam_declaration1583 specparam_declaration_instance1583();
    specparam_declaration1584 specparam_declaration_instance1584();
    specparam_declaration1585 specparam_declaration_instance1585();
    specparam_declaration1586 specparam_declaration_instance1586();
    specparam_declaration1587 specparam_declaration_instance1587();
    specparam_declaration1588 specparam_declaration_instance1588();
    specparam_declaration1589 specparam_declaration_instance1589();
    specparam_declaration1590 specparam_declaration_instance1590();
    specparam_declaration1591 specparam_declaration_instance1591();
    specparam_declaration1592 specparam_declaration_instance1592();
    specparam_declaration1593 specparam_declaration_instance1593();
    specparam_declaration1594 specparam_declaration_instance1594();
    specparam_declaration1595 specparam_declaration_instance1595();
    specparam_declaration1596 specparam_declaration_instance1596();
    specparam_declaration1597 specparam_declaration_instance1597();
    specparam_declaration1598 specparam_declaration_instance1598();
    specparam_declaration1599 specparam_declaration_instance1599();
    specparam_declaration1600 specparam_declaration_instance1600();
    specparam_declaration1601 specparam_declaration_instance1601();
    specparam_declaration1602 specparam_declaration_instance1602();
    specparam_declaration1603 specparam_declaration_instance1603();
    specparam_declaration1604 specparam_declaration_instance1604();
    specparam_declaration1605 specparam_declaration_instance1605();
    specparam_declaration1606 specparam_declaration_instance1606();
    specparam_declaration1607 specparam_declaration_instance1607();
    specparam_declaration1608 specparam_declaration_instance1608();
    specparam_declaration1609 specparam_declaration_instance1609();
    specparam_declaration1610 specparam_declaration_instance1610();
    specparam_declaration1611 specparam_declaration_instance1611();
    specparam_declaration1612 specparam_declaration_instance1612();
    specparam_declaration1613 specparam_declaration_instance1613();
    specparam_declaration1614 specparam_declaration_instance1614();
    specparam_declaration1615 specparam_declaration_instance1615();
    specparam_declaration1616 specparam_declaration_instance1616();
    specparam_declaration1617 specparam_declaration_instance1617();
    specparam_declaration1618 specparam_declaration_instance1618();
    specparam_declaration1619 specparam_declaration_instance1619();
    specparam_declaration1620 specparam_declaration_instance1620();
    specparam_declaration1621 specparam_declaration_instance1621();
    specparam_declaration1622 specparam_declaration_instance1622();
    specparam_declaration1623 specparam_declaration_instance1623();
    specparam_declaration1624 specparam_declaration_instance1624();
    specparam_declaration1625 specparam_declaration_instance1625();
    specparam_declaration1626 specparam_declaration_instance1626();
    specparam_declaration1627 specparam_declaration_instance1627();
    specparam_declaration1628 specparam_declaration_instance1628();
    specparam_declaration1629 specparam_declaration_instance1629();
    specparam_declaration1630 specparam_declaration_instance1630();
    specparam_declaration1631 specparam_declaration_instance1631();
    specparam_declaration1632 specparam_declaration_instance1632();
    specparam_declaration1633 specparam_declaration_instance1633();
    specparam_declaration1634 specparam_declaration_instance1634();
    specparam_declaration1635 specparam_declaration_instance1635();
    specparam_declaration1636 specparam_declaration_instance1636();
    specparam_declaration1637 specparam_declaration_instance1637();
    specparam_declaration1638 specparam_declaration_instance1638();
    specparam_declaration1639 specparam_declaration_instance1639();
    specparam_declaration1640 specparam_declaration_instance1640();
    specparam_declaration1641 specparam_declaration_instance1641();
    specparam_declaration1642 specparam_declaration_instance1642();
    specparam_declaration1643 specparam_declaration_instance1643();
    specparam_declaration1644 specparam_declaration_instance1644();
    specparam_declaration1645 specparam_declaration_instance1645();
    specparam_declaration1646 specparam_declaration_instance1646();
    specparam_declaration1647 specparam_declaration_instance1647();
    specparam_declaration1648 specparam_declaration_instance1648();
    specparam_declaration1649 specparam_declaration_instance1649();
    specparam_declaration1650 specparam_declaration_instance1650();
    specparam_declaration1651 specparam_declaration_instance1651();
    specparam_declaration1652 specparam_declaration_instance1652();
    specparam_declaration1653 specparam_declaration_instance1653();
    specparam_declaration1654 specparam_declaration_instance1654();
    specparam_declaration1655 specparam_declaration_instance1655();
    specparam_declaration1656 specparam_declaration_instance1656();
    specparam_declaration1657 specparam_declaration_instance1657();
    specparam_declaration1658 specparam_declaration_instance1658();
    specparam_declaration1659 specparam_declaration_instance1659();
    specparam_declaration1660 specparam_declaration_instance1660();
    specparam_declaration1661 specparam_declaration_instance1661();
    specparam_declaration1662 specparam_declaration_instance1662();
    specparam_declaration1663 specparam_declaration_instance1663();
    specparam_declaration1664 specparam_declaration_instance1664();
    specparam_declaration1665 specparam_declaration_instance1665();
    specparam_declaration1666 specparam_declaration_instance1666();
    specparam_declaration1667 specparam_declaration_instance1667();
    specparam_declaration1668 specparam_declaration_instance1668();
    specparam_declaration1669 specparam_declaration_instance1669();
    specparam_declaration1670 specparam_declaration_instance1670();
    specparam_declaration1671 specparam_declaration_instance1671();
    specparam_declaration1672 specparam_declaration_instance1672();
    specparam_declaration1673 specparam_declaration_instance1673();
    specparam_declaration1674 specparam_declaration_instance1674();
    specparam_declaration1675 specparam_declaration_instance1675();
    specparam_declaration1676 specparam_declaration_instance1676();
    specparam_declaration1677 specparam_declaration_instance1677();
    specparam_declaration1678 specparam_declaration_instance1678();
    specparam_declaration1679 specparam_declaration_instance1679();
    specparam_declaration1680 specparam_declaration_instance1680();
    specparam_declaration1681 specparam_declaration_instance1681();
    specparam_declaration1682 specparam_declaration_instance1682();
    specparam_declaration1683 specparam_declaration_instance1683();
    specparam_declaration1684 specparam_declaration_instance1684();
    specparam_declaration1685 specparam_declaration_instance1685();
    specparam_declaration1686 specparam_declaration_instance1686();
    specparam_declaration1687 specparam_declaration_instance1687();
    specparam_declaration1688 specparam_declaration_instance1688();
    specparam_declaration1689 specparam_declaration_instance1689();
    specparam_declaration1690 specparam_declaration_instance1690();
    specparam_declaration1691 specparam_declaration_instance1691();
    specparam_declaration1692 specparam_declaration_instance1692();
    specparam_declaration1693 specparam_declaration_instance1693();
    specparam_declaration1694 specparam_declaration_instance1694();
    specparam_declaration1695 specparam_declaration_instance1695();
    specparam_declaration1696 specparam_declaration_instance1696();
    specparam_declaration1697 specparam_declaration_instance1697();
    specparam_declaration1698 specparam_declaration_instance1698();
    specparam_declaration1699 specparam_declaration_instance1699();
    specparam_declaration1700 specparam_declaration_instance1700();
    specparam_declaration1701 specparam_declaration_instance1701();
    specparam_declaration1702 specparam_declaration_instance1702();
    specparam_declaration1703 specparam_declaration_instance1703();
    specparam_declaration1704 specparam_declaration_instance1704();
    specparam_declaration1705 specparam_declaration_instance1705();
    specparam_declaration1706 specparam_declaration_instance1706();
    specparam_declaration1707 specparam_declaration_instance1707();
    specparam_declaration1708 specparam_declaration_instance1708();
    specparam_declaration1709 specparam_declaration_instance1709();
    specparam_declaration1710 specparam_declaration_instance1710();
    specparam_declaration1711 specparam_declaration_instance1711();
    specparam_declaration1712 specparam_declaration_instance1712();
    specparam_declaration1713 specparam_declaration_instance1713();
    specparam_declaration1714 specparam_declaration_instance1714();
    specparam_declaration1715 specparam_declaration_instance1715();
    specparam_declaration1716 specparam_declaration_instance1716();
    specparam_declaration1717 specparam_declaration_instance1717();
    specparam_declaration1718 specparam_declaration_instance1718();
    specparam_declaration1719 specparam_declaration_instance1719();
    specparam_declaration1720 specparam_declaration_instance1720();
    specparam_declaration1721 specparam_declaration_instance1721();
    specparam_declaration1722 specparam_declaration_instance1722();
    specparam_declaration1723 specparam_declaration_instance1723();
    specparam_declaration1724 specparam_declaration_instance1724();
    specparam_declaration1725 specparam_declaration_instance1725();
    specparam_declaration1726 specparam_declaration_instance1726();
    specparam_declaration1727 specparam_declaration_instance1727();
    specparam_declaration1728 specparam_declaration_instance1728();
    specparam_declaration1729 specparam_declaration_instance1729();
    specparam_declaration1730 specparam_declaration_instance1730();
    specparam_declaration1731 specparam_declaration_instance1731();
    specparam_declaration1732 specparam_declaration_instance1732();
    specparam_declaration1733 specparam_declaration_instance1733();
    specparam_declaration1734 specparam_declaration_instance1734();
    specparam_declaration1735 specparam_declaration_instance1735();
    specparam_declaration1736 specparam_declaration_instance1736();
    specparam_declaration1737 specparam_declaration_instance1737();
    specparam_declaration1738 specparam_declaration_instance1738();
    specparam_declaration1739 specparam_declaration_instance1739();
    specparam_declaration1740 specparam_declaration_instance1740();
    specparam_declaration1741 specparam_declaration_instance1741();
    specparam_declaration1742 specparam_declaration_instance1742();
    specparam_declaration1743 specparam_declaration_instance1743();
    specparam_declaration1744 specparam_declaration_instance1744();
    specparam_declaration1745 specparam_declaration_instance1745();
    specparam_declaration1746 specparam_declaration_instance1746();
    specparam_declaration1747 specparam_declaration_instance1747();
    specparam_declaration1748 specparam_declaration_instance1748();
    specparam_declaration1749 specparam_declaration_instance1749();
    specparam_declaration1750 specparam_declaration_instance1750();
    specparam_declaration1751 specparam_declaration_instance1751();
    specparam_declaration1752 specparam_declaration_instance1752();
    specparam_declaration1753 specparam_declaration_instance1753();
    specparam_declaration1754 specparam_declaration_instance1754();
    specparam_declaration1755 specparam_declaration_instance1755();
    specparam_declaration1756 specparam_declaration_instance1756();
    specparam_declaration1757 specparam_declaration_instance1757();
    specparam_declaration1758 specparam_declaration_instance1758();
    specparam_declaration1759 specparam_declaration_instance1759();
    specparam_declaration1760 specparam_declaration_instance1760();
    specparam_declaration1761 specparam_declaration_instance1761();
    specparam_declaration1762 specparam_declaration_instance1762();
    specparam_declaration1763 specparam_declaration_instance1763();
    specparam_declaration1764 specparam_declaration_instance1764();
    specparam_declaration1765 specparam_declaration_instance1765();
    specparam_declaration1766 specparam_declaration_instance1766();
    specparam_declaration1767 specparam_declaration_instance1767();
    specparam_declaration1768 specparam_declaration_instance1768();
    specparam_declaration1769 specparam_declaration_instance1769();
    specparam_declaration1770 specparam_declaration_instance1770();
    specparam_declaration1771 specparam_declaration_instance1771();
    specparam_declaration1772 specparam_declaration_instance1772();
    specparam_declaration1773 specparam_declaration_instance1773();
    specparam_declaration1774 specparam_declaration_instance1774();
    specparam_declaration1775 specparam_declaration_instance1775();
    specparam_declaration1776 specparam_declaration_instance1776();
    specparam_declaration1777 specparam_declaration_instance1777();
    specparam_declaration1778 specparam_declaration_instance1778();
    specparam_declaration1779 specparam_declaration_instance1779();
    specparam_declaration1780 specparam_declaration_instance1780();
    specparam_declaration1781 specparam_declaration_instance1781();
    specparam_declaration1782 specparam_declaration_instance1782();
    specparam_declaration1783 specparam_declaration_instance1783();
    specparam_declaration1784 specparam_declaration_instance1784();
    specparam_declaration1785 specparam_declaration_instance1785();
    specparam_declaration1786 specparam_declaration_instance1786();
    specparam_declaration1787 specparam_declaration_instance1787();
    specparam_declaration1788 specparam_declaration_instance1788();
    specparam_declaration1789 specparam_declaration_instance1789();
    specparam_declaration1790 specparam_declaration_instance1790();
    specparam_declaration1791 specparam_declaration_instance1791();
    specparam_declaration1792 specparam_declaration_instance1792();
    specparam_declaration1793 specparam_declaration_instance1793();
    specparam_declaration1794 specparam_declaration_instance1794();
    specparam_declaration1795 specparam_declaration_instance1795();
    specparam_declaration1796 specparam_declaration_instance1796();
    specparam_declaration1797 specparam_declaration_instance1797();
    specparam_declaration1798 specparam_declaration_instance1798();
    specparam_declaration1799 specparam_declaration_instance1799();
    specparam_declaration1800 specparam_declaration_instance1800();
    specparam_declaration1801 specparam_declaration_instance1801();
    specparam_declaration1802 specparam_declaration_instance1802();
    specparam_declaration1803 specparam_declaration_instance1803();
    specparam_declaration1804 specparam_declaration_instance1804();
    specparam_declaration1805 specparam_declaration_instance1805();
    specparam_declaration1806 specparam_declaration_instance1806();
    specparam_declaration1807 specparam_declaration_instance1807();
    specparam_declaration1808 specparam_declaration_instance1808();
    specparam_declaration1809 specparam_declaration_instance1809();
    specparam_declaration1810 specparam_declaration_instance1810();
    specparam_declaration1811 specparam_declaration_instance1811();
    specparam_declaration1812 specparam_declaration_instance1812();
    specparam_declaration1813 specparam_declaration_instance1813();
    specparam_declaration1814 specparam_declaration_instance1814();
    specparam_declaration1815 specparam_declaration_instance1815();
    specparam_declaration1816 specparam_declaration_instance1816();
    specparam_declaration1817 specparam_declaration_instance1817();
    specparam_declaration1818 specparam_declaration_instance1818();
    specparam_declaration1819 specparam_declaration_instance1819();
    specparam_declaration1820 specparam_declaration_instance1820();
    specparam_declaration1821 specparam_declaration_instance1821();
    specparam_declaration1822 specparam_declaration_instance1822();
    specparam_declaration1823 specparam_declaration_instance1823();
    specparam_declaration1824 specparam_declaration_instance1824();
    specparam_declaration1825 specparam_declaration_instance1825();
    specparam_declaration1826 specparam_declaration_instance1826();
    specparam_declaration1827 specparam_declaration_instance1827();
    specparam_declaration1828 specparam_declaration_instance1828();
    specparam_declaration1829 specparam_declaration_instance1829();
    specparam_declaration1830 specparam_declaration_instance1830();
    specparam_declaration1831 specparam_declaration_instance1831();
    specparam_declaration1832 specparam_declaration_instance1832();
    specparam_declaration1833 specparam_declaration_instance1833();
    specparam_declaration1834 specparam_declaration_instance1834();
    specparam_declaration1835 specparam_declaration_instance1835();
    specparam_declaration1836 specparam_declaration_instance1836();
    specparam_declaration1837 specparam_declaration_instance1837();
    specparam_declaration1838 specparam_declaration_instance1838();
    specparam_declaration1839 specparam_declaration_instance1839();
    specparam_declaration1840 specparam_declaration_instance1840();
    specparam_declaration1841 specparam_declaration_instance1841();
    specparam_declaration1842 specparam_declaration_instance1842();
    specparam_declaration1843 specparam_declaration_instance1843();
    specparam_declaration1844 specparam_declaration_instance1844();
    specparam_declaration1845 specparam_declaration_instance1845();
    specparam_declaration1846 specparam_declaration_instance1846();
    specparam_declaration1847 specparam_declaration_instance1847();
    specparam_declaration1848 specparam_declaration_instance1848();
    specparam_declaration1849 specparam_declaration_instance1849();
    specparam_declaration1850 specparam_declaration_instance1850();
    specparam_declaration1851 specparam_declaration_instance1851();
    specparam_declaration1852 specparam_declaration_instance1852();
    specparam_declaration1853 specparam_declaration_instance1853();
    specparam_declaration1854 specparam_declaration_instance1854();
    specparam_declaration1855 specparam_declaration_instance1855();
    specparam_declaration1856 specparam_declaration_instance1856();
    specparam_declaration1857 specparam_declaration_instance1857();
    specparam_declaration1858 specparam_declaration_instance1858();
    specparam_declaration1859 specparam_declaration_instance1859();
    specparam_declaration1860 specparam_declaration_instance1860();
    specparam_declaration1861 specparam_declaration_instance1861();
    specparam_declaration1862 specparam_declaration_instance1862();
    specparam_declaration1863 specparam_declaration_instance1863();
    specparam_declaration1864 specparam_declaration_instance1864();
    specparam_declaration1865 specparam_declaration_instance1865();
    specparam_declaration1866 specparam_declaration_instance1866();
    specparam_declaration1867 specparam_declaration_instance1867();
    specparam_declaration1868 specparam_declaration_instance1868();
    specparam_declaration1869 specparam_declaration_instance1869();
    specparam_declaration1870 specparam_declaration_instance1870();
    specparam_declaration1871 specparam_declaration_instance1871();
    specparam_declaration1872 specparam_declaration_instance1872();
    specparam_declaration1873 specparam_declaration_instance1873();
    specparam_declaration1874 specparam_declaration_instance1874();
    specparam_declaration1875 specparam_declaration_instance1875();
    specparam_declaration1876 specparam_declaration_instance1876();
    specparam_declaration1877 specparam_declaration_instance1877();
    specparam_declaration1878 specparam_declaration_instance1878();
    specparam_declaration1879 specparam_declaration_instance1879();
    specparam_declaration1880 specparam_declaration_instance1880();
    specparam_declaration1881 specparam_declaration_instance1881();
    specparam_declaration1882 specparam_declaration_instance1882();
    specparam_declaration1883 specparam_declaration_instance1883();
    specparam_declaration1884 specparam_declaration_instance1884();
    specparam_declaration1885 specparam_declaration_instance1885();
    specparam_declaration1886 specparam_declaration_instance1886();
    specparam_declaration1887 specparam_declaration_instance1887();
    specparam_declaration1888 specparam_declaration_instance1888();
    specparam_declaration1889 specparam_declaration_instance1889();
    specparam_declaration1890 specparam_declaration_instance1890();
    specparam_declaration1891 specparam_declaration_instance1891();
    specparam_declaration1892 specparam_declaration_instance1892();
    specparam_declaration1893 specparam_declaration_instance1893();
    specparam_declaration1894 specparam_declaration_instance1894();
    specparam_declaration1895 specparam_declaration_instance1895();
    specparam_declaration1896 specparam_declaration_instance1896();
    specparam_declaration1897 specparam_declaration_instance1897();
    specparam_declaration1898 specparam_declaration_instance1898();
    specparam_declaration1899 specparam_declaration_instance1899();
    specparam_declaration1900 specparam_declaration_instance1900();
    specparam_declaration1901 specparam_declaration_instance1901();
    specparam_declaration1902 specparam_declaration_instance1902();
    specparam_declaration1903 specparam_declaration_instance1903();
    specparam_declaration1904 specparam_declaration_instance1904();
    specparam_declaration1905 specparam_declaration_instance1905();
    specparam_declaration1906 specparam_declaration_instance1906();
    specparam_declaration1907 specparam_declaration_instance1907();
    specparam_declaration1908 specparam_declaration_instance1908();
    specparam_declaration1909 specparam_declaration_instance1909();
    specparam_declaration1910 specparam_declaration_instance1910();
    specparam_declaration1911 specparam_declaration_instance1911();
    specparam_declaration1912 specparam_declaration_instance1912();
    specparam_declaration1913 specparam_declaration_instance1913();
    specparam_declaration1914 specparam_declaration_instance1914();
    specparam_declaration1915 specparam_declaration_instance1915();
    specparam_declaration1916 specparam_declaration_instance1916();
    specparam_declaration1917 specparam_declaration_instance1917();
    specparam_declaration1918 specparam_declaration_instance1918();
    specparam_declaration1919 specparam_declaration_instance1919();
    specparam_declaration1920 specparam_declaration_instance1920();
    specparam_declaration1921 specparam_declaration_instance1921();
    specparam_declaration1922 specparam_declaration_instance1922();
    specparam_declaration1923 specparam_declaration_instance1923();
    specparam_declaration1924 specparam_declaration_instance1924();
    specparam_declaration1925 specparam_declaration_instance1925();
    specparam_declaration1926 specparam_declaration_instance1926();
    specparam_declaration1927 specparam_declaration_instance1927();
    specparam_declaration1928 specparam_declaration_instance1928();
    specparam_declaration1929 specparam_declaration_instance1929();
    specparam_declaration1930 specparam_declaration_instance1930();
    specparam_declaration1931 specparam_declaration_instance1931();
    specparam_declaration1932 specparam_declaration_instance1932();
    specparam_declaration1933 specparam_declaration_instance1933();
    specparam_declaration1934 specparam_declaration_instance1934();
    specparam_declaration1935 specparam_declaration_instance1935();
    specparam_declaration1936 specparam_declaration_instance1936();
    specparam_declaration1937 specparam_declaration_instance1937();
    specparam_declaration1938 specparam_declaration_instance1938();
    specparam_declaration1939 specparam_declaration_instance1939();
    specparam_declaration1940 specparam_declaration_instance1940();
    specparam_declaration1941 specparam_declaration_instance1941();
    specparam_declaration1942 specparam_declaration_instance1942();
    specparam_declaration1943 specparam_declaration_instance1943();
    specparam_declaration1944 specparam_declaration_instance1944();
    specparam_declaration1945 specparam_declaration_instance1945();
    specparam_declaration1946 specparam_declaration_instance1946();
    specparam_declaration1947 specparam_declaration_instance1947();
    specparam_declaration1948 specparam_declaration_instance1948();
    specparam_declaration1949 specparam_declaration_instance1949();
    specparam_declaration1950 specparam_declaration_instance1950();
    specparam_declaration1951 specparam_declaration_instance1951();
    specparam_declaration1952 specparam_declaration_instance1952();
    specparam_declaration1953 specparam_declaration_instance1953();
    specparam_declaration1954 specparam_declaration_instance1954();
    specparam_declaration1955 specparam_declaration_instance1955();
    specparam_declaration1956 specparam_declaration_instance1956();
    specparam_declaration1957 specparam_declaration_instance1957();
    specparam_declaration1958 specparam_declaration_instance1958();
    specparam_declaration1959 specparam_declaration_instance1959();
    specparam_declaration1960 specparam_declaration_instance1960();
    specparam_declaration1961 specparam_declaration_instance1961();
    specparam_declaration1962 specparam_declaration_instance1962();
    specparam_declaration1963 specparam_declaration_instance1963();
    specparam_declaration1964 specparam_declaration_instance1964();
    specparam_declaration1965 specparam_declaration_instance1965();
    specparam_declaration1966 specparam_declaration_instance1966();
    specparam_declaration1967 specparam_declaration_instance1967();
    specparam_declaration1968 specparam_declaration_instance1968();
    specparam_declaration1969 specparam_declaration_instance1969();
    specparam_declaration1970 specparam_declaration_instance1970();
    specparam_declaration1971 specparam_declaration_instance1971();
    specparam_declaration1972 specparam_declaration_instance1972();
    specparam_declaration1973 specparam_declaration_instance1973();
    specparam_declaration1974 specparam_declaration_instance1974();
    specparam_declaration1975 specparam_declaration_instance1975();
    specparam_declaration1976 specparam_declaration_instance1976();
    specparam_declaration1977 specparam_declaration_instance1977();
    specparam_declaration1978 specparam_declaration_instance1978();
    specparam_declaration1979 specparam_declaration_instance1979();
    specparam_declaration1980 specparam_declaration_instance1980();
    specparam_declaration1981 specparam_declaration_instance1981();
    specparam_declaration1982 specparam_declaration_instance1982();
    specparam_declaration1983 specparam_declaration_instance1983();
    specparam_declaration1984 specparam_declaration_instance1984();
    specparam_declaration1985 specparam_declaration_instance1985();
    specparam_declaration1986 specparam_declaration_instance1986();
    specparam_declaration1987 specparam_declaration_instance1987();
    specparam_declaration1988 specparam_declaration_instance1988();
    specparam_declaration1989 specparam_declaration_instance1989();
    specparam_declaration1990 specparam_declaration_instance1990();
    specparam_declaration1991 specparam_declaration_instance1991();
    specparam_declaration1992 specparam_declaration_instance1992();
    specparam_declaration1993 specparam_declaration_instance1993();
    specparam_declaration1994 specparam_declaration_instance1994();
    specparam_declaration1995 specparam_declaration_instance1995();
    specparam_declaration1996 specparam_declaration_instance1996();
    specparam_declaration1997 specparam_declaration_instance1997();
    specparam_declaration1998 specparam_declaration_instance1998();
    specparam_declaration1999 specparam_declaration_instance1999();
    specparam_declaration2000 specparam_declaration_instance2000();
    specparam_declaration2001 specparam_declaration_instance2001();
    specparam_declaration2002 specparam_declaration_instance2002();
    specparam_declaration2003 specparam_declaration_instance2003();
    specparam_declaration2004 specparam_declaration_instance2004();
    specparam_declaration2005 specparam_declaration_instance2005();
    specparam_declaration2006 specparam_declaration_instance2006();
    specparam_declaration2007 specparam_declaration_instance2007();
    specparam_declaration2008 specparam_declaration_instance2008();
    specparam_declaration2009 specparam_declaration_instance2009();
    specparam_declaration2010 specparam_declaration_instance2010();
    specparam_declaration2011 specparam_declaration_instance2011();
    specparam_declaration2012 specparam_declaration_instance2012();
    specparam_declaration2013 specparam_declaration_instance2013();
    specparam_declaration2014 specparam_declaration_instance2014();
    specparam_declaration2015 specparam_declaration_instance2015();
    specparam_declaration2016 specparam_declaration_instance2016();
    specparam_declaration2017 specparam_declaration_instance2017();
    specparam_declaration2018 specparam_declaration_instance2018();
    specparam_declaration2019 specparam_declaration_instance2019();
    specparam_declaration2020 specparam_declaration_instance2020();
    specparam_declaration2021 specparam_declaration_instance2021();
    specparam_declaration2022 specparam_declaration_instance2022();
    specparam_declaration2023 specparam_declaration_instance2023();
    specparam_declaration2024 specparam_declaration_instance2024();
    specparam_declaration2025 specparam_declaration_instance2025();
    specparam_declaration2026 specparam_declaration_instance2026();
    specparam_declaration2027 specparam_declaration_instance2027();
    specparam_declaration2028 specparam_declaration_instance2028();
    specparam_declaration2029 specparam_declaration_instance2029();
    specparam_declaration2030 specparam_declaration_instance2030();
    specparam_declaration2031 specparam_declaration_instance2031();
    specparam_declaration2032 specparam_declaration_instance2032();
    specparam_declaration2033 specparam_declaration_instance2033();
    specparam_declaration2034 specparam_declaration_instance2034();
    specparam_declaration2035 specparam_declaration_instance2035();
    specparam_declaration2036 specparam_declaration_instance2036();
    specparam_declaration2037 specparam_declaration_instance2037();
    specparam_declaration2038 specparam_declaration_instance2038();
    specparam_declaration2039 specparam_declaration_instance2039();
    specparam_declaration2040 specparam_declaration_instance2040();
    specparam_declaration2041 specparam_declaration_instance2041();
    specparam_declaration2042 specparam_declaration_instance2042();
    specparam_declaration2043 specparam_declaration_instance2043();
    specparam_declaration2044 specparam_declaration_instance2044();
    specparam_declaration2045 specparam_declaration_instance2045();
    specparam_declaration2046 specparam_declaration_instance2046();
    specparam_declaration2047 specparam_declaration_instance2047();
    specparam_declaration2048 specparam_declaration_instance2048();
    specparam_declaration2049 specparam_declaration_instance2049();
    specparam_declaration2050 specparam_declaration_instance2050();
    specparam_declaration2051 specparam_declaration_instance2051();
    specparam_declaration2052 specparam_declaration_instance2052();
    specparam_declaration2053 specparam_declaration_instance2053();
    specparam_declaration2054 specparam_declaration_instance2054();
    specparam_declaration2055 specparam_declaration_instance2055();
    specparam_declaration2056 specparam_declaration_instance2056();
    specparam_declaration2057 specparam_declaration_instance2057();
    specparam_declaration2058 specparam_declaration_instance2058();
    specparam_declaration2059 specparam_declaration_instance2059();
    specparam_declaration2060 specparam_declaration_instance2060();
    specparam_declaration2061 specparam_declaration_instance2061();
    specparam_declaration2062 specparam_declaration_instance2062();
    specparam_declaration2063 specparam_declaration_instance2063();
    specparam_declaration2064 specparam_declaration_instance2064();
    specparam_declaration2065 specparam_declaration_instance2065();
    specparam_declaration2066 specparam_declaration_instance2066();
    specparam_declaration2067 specparam_declaration_instance2067();
    specparam_declaration2068 specparam_declaration_instance2068();
    specparam_declaration2069 specparam_declaration_instance2069();
    specparam_declaration2070 specparam_declaration_instance2070();
    specparam_declaration2071 specparam_declaration_instance2071();
    specparam_declaration2072 specparam_declaration_instance2072();
    specparam_declaration2073 specparam_declaration_instance2073();
    specparam_declaration2074 specparam_declaration_instance2074();
    specparam_declaration2075 specparam_declaration_instance2075();
    specparam_declaration2076 specparam_declaration_instance2076();
    specparam_declaration2077 specparam_declaration_instance2077();
    specparam_declaration2078 specparam_declaration_instance2078();
    specparam_declaration2079 specparam_declaration_instance2079();
    specparam_declaration2080 specparam_declaration_instance2080();
    specparam_declaration2081 specparam_declaration_instance2081();
    specparam_declaration2082 specparam_declaration_instance2082();
    specparam_declaration2083 specparam_declaration_instance2083();
    specparam_declaration2084 specparam_declaration_instance2084();
    specparam_declaration2085 specparam_declaration_instance2085();
    specparam_declaration2086 specparam_declaration_instance2086();
    specparam_declaration2087 specparam_declaration_instance2087();
    specparam_declaration2088 specparam_declaration_instance2088();
    specparam_declaration2089 specparam_declaration_instance2089();
    specparam_declaration2090 specparam_declaration_instance2090();
    specparam_declaration2091 specparam_declaration_instance2091();
    specparam_declaration2092 specparam_declaration_instance2092();
    specparam_declaration2093 specparam_declaration_instance2093();
    specparam_declaration2094 specparam_declaration_instance2094();
    specparam_declaration2095 specparam_declaration_instance2095();
    specparam_declaration2096 specparam_declaration_instance2096();
    specparam_declaration2097 specparam_declaration_instance2097();
    specparam_declaration2098 specparam_declaration_instance2098();
    specparam_declaration2099 specparam_declaration_instance2099();
    specparam_declaration2100 specparam_declaration_instance2100();
    specparam_declaration2101 specparam_declaration_instance2101();
    specparam_declaration2102 specparam_declaration_instance2102();
    specparam_declaration2103 specparam_declaration_instance2103();
    specparam_declaration2104 specparam_declaration_instance2104();
    specparam_declaration2105 specparam_declaration_instance2105();
    specparam_declaration2106 specparam_declaration_instance2106();
    specparam_declaration2107 specparam_declaration_instance2107();
    specparam_declaration2108 specparam_declaration_instance2108();
    specparam_declaration2109 specparam_declaration_instance2109();
    specparam_declaration2110 specparam_declaration_instance2110();
    specparam_declaration2111 specparam_declaration_instance2111();
    specparam_declaration2112 specparam_declaration_instance2112();
    specparam_declaration2113 specparam_declaration_instance2113();
    specparam_declaration2114 specparam_declaration_instance2114();
    specparam_declaration2115 specparam_declaration_instance2115();
    specparam_declaration2116 specparam_declaration_instance2116();
    specparam_declaration2117 specparam_declaration_instance2117();
    specparam_declaration2118 specparam_declaration_instance2118();
    specparam_declaration2119 specparam_declaration_instance2119();
    specparam_declaration2120 specparam_declaration_instance2120();
    specparam_declaration2121 specparam_declaration_instance2121();
    specparam_declaration2122 specparam_declaration_instance2122();
    specparam_declaration2123 specparam_declaration_instance2123();
    specparam_declaration2124 specparam_declaration_instance2124();
    specparam_declaration2125 specparam_declaration_instance2125();
    specparam_declaration2126 specparam_declaration_instance2126();
    specparam_declaration2127 specparam_declaration_instance2127();
    specparam_declaration2128 specparam_declaration_instance2128();
    specparam_declaration2129 specparam_declaration_instance2129();
    specparam_declaration2130 specparam_declaration_instance2130();
    specparam_declaration2131 specparam_declaration_instance2131();
    specparam_declaration2132 specparam_declaration_instance2132();
    specparam_declaration2133 specparam_declaration_instance2133();
    specparam_declaration2134 specparam_declaration_instance2134();
    specparam_declaration2135 specparam_declaration_instance2135();
    specparam_declaration2136 specparam_declaration_instance2136();
    specparam_declaration2137 specparam_declaration_instance2137();
    specparam_declaration2138 specparam_declaration_instance2138();
    specparam_declaration2139 specparam_declaration_instance2139();
    specparam_declaration2140 specparam_declaration_instance2140();
    specparam_declaration2141 specparam_declaration_instance2141();
    specparam_declaration2142 specparam_declaration_instance2142();
    specparam_declaration2143 specparam_declaration_instance2143();
    specparam_declaration2144 specparam_declaration_instance2144();
    specparam_declaration2145 specparam_declaration_instance2145();
    specparam_declaration2146 specparam_declaration_instance2146();
    specparam_declaration2147 specparam_declaration_instance2147();
    specparam_declaration2148 specparam_declaration_instance2148();
    specparam_declaration2149 specparam_declaration_instance2149();
    specparam_declaration2150 specparam_declaration_instance2150();
    specparam_declaration2151 specparam_declaration_instance2151();
    specparam_declaration2152 specparam_declaration_instance2152();
    specparam_declaration2153 specparam_declaration_instance2153();
    specparam_declaration2154 specparam_declaration_instance2154();
    specparam_declaration2155 specparam_declaration_instance2155();
    specparam_declaration2156 specparam_declaration_instance2156();
    specparam_declaration2157 specparam_declaration_instance2157();
    specparam_declaration2158 specparam_declaration_instance2158();
    specparam_declaration2159 specparam_declaration_instance2159();
    specparam_declaration2160 specparam_declaration_instance2160();
    specparam_declaration2161 specparam_declaration_instance2161();
    specparam_declaration2162 specparam_declaration_instance2162();
    specparam_declaration2163 specparam_declaration_instance2163();
    specparam_declaration2164 specparam_declaration_instance2164();
    specparam_declaration2165 specparam_declaration_instance2165();
    specparam_declaration2166 specparam_declaration_instance2166();
    specparam_declaration2167 specparam_declaration_instance2167();
    specparam_declaration2168 specparam_declaration_instance2168();
    specparam_declaration2169 specparam_declaration_instance2169();
    specparam_declaration2170 specparam_declaration_instance2170();
    specparam_declaration2171 specparam_declaration_instance2171();
    specparam_declaration2172 specparam_declaration_instance2172();
    specparam_declaration2173 specparam_declaration_instance2173();
    specparam_declaration2174 specparam_declaration_instance2174();
    specparam_declaration2175 specparam_declaration_instance2175();
    specparam_declaration2176 specparam_declaration_instance2176();
    specparam_declaration2177 specparam_declaration_instance2177();
    specparam_declaration2178 specparam_declaration_instance2178();
    specparam_declaration2179 specparam_declaration_instance2179();
    specparam_declaration2180 specparam_declaration_instance2180();
    specparam_declaration2181 specparam_declaration_instance2181();
    specparam_declaration2182 specparam_declaration_instance2182();
    specparam_declaration2183 specparam_declaration_instance2183();
    specparam_declaration2184 specparam_declaration_instance2184();
    specparam_declaration2185 specparam_declaration_instance2185();
    specparam_declaration2186 specparam_declaration_instance2186();
    specparam_declaration2187 specparam_declaration_instance2187();
    specparam_declaration2188 specparam_declaration_instance2188();
    specparam_declaration2189 specparam_declaration_instance2189();
    specparam_declaration2190 specparam_declaration_instance2190();
    specparam_declaration2191 specparam_declaration_instance2191();
    specparam_declaration2192 specparam_declaration_instance2192();
    specparam_declaration2193 specparam_declaration_instance2193();
    specparam_declaration2194 specparam_declaration_instance2194();
    specparam_declaration2195 specparam_declaration_instance2195();
    specparam_declaration2196 specparam_declaration_instance2196();
    specparam_declaration2197 specparam_declaration_instance2197();
    specparam_declaration2198 specparam_declaration_instance2198();
    specparam_declaration2199 specparam_declaration_instance2199();
    specparam_declaration2200 specparam_declaration_instance2200();
    specparam_declaration2201 specparam_declaration_instance2201();
    specparam_declaration2202 specparam_declaration_instance2202();
    specparam_declaration2203 specparam_declaration_instance2203();
    specparam_declaration2204 specparam_declaration_instance2204();
    specparam_declaration2205 specparam_declaration_instance2205();
    specparam_declaration2206 specparam_declaration_instance2206();
    specparam_declaration2207 specparam_declaration_instance2207();
    specparam_declaration2208 specparam_declaration_instance2208();
    specparam_declaration2209 specparam_declaration_instance2209();
    specparam_declaration2210 specparam_declaration_instance2210();
    specparam_declaration2211 specparam_declaration_instance2211();
    specparam_declaration2212 specparam_declaration_instance2212();
    specparam_declaration2213 specparam_declaration_instance2213();
    specparam_declaration2214 specparam_declaration_instance2214();
    specparam_declaration2215 specparam_declaration_instance2215();
    specparam_declaration2216 specparam_declaration_instance2216();
    specparam_declaration2217 specparam_declaration_instance2217();
    specparam_declaration2218 specparam_declaration_instance2218();
    specparam_declaration2219 specparam_declaration_instance2219();
    specparam_declaration2220 specparam_declaration_instance2220();
    specparam_declaration2221 specparam_declaration_instance2221();
    specparam_declaration2222 specparam_declaration_instance2222();
    specparam_declaration2223 specparam_declaration_instance2223();
    specparam_declaration2224 specparam_declaration_instance2224();
    specparam_declaration2225 specparam_declaration_instance2225();
    specparam_declaration2226 specparam_declaration_instance2226();
    specparam_declaration2227 specparam_declaration_instance2227();
    specparam_declaration2228 specparam_declaration_instance2228();
    specparam_declaration2229 specparam_declaration_instance2229();
    specparam_declaration2230 specparam_declaration_instance2230();
    specparam_declaration2231 specparam_declaration_instance2231();
    specparam_declaration2232 specparam_declaration_instance2232();
    specparam_declaration2233 specparam_declaration_instance2233();
    specparam_declaration2234 specparam_declaration_instance2234();
    specparam_declaration2235 specparam_declaration_instance2235();
    specparam_declaration2236 specparam_declaration_instance2236();
    specparam_declaration2237 specparam_declaration_instance2237();
    specparam_declaration2238 specparam_declaration_instance2238();
    specparam_declaration2239 specparam_declaration_instance2239();
    specparam_declaration2240 specparam_declaration_instance2240();
    specparam_declaration2241 specparam_declaration_instance2241();
    specparam_declaration2242 specparam_declaration_instance2242();
    specparam_declaration2243 specparam_declaration_instance2243();
    specparam_declaration2244 specparam_declaration_instance2244();
    specparam_declaration2245 specparam_declaration_instance2245();
    specparam_declaration2246 specparam_declaration_instance2246();
    specparam_declaration2247 specparam_declaration_instance2247();
    specparam_declaration2248 specparam_declaration_instance2248();
    specparam_declaration2249 specparam_declaration_instance2249();
    specparam_declaration2250 specparam_declaration_instance2250();
    specparam_declaration2251 specparam_declaration_instance2251();
    specparam_declaration2252 specparam_declaration_instance2252();
    specparam_declaration2253 specparam_declaration_instance2253();
    specparam_declaration2254 specparam_declaration_instance2254();
    specparam_declaration2255 specparam_declaration_instance2255();
    specparam_declaration2256 specparam_declaration_instance2256();
    specparam_declaration2257 specparam_declaration_instance2257();
    specparam_declaration2258 specparam_declaration_instance2258();
    specparam_declaration2259 specparam_declaration_instance2259();
    specparam_declaration2260 specparam_declaration_instance2260();
    specparam_declaration2261 specparam_declaration_instance2261();
    specparam_declaration2262 specparam_declaration_instance2262();
    specparam_declaration2263 specparam_declaration_instance2263();
    specparam_declaration2264 specparam_declaration_instance2264();
    specparam_declaration2265 specparam_declaration_instance2265();
    specparam_declaration2266 specparam_declaration_instance2266();
    specparam_declaration2267 specparam_declaration_instance2267();
    specparam_declaration2268 specparam_declaration_instance2268();
    specparam_declaration2269 specparam_declaration_instance2269();
    specparam_declaration2270 specparam_declaration_instance2270();
    specparam_declaration2271 specparam_declaration_instance2271();
    specparam_declaration2272 specparam_declaration_instance2272();
    specparam_declaration2273 specparam_declaration_instance2273();
    specparam_declaration2274 specparam_declaration_instance2274();
    specparam_declaration2275 specparam_declaration_instance2275();
    specparam_declaration2276 specparam_declaration_instance2276();
    specparam_declaration2277 specparam_declaration_instance2277();
    specparam_declaration2278 specparam_declaration_instance2278();
    specparam_declaration2279 specparam_declaration_instance2279();
    specparam_declaration2280 specparam_declaration_instance2280();
    specparam_declaration2281 specparam_declaration_instance2281();
    specparam_declaration2282 specparam_declaration_instance2282();
    specparam_declaration2283 specparam_declaration_instance2283();
    specparam_declaration2284 specparam_declaration_instance2284();
    specparam_declaration2285 specparam_declaration_instance2285();
    specparam_declaration2286 specparam_declaration_instance2286();
    specparam_declaration2287 specparam_declaration_instance2287();
    specparam_declaration2288 specparam_declaration_instance2288();
    specparam_declaration2289 specparam_declaration_instance2289();
    specparam_declaration2290 specparam_declaration_instance2290();
    specparam_declaration2291 specparam_declaration_instance2291();
    specparam_declaration2292 specparam_declaration_instance2292();
    specparam_declaration2293 specparam_declaration_instance2293();
    specparam_declaration2294 specparam_declaration_instance2294();
    specparam_declaration2295 specparam_declaration_instance2295();
    specparam_declaration2296 specparam_declaration_instance2296();
    specparam_declaration2297 specparam_declaration_instance2297();
    specparam_declaration2298 specparam_declaration_instance2298();
    specparam_declaration2299 specparam_declaration_instance2299();
    specparam_declaration2300 specparam_declaration_instance2300();
    specparam_declaration2301 specparam_declaration_instance2301();
    specparam_declaration2302 specparam_declaration_instance2302();
    specparam_declaration2303 specparam_declaration_instance2303();
    specparam_declaration2304 specparam_declaration_instance2304();
    specparam_declaration2305 specparam_declaration_instance2305();
    specparam_declaration2306 specparam_declaration_instance2306();
    specparam_declaration2307 specparam_declaration_instance2307();
    specparam_declaration2308 specparam_declaration_instance2308();
    specparam_declaration2309 specparam_declaration_instance2309();
    specparam_declaration2310 specparam_declaration_instance2310();
    specparam_declaration2311 specparam_declaration_instance2311();
    specparam_declaration2312 specparam_declaration_instance2312();
    specparam_declaration2313 specparam_declaration_instance2313();
    specparam_declaration2314 specparam_declaration_instance2314();
    specparam_declaration2315 specparam_declaration_instance2315();
    specparam_declaration2316 specparam_declaration_instance2316();
    specparam_declaration2317 specparam_declaration_instance2317();
    specparam_declaration2318 specparam_declaration_instance2318();
    specparam_declaration2319 specparam_declaration_instance2319();
    specparam_declaration2320 specparam_declaration_instance2320();
    specparam_declaration2321 specparam_declaration_instance2321();
    specparam_declaration2322 specparam_declaration_instance2322();
    specparam_declaration2323 specparam_declaration_instance2323();
    specparam_declaration2324 specparam_declaration_instance2324();
    specparam_declaration2325 specparam_declaration_instance2325();
    specparam_declaration2326 specparam_declaration_instance2326();
    specparam_declaration2327 specparam_declaration_instance2327();
    specparam_declaration2328 specparam_declaration_instance2328();
    specparam_declaration2329 specparam_declaration_instance2329();
    specparam_declaration2330 specparam_declaration_instance2330();
    specparam_declaration2331 specparam_declaration_instance2331();
    specparam_declaration2332 specparam_declaration_instance2332();
    specparam_declaration2333 specparam_declaration_instance2333();
    specparam_declaration2334 specparam_declaration_instance2334();
    specparam_declaration2335 specparam_declaration_instance2335();
    specparam_declaration2336 specparam_declaration_instance2336();
    specparam_declaration2337 specparam_declaration_instance2337();
    specparam_declaration2338 specparam_declaration_instance2338();
    specparam_declaration2339 specparam_declaration_instance2339();
    specparam_declaration2340 specparam_declaration_instance2340();
    specparam_declaration2341 specparam_declaration_instance2341();
    specparam_declaration2342 specparam_declaration_instance2342();
    specparam_declaration2343 specparam_declaration_instance2343();
    specparam_declaration2344 specparam_declaration_instance2344();
    specparam_declaration2345 specparam_declaration_instance2345();
    specparam_declaration2346 specparam_declaration_instance2346();
    specparam_declaration2347 specparam_declaration_instance2347();
    specparam_declaration2348 specparam_declaration_instance2348();
    specparam_declaration2349 specparam_declaration_instance2349();
    specparam_declaration2350 specparam_declaration_instance2350();
    specparam_declaration2351 specparam_declaration_instance2351();
    specparam_declaration2352 specparam_declaration_instance2352();
    specparam_declaration2353 specparam_declaration_instance2353();
    specparam_declaration2354 specparam_declaration_instance2354();
    specparam_declaration2355 specparam_declaration_instance2355();
    specparam_declaration2356 specparam_declaration_instance2356();
    specparam_declaration2357 specparam_declaration_instance2357();
    specparam_declaration2358 specparam_declaration_instance2358();
    specparam_declaration2359 specparam_declaration_instance2359();
    specparam_declaration2360 specparam_declaration_instance2360();
    specparam_declaration2361 specparam_declaration_instance2361();
    specparam_declaration2362 specparam_declaration_instance2362();
    specparam_declaration2363 specparam_declaration_instance2363();
    specparam_declaration2364 specparam_declaration_instance2364();
    specparam_declaration2365 specparam_declaration_instance2365();
    specparam_declaration2366 specparam_declaration_instance2366();
    specparam_declaration2367 specparam_declaration_instance2367();
    specparam_declaration2368 specparam_declaration_instance2368();
    specparam_declaration2369 specparam_declaration_instance2369();
    specparam_declaration2370 specparam_declaration_instance2370();
    specparam_declaration2371 specparam_declaration_instance2371();
    specparam_declaration2372 specparam_declaration_instance2372();
    specparam_declaration2373 specparam_declaration_instance2373();
    specparam_declaration2374 specparam_declaration_instance2374();
    specparam_declaration2375 specparam_declaration_instance2375();
    specparam_declaration2376 specparam_declaration_instance2376();
    specparam_declaration2377 specparam_declaration_instance2377();
    specparam_declaration2378 specparam_declaration_instance2378();
    specparam_declaration2379 specparam_declaration_instance2379();
    specparam_declaration2380 specparam_declaration_instance2380();
    specparam_declaration2381 specparam_declaration_instance2381();
    specparam_declaration2382 specparam_declaration_instance2382();
    specparam_declaration2383 specparam_declaration_instance2383();
    specparam_declaration2384 specparam_declaration_instance2384();
    specparam_declaration2385 specparam_declaration_instance2385();
    specparam_declaration2386 specparam_declaration_instance2386();
    specparam_declaration2387 specparam_declaration_instance2387();
    specparam_declaration2388 specparam_declaration_instance2388();
    specparam_declaration2389 specparam_declaration_instance2389();
    specparam_declaration2390 specparam_declaration_instance2390();
    specparam_declaration2391 specparam_declaration_instance2391();
    specparam_declaration2392 specparam_declaration_instance2392();
    specparam_declaration2393 specparam_declaration_instance2393();
    specparam_declaration2394 specparam_declaration_instance2394();
    specparam_declaration2395 specparam_declaration_instance2395();
    specparam_declaration2396 specparam_declaration_instance2396();
    specparam_declaration2397 specparam_declaration_instance2397();
    specparam_declaration2398 specparam_declaration_instance2398();
    specparam_declaration2399 specparam_declaration_instance2399();
    specparam_declaration2400 specparam_declaration_instance2400();
    specparam_declaration2401 specparam_declaration_instance2401();
    specparam_declaration2402 specparam_declaration_instance2402();
    specparam_declaration2403 specparam_declaration_instance2403();
    specparam_declaration2404 specparam_declaration_instance2404();
    specparam_declaration2405 specparam_declaration_instance2405();
    specparam_declaration2406 specparam_declaration_instance2406();
    specparam_declaration2407 specparam_declaration_instance2407();
    specparam_declaration2408 specparam_declaration_instance2408();
    specparam_declaration2409 specparam_declaration_instance2409();
    specparam_declaration2410 specparam_declaration_instance2410();
    specparam_declaration2411 specparam_declaration_instance2411();
    specparam_declaration2412 specparam_declaration_instance2412();
    specparam_declaration2413 specparam_declaration_instance2413();
    specparam_declaration2414 specparam_declaration_instance2414();
    specparam_declaration2415 specparam_declaration_instance2415();
    specparam_declaration2416 specparam_declaration_instance2416();
    specparam_declaration2417 specparam_declaration_instance2417();
    specparam_declaration2418 specparam_declaration_instance2418();
    specparam_declaration2419 specparam_declaration_instance2419();
    specparam_declaration2420 specparam_declaration_instance2420();
    specparam_declaration2421 specparam_declaration_instance2421();
    specparam_declaration2422 specparam_declaration_instance2422();
    specparam_declaration2423 specparam_declaration_instance2423();
    specparam_declaration2424 specparam_declaration_instance2424();
    specparam_declaration2425 specparam_declaration_instance2425();
    specparam_declaration2426 specparam_declaration_instance2426();
    specparam_declaration2427 specparam_declaration_instance2427();
    specparam_declaration2428 specparam_declaration_instance2428();
    specparam_declaration2429 specparam_declaration_instance2429();
    specparam_declaration2430 specparam_declaration_instance2430();
    specparam_declaration2431 specparam_declaration_instance2431();
    specparam_declaration2432 specparam_declaration_instance2432();
    specparam_declaration2433 specparam_declaration_instance2433();
    specparam_declaration2434 specparam_declaration_instance2434();
    specparam_declaration2435 specparam_declaration_instance2435();
    specparam_declaration2436 specparam_declaration_instance2436();
    specparam_declaration2437 specparam_declaration_instance2437();
    specparam_declaration2438 specparam_declaration_instance2438();
    specparam_declaration2439 specparam_declaration_instance2439();
    specparam_declaration2440 specparam_declaration_instance2440();
    specparam_declaration2441 specparam_declaration_instance2441();
    specparam_declaration2442 specparam_declaration_instance2442();
    specparam_declaration2443 specparam_declaration_instance2443();
    specparam_declaration2444 specparam_declaration_instance2444();
    specparam_declaration2445 specparam_declaration_instance2445();
    specparam_declaration2446 specparam_declaration_instance2446();
    specparam_declaration2447 specparam_declaration_instance2447();
    specparam_declaration2448 specparam_declaration_instance2448();
    specparam_declaration2449 specparam_declaration_instance2449();
    specparam_declaration2450 specparam_declaration_instance2450();
    specparam_declaration2451 specparam_declaration_instance2451();
    specparam_declaration2452 specparam_declaration_instance2452();
    specparam_declaration2453 specparam_declaration_instance2453();
    specparam_declaration2454 specparam_declaration_instance2454();
    specparam_declaration2455 specparam_declaration_instance2455();
    specparam_declaration2456 specparam_declaration_instance2456();
    specparam_declaration2457 specparam_declaration_instance2457();
    specparam_declaration2458 specparam_declaration_instance2458();
    specparam_declaration2459 specparam_declaration_instance2459();
    specparam_declaration2460 specparam_declaration_instance2460();
    specparam_declaration2461 specparam_declaration_instance2461();
    specparam_declaration2462 specparam_declaration_instance2462();
    specparam_declaration2463 specparam_declaration_instance2463();
    specparam_declaration2464 specparam_declaration_instance2464();
    specparam_declaration2465 specparam_declaration_instance2465();
    specparam_declaration2466 specparam_declaration_instance2466();
    specparam_declaration2467 specparam_declaration_instance2467();
    specparam_declaration2468 specparam_declaration_instance2468();
    specparam_declaration2469 specparam_declaration_instance2469();
    specparam_declaration2470 specparam_declaration_instance2470();
    specparam_declaration2471 specparam_declaration_instance2471();
    specparam_declaration2472 specparam_declaration_instance2472();
    specparam_declaration2473 specparam_declaration_instance2473();
    specparam_declaration2474 specparam_declaration_instance2474();
    specparam_declaration2475 specparam_declaration_instance2475();
    specparam_declaration2476 specparam_declaration_instance2476();
    specparam_declaration2477 specparam_declaration_instance2477();
    specparam_declaration2478 specparam_declaration_instance2478();
    specparam_declaration2479 specparam_declaration_instance2479();
    specparam_declaration2480 specparam_declaration_instance2480();
    specparam_declaration2481 specparam_declaration_instance2481();
    specparam_declaration2482 specparam_declaration_instance2482();
    specparam_declaration2483 specparam_declaration_instance2483();
    specparam_declaration2484 specparam_declaration_instance2484();
    specparam_declaration2485 specparam_declaration_instance2485();
    specparam_declaration2486 specparam_declaration_instance2486();
    specparam_declaration2487 specparam_declaration_instance2487();
    specparam_declaration2488 specparam_declaration_instance2488();
    specparam_declaration2489 specparam_declaration_instance2489();
    specparam_declaration2490 specparam_declaration_instance2490();
    specparam_declaration2491 specparam_declaration_instance2491();
    specparam_declaration2492 specparam_declaration_instance2492();
    specparam_declaration2493 specparam_declaration_instance2493();
    specparam_declaration2494 specparam_declaration_instance2494();
    specparam_declaration2495 specparam_declaration_instance2495();
    specparam_declaration2496 specparam_declaration_instance2496();
    specparam_declaration2497 specparam_declaration_instance2497();
    specparam_declaration2498 specparam_declaration_instance2498();
    specparam_declaration2499 specparam_declaration_instance2499();
    specparam_declaration2500 specparam_declaration_instance2500();
    specparam_declaration2501 specparam_declaration_instance2501();
    specparam_declaration2502 specparam_declaration_instance2502();
    specparam_declaration2503 specparam_declaration_instance2503();
    specparam_declaration2504 specparam_declaration_instance2504();
    specparam_declaration2505 specparam_declaration_instance2505();
    specparam_declaration2506 specparam_declaration_instance2506();
    specparam_declaration2507 specparam_declaration_instance2507();
    specparam_declaration2508 specparam_declaration_instance2508();
    specparam_declaration2509 specparam_declaration_instance2509();
    specparam_declaration2510 specparam_declaration_instance2510();
    specparam_declaration2511 specparam_declaration_instance2511();
    specparam_declaration2512 specparam_declaration_instance2512();
    specparam_declaration2513 specparam_declaration_instance2513();
    specparam_declaration2514 specparam_declaration_instance2514();
    specparam_declaration2515 specparam_declaration_instance2515();
    specparam_declaration2516 specparam_declaration_instance2516();
    specparam_declaration2517 specparam_declaration_instance2517();
    specparam_declaration2518 specparam_declaration_instance2518();
    specparam_declaration2519 specparam_declaration_instance2519();
    specparam_declaration2520 specparam_declaration_instance2520();
    specparam_declaration2521 specparam_declaration_instance2521();
    specparam_declaration2522 specparam_declaration_instance2522();
    specparam_declaration2523 specparam_declaration_instance2523();
    specparam_declaration2524 specparam_declaration_instance2524();
    specparam_declaration2525 specparam_declaration_instance2525();
    specparam_declaration2526 specparam_declaration_instance2526();
    specparam_declaration2527 specparam_declaration_instance2527();
    specparam_declaration2528 specparam_declaration_instance2528();
    specparam_declaration2529 specparam_declaration_instance2529();
    specparam_declaration2530 specparam_declaration_instance2530();
    specparam_declaration2531 specparam_declaration_instance2531();
    specparam_declaration2532 specparam_declaration_instance2532();
    specparam_declaration2533 specparam_declaration_instance2533();
    specparam_declaration2534 specparam_declaration_instance2534();
    specparam_declaration2535 specparam_declaration_instance2535();
    specparam_declaration2536 specparam_declaration_instance2536();
    specparam_declaration2537 specparam_declaration_instance2537();
    specparam_declaration2538 specparam_declaration_instance2538();
    specparam_declaration2539 specparam_declaration_instance2539();
    specparam_declaration2540 specparam_declaration_instance2540();
    specparam_declaration2541 specparam_declaration_instance2541();
    specparam_declaration2542 specparam_declaration_instance2542();
    specparam_declaration2543 specparam_declaration_instance2543();
    specparam_declaration2544 specparam_declaration_instance2544();
    specparam_declaration2545 specparam_declaration_instance2545();
    specparam_declaration2546 specparam_declaration_instance2546();
    specparam_declaration2547 specparam_declaration_instance2547();
    specparam_declaration2548 specparam_declaration_instance2548();
    specparam_declaration2549 specparam_declaration_instance2549();
    specparam_declaration2550 specparam_declaration_instance2550();
    specparam_declaration2551 specparam_declaration_instance2551();
    specparam_declaration2552 specparam_declaration_instance2552();
    specparam_declaration2553 specparam_declaration_instance2553();
    specparam_declaration2554 specparam_declaration_instance2554();
    specparam_declaration2555 specparam_declaration_instance2555();
    specparam_declaration2556 specparam_declaration_instance2556();
    specparam_declaration2557 specparam_declaration_instance2557();
    specparam_declaration2558 specparam_declaration_instance2558();
    specparam_declaration2559 specparam_declaration_instance2559();
    specparam_declaration2560 specparam_declaration_instance2560();
    specparam_declaration2561 specparam_declaration_instance2561();
    specparam_declaration2562 specparam_declaration_instance2562();
    specparam_declaration2563 specparam_declaration_instance2563();
    specparam_declaration2564 specparam_declaration_instance2564();
    specparam_declaration2565 specparam_declaration_instance2565();
    specparam_declaration2566 specparam_declaration_instance2566();
    specparam_declaration2567 specparam_declaration_instance2567();
    specparam_declaration2568 specparam_declaration_instance2568();
    specparam_declaration2569 specparam_declaration_instance2569();
    specparam_declaration2570 specparam_declaration_instance2570();
    specparam_declaration2571 specparam_declaration_instance2571();
    specparam_declaration2572 specparam_declaration_instance2572();
    specparam_declaration2573 specparam_declaration_instance2573();
    specparam_declaration2574 specparam_declaration_instance2574();
    specparam_declaration2575 specparam_declaration_instance2575();
    specparam_declaration2576 specparam_declaration_instance2576();
    specparam_declaration2577 specparam_declaration_instance2577();
    specparam_declaration2578 specparam_declaration_instance2578();
    specparam_declaration2579 specparam_declaration_instance2579();
    specparam_declaration2580 specparam_declaration_instance2580();
    specparam_declaration2581 specparam_declaration_instance2581();
    specparam_declaration2582 specparam_declaration_instance2582();
    specparam_declaration2583 specparam_declaration_instance2583();
    specparam_declaration2584 specparam_declaration_instance2584();
    specparam_declaration2585 specparam_declaration_instance2585();
    specparam_declaration2586 specparam_declaration_instance2586();
    specparam_declaration2587 specparam_declaration_instance2587();
    specparam_declaration2588 specparam_declaration_instance2588();
    specparam_declaration2589 specparam_declaration_instance2589();
    specparam_declaration2590 specparam_declaration_instance2590();
    specparam_declaration2591 specparam_declaration_instance2591();
    specparam_declaration2592 specparam_declaration_instance2592();
    specparam_declaration2593 specparam_declaration_instance2593();
    specparam_declaration2594 specparam_declaration_instance2594();
    specparam_declaration2595 specparam_declaration_instance2595();
    specparam_declaration2596 specparam_declaration_instance2596();
    specparam_declaration2597 specparam_declaration_instance2597();
    specparam_declaration2598 specparam_declaration_instance2598();
    specparam_declaration2599 specparam_declaration_instance2599();
    specparam_declaration2600 specparam_declaration_instance2600();
    specparam_declaration2601 specparam_declaration_instance2601();
    specparam_declaration2602 specparam_declaration_instance2602();
    specparam_declaration2603 specparam_declaration_instance2603();
    specparam_declaration2604 specparam_declaration_instance2604();
    specparam_declaration2605 specparam_declaration_instance2605();
    specparam_declaration2606 specparam_declaration_instance2606();
    specparam_declaration2607 specparam_declaration_instance2607();
    specparam_declaration2608 specparam_declaration_instance2608();
    specparam_declaration2609 specparam_declaration_instance2609();
    specparam_declaration2610 specparam_declaration_instance2610();
    specparam_declaration2611 specparam_declaration_instance2611();
    specparam_declaration2612 specparam_declaration_instance2612();
    specparam_declaration2613 specparam_declaration_instance2613();
    specparam_declaration2614 specparam_declaration_instance2614();
    specparam_declaration2615 specparam_declaration_instance2615();
    specparam_declaration2616 specparam_declaration_instance2616();
    specparam_declaration2617 specparam_declaration_instance2617();
    specparam_declaration2618 specparam_declaration_instance2618();
    specparam_declaration2619 specparam_declaration_instance2619();
    specparam_declaration2620 specparam_declaration_instance2620();
    specparam_declaration2621 specparam_declaration_instance2621();
    specparam_declaration2622 specparam_declaration_instance2622();
    specparam_declaration2623 specparam_declaration_instance2623();
    specparam_declaration2624 specparam_declaration_instance2624();
    specparam_declaration2625 specparam_declaration_instance2625();
    specparam_declaration2626 specparam_declaration_instance2626();
    specparam_declaration2627 specparam_declaration_instance2627();
    specparam_declaration2628 specparam_declaration_instance2628();
    specparam_declaration2629 specparam_declaration_instance2629();
    specparam_declaration2630 specparam_declaration_instance2630();
    specparam_declaration2631 specparam_declaration_instance2631();
    specparam_declaration2632 specparam_declaration_instance2632();
    specparam_declaration2633 specparam_declaration_instance2633();
    specparam_declaration2634 specparam_declaration_instance2634();
    specparam_declaration2635 specparam_declaration_instance2635();
    specparam_declaration2636 specparam_declaration_instance2636();
    specparam_declaration2637 specparam_declaration_instance2637();
    specparam_declaration2638 specparam_declaration_instance2638();
    specparam_declaration2639 specparam_declaration_instance2639();
    specparam_declaration2640 specparam_declaration_instance2640();
    specparam_declaration2641 specparam_declaration_instance2641();
    specparam_declaration2642 specparam_declaration_instance2642();
    specparam_declaration2643 specparam_declaration_instance2643();
    specparam_declaration2644 specparam_declaration_instance2644();
    specparam_declaration2645 specparam_declaration_instance2645();
    specparam_declaration2646 specparam_declaration_instance2646();
    specparam_declaration2647 specparam_declaration_instance2647();
    specparam_declaration2648 specparam_declaration_instance2648();
    specparam_declaration2649 specparam_declaration_instance2649();
    specparam_declaration2650 specparam_declaration_instance2650();
    specparam_declaration2651 specparam_declaration_instance2651();
    specparam_declaration2652 specparam_declaration_instance2652();
    specparam_declaration2653 specparam_declaration_instance2653();
    specparam_declaration2654 specparam_declaration_instance2654();
    specparam_declaration2655 specparam_declaration_instance2655();
    specparam_declaration2656 specparam_declaration_instance2656();
    specparam_declaration2657 specparam_declaration_instance2657();
    specparam_declaration2658 specparam_declaration_instance2658();
    specparam_declaration2659 specparam_declaration_instance2659();
    specparam_declaration2660 specparam_declaration_instance2660();
    specparam_declaration2661 specparam_declaration_instance2661();
    specparam_declaration2662 specparam_declaration_instance2662();
    specparam_declaration2663 specparam_declaration_instance2663();
    specparam_declaration2664 specparam_declaration_instance2664();
    specparam_declaration2665 specparam_declaration_instance2665();
    specparam_declaration2666 specparam_declaration_instance2666();
    specparam_declaration2667 specparam_declaration_instance2667();
    specparam_declaration2668 specparam_declaration_instance2668();
    specparam_declaration2669 specparam_declaration_instance2669();
    specparam_declaration2670 specparam_declaration_instance2670();
    specparam_declaration2671 specparam_declaration_instance2671();
    specparam_declaration2672 specparam_declaration_instance2672();
    specparam_declaration2673 specparam_declaration_instance2673();
    specparam_declaration2674 specparam_declaration_instance2674();
    specparam_declaration2675 specparam_declaration_instance2675();
    specparam_declaration2676 specparam_declaration_instance2676();
    specparam_declaration2677 specparam_declaration_instance2677();
    specparam_declaration2678 specparam_declaration_instance2678();
    specparam_declaration2679 specparam_declaration_instance2679();
    specparam_declaration2680 specparam_declaration_instance2680();
    specparam_declaration2681 specparam_declaration_instance2681();
    specparam_declaration2682 specparam_declaration_instance2682();
    specparam_declaration2683 specparam_declaration_instance2683();
    specparam_declaration2684 specparam_declaration_instance2684();
    specparam_declaration2685 specparam_declaration_instance2685();
    specparam_declaration2686 specparam_declaration_instance2686();
    specparam_declaration2687 specparam_declaration_instance2687();
    specparam_declaration2688 specparam_declaration_instance2688();
    specparam_declaration2689 specparam_declaration_instance2689();
    specparam_declaration2690 specparam_declaration_instance2690();
    specparam_declaration2691 specparam_declaration_instance2691();
    specparam_declaration2692 specparam_declaration_instance2692();
    specparam_declaration2693 specparam_declaration_instance2693();
    specparam_declaration2694 specparam_declaration_instance2694();
    specparam_declaration2695 specparam_declaration_instance2695();
    specparam_declaration2696 specparam_declaration_instance2696();
    specparam_declaration2697 specparam_declaration_instance2697();
    specparam_declaration2698 specparam_declaration_instance2698();
    specparam_declaration2699 specparam_declaration_instance2699();
    specparam_declaration2700 specparam_declaration_instance2700();
    specparam_declaration2701 specparam_declaration_instance2701();
    specparam_declaration2702 specparam_declaration_instance2702();
    specparam_declaration2703 specparam_declaration_instance2703();
    specparam_declaration2704 specparam_declaration_instance2704();
    specparam_declaration2705 specparam_declaration_instance2705();
    specparam_declaration2706 specparam_declaration_instance2706();
    specparam_declaration2707 specparam_declaration_instance2707();
    specparam_declaration2708 specparam_declaration_instance2708();
    specparam_declaration2709 specparam_declaration_instance2709();
    specparam_declaration2710 specparam_declaration_instance2710();
    specparam_declaration2711 specparam_declaration_instance2711();
    specparam_declaration2712 specparam_declaration_instance2712();
    specparam_declaration2713 specparam_declaration_instance2713();
    specparam_declaration2714 specparam_declaration_instance2714();
    specparam_declaration2715 specparam_declaration_instance2715();
    specparam_declaration2716 specparam_declaration_instance2716();
    specparam_declaration2717 specparam_declaration_instance2717();
    specparam_declaration2718 specparam_declaration_instance2718();
    specparam_declaration2719 specparam_declaration_instance2719();
    specparam_declaration2720 specparam_declaration_instance2720();
    specparam_declaration2721 specparam_declaration_instance2721();
    specparam_declaration2722 specparam_declaration_instance2722();
    specparam_declaration2723 specparam_declaration_instance2723();
    specparam_declaration2724 specparam_declaration_instance2724();
    specparam_declaration2725 specparam_declaration_instance2725();
    specparam_declaration2726 specparam_declaration_instance2726();
    specparam_declaration2727 specparam_declaration_instance2727();
    specparam_declaration2728 specparam_declaration_instance2728();
    specparam_declaration2729 specparam_declaration_instance2729();
    specparam_declaration2730 specparam_declaration_instance2730();
    specparam_declaration2731 specparam_declaration_instance2731();
    specparam_declaration2732 specparam_declaration_instance2732();
    specparam_declaration2733 specparam_declaration_instance2733();
    specparam_declaration2734 specparam_declaration_instance2734();
    specparam_declaration2735 specparam_declaration_instance2735();
    specparam_declaration2736 specparam_declaration_instance2736();
    specparam_declaration2737 specparam_declaration_instance2737();
    specparam_declaration2738 specparam_declaration_instance2738();
    specparam_declaration2739 specparam_declaration_instance2739();
    specparam_declaration2740 specparam_declaration_instance2740();
    specparam_declaration2741 specparam_declaration_instance2741();
    specparam_declaration2742 specparam_declaration_instance2742();
    specparam_declaration2743 specparam_declaration_instance2743();
    specparam_declaration2744 specparam_declaration_instance2744();
    specparam_declaration2745 specparam_declaration_instance2745();
    specparam_declaration2746 specparam_declaration_instance2746();
    specparam_declaration2747 specparam_declaration_instance2747();
    specparam_declaration2748 specparam_declaration_instance2748();
    specparam_declaration2749 specparam_declaration_instance2749();
    specparam_declaration2750 specparam_declaration_instance2750();
    specparam_declaration2751 specparam_declaration_instance2751();
    specparam_declaration2752 specparam_declaration_instance2752();
    specparam_declaration2753 specparam_declaration_instance2753();
    specparam_declaration2754 specparam_declaration_instance2754();
    specparam_declaration2755 specparam_declaration_instance2755();
    specparam_declaration2756 specparam_declaration_instance2756();
    specparam_declaration2757 specparam_declaration_instance2757();
    specparam_declaration2758 specparam_declaration_instance2758();
    specparam_declaration2759 specparam_declaration_instance2759();
    specparam_declaration2760 specparam_declaration_instance2760();
    specparam_declaration2761 specparam_declaration_instance2761();
    specparam_declaration2762 specparam_declaration_instance2762();
    specparam_declaration2763 specparam_declaration_instance2763();
    specparam_declaration2764 specparam_declaration_instance2764();
    specparam_declaration2765 specparam_declaration_instance2765();
    specparam_declaration2766 specparam_declaration_instance2766();
    specparam_declaration2767 specparam_declaration_instance2767();
    specparam_declaration2768 specparam_declaration_instance2768();
    specparam_declaration2769 specparam_declaration_instance2769();
    specparam_declaration2770 specparam_declaration_instance2770();
    specparam_declaration2771 specparam_declaration_instance2771();
    specparam_declaration2772 specparam_declaration_instance2772();
    specparam_declaration2773 specparam_declaration_instance2773();
    specparam_declaration2774 specparam_declaration_instance2774();
    specparam_declaration2775 specparam_declaration_instance2775();
    specparam_declaration2776 specparam_declaration_instance2776();
    specparam_declaration2777 specparam_declaration_instance2777();
    specparam_declaration2778 specparam_declaration_instance2778();
    specparam_declaration2779 specparam_declaration_instance2779();
    specparam_declaration2780 specparam_declaration_instance2780();
    specparam_declaration2781 specparam_declaration_instance2781();
    specparam_declaration2782 specparam_declaration_instance2782();
    specparam_declaration2783 specparam_declaration_instance2783();
    specparam_declaration2784 specparam_declaration_instance2784();
    specparam_declaration2785 specparam_declaration_instance2785();
    specparam_declaration2786 specparam_declaration_instance2786();
    specparam_declaration2787 specparam_declaration_instance2787();
    specparam_declaration2788 specparam_declaration_instance2788();
    specparam_declaration2789 specparam_declaration_instance2789();
    specparam_declaration2790 specparam_declaration_instance2790();
    specparam_declaration2791 specparam_declaration_instance2791();
    specparam_declaration2792 specparam_declaration_instance2792();
    specparam_declaration2793 specparam_declaration_instance2793();
    specparam_declaration2794 specparam_declaration_instance2794();
    specparam_declaration2795 specparam_declaration_instance2795();
    specparam_declaration2796 specparam_declaration_instance2796();
    specparam_declaration2797 specparam_declaration_instance2797();
    specparam_declaration2798 specparam_declaration_instance2798();
    specparam_declaration2799 specparam_declaration_instance2799();
    specparam_declaration2800 specparam_declaration_instance2800();
    specparam_declaration2801 specparam_declaration_instance2801();
    specparam_declaration2802 specparam_declaration_instance2802();
    specparam_declaration2803 specparam_declaration_instance2803();
    specparam_declaration2804 specparam_declaration_instance2804();
    specparam_declaration2805 specparam_declaration_instance2805();
    specparam_declaration2806 specparam_declaration_instance2806();
    specparam_declaration2807 specparam_declaration_instance2807();
    specparam_declaration2808 specparam_declaration_instance2808();
    specparam_declaration2809 specparam_declaration_instance2809();
    specparam_declaration2810 specparam_declaration_instance2810();
    specparam_declaration2811 specparam_declaration_instance2811();
    specparam_declaration2812 specparam_declaration_instance2812();
    specparam_declaration2813 specparam_declaration_instance2813();
    specparam_declaration2814 specparam_declaration_instance2814();
    specparam_declaration2815 specparam_declaration_instance2815();
    specparam_declaration2816 specparam_declaration_instance2816();
    specparam_declaration2817 specparam_declaration_instance2817();
    specparam_declaration2818 specparam_declaration_instance2818();
    specparam_declaration2819 specparam_declaration_instance2819();
    specparam_declaration2820 specparam_declaration_instance2820();
    specparam_declaration2821 specparam_declaration_instance2821();
    specparam_declaration2822 specparam_declaration_instance2822();
    specparam_declaration2823 specparam_declaration_instance2823();
    specparam_declaration2824 specparam_declaration_instance2824();
    specparam_declaration2825 specparam_declaration_instance2825();
    specparam_declaration2826 specparam_declaration_instance2826();
    specparam_declaration2827 specparam_declaration_instance2827();
    specparam_declaration2828 specparam_declaration_instance2828();
    specparam_declaration2829 specparam_declaration_instance2829();
    specparam_declaration2830 specparam_declaration_instance2830();
    specparam_declaration2831 specparam_declaration_instance2831();
    specparam_declaration2832 specparam_declaration_instance2832();
    specparam_declaration2833 specparam_declaration_instance2833();
    specparam_declaration2834 specparam_declaration_instance2834();
    specparam_declaration2835 specparam_declaration_instance2835();
    specparam_declaration2836 specparam_declaration_instance2836();
    specparam_declaration2837 specparam_declaration_instance2837();
    specparam_declaration2838 specparam_declaration_instance2838();
    specparam_declaration2839 specparam_declaration_instance2839();
    specparam_declaration2840 specparam_declaration_instance2840();
    specparam_declaration2841 specparam_declaration_instance2841();
    specparam_declaration2842 specparam_declaration_instance2842();
    specparam_declaration2843 specparam_declaration_instance2843();
    specparam_declaration2844 specparam_declaration_instance2844();
    specparam_declaration2845 specparam_declaration_instance2845();
    specparam_declaration2846 specparam_declaration_instance2846();
    specparam_declaration2847 specparam_declaration_instance2847();
    specparam_declaration2848 specparam_declaration_instance2848();
    specparam_declaration2849 specparam_declaration_instance2849();
    specparam_declaration2850 specparam_declaration_instance2850();
    specparam_declaration2851 specparam_declaration_instance2851();
    specparam_declaration2852 specparam_declaration_instance2852();
    specparam_declaration2853 specparam_declaration_instance2853();
    specparam_declaration2854 specparam_declaration_instance2854();
    specparam_declaration2855 specparam_declaration_instance2855();
    specparam_declaration2856 specparam_declaration_instance2856();
    specparam_declaration2857 specparam_declaration_instance2857();
    specparam_declaration2858 specparam_declaration_instance2858();
    specparam_declaration2859 specparam_declaration_instance2859();
    specparam_declaration2860 specparam_declaration_instance2860();
    specparam_declaration2861 specparam_declaration_instance2861();
    specparam_declaration2862 specparam_declaration_instance2862();
    specparam_declaration2863 specparam_declaration_instance2863();
    specparam_declaration2864 specparam_declaration_instance2864();
    specparam_declaration2865 specparam_declaration_instance2865();
    specparam_declaration2866 specparam_declaration_instance2866();
    specparam_declaration2867 specparam_declaration_instance2867();
    specparam_declaration2868 specparam_declaration_instance2868();
    specparam_declaration2869 specparam_declaration_instance2869();
    specparam_declaration2870 specparam_declaration_instance2870();
    specparam_declaration2871 specparam_declaration_instance2871();
    specparam_declaration2872 specparam_declaration_instance2872();
    specparam_declaration2873 specparam_declaration_instance2873();
    specparam_declaration2874 specparam_declaration_instance2874();
    specparam_declaration2875 specparam_declaration_instance2875();
    specparam_declaration2876 specparam_declaration_instance2876();
    specparam_declaration2877 specparam_declaration_instance2877();
    specparam_declaration2878 specparam_declaration_instance2878();
    specparam_declaration2879 specparam_declaration_instance2879();
    specparam_declaration2880 specparam_declaration_instance2880();
    specparam_declaration2881 specparam_declaration_instance2881();
    specparam_declaration2882 specparam_declaration_instance2882();
    specparam_declaration2883 specparam_declaration_instance2883();
    specparam_declaration2884 specparam_declaration_instance2884();
    specparam_declaration2885 specparam_declaration_instance2885();
    specparam_declaration2886 specparam_declaration_instance2886();
    specparam_declaration2887 specparam_declaration_instance2887();
    specparam_declaration2888 specparam_declaration_instance2888();
    specparam_declaration2889 specparam_declaration_instance2889();
    specparam_declaration2890 specparam_declaration_instance2890();
    specparam_declaration2891 specparam_declaration_instance2891();
    specparam_declaration2892 specparam_declaration_instance2892();
    specparam_declaration2893 specparam_declaration_instance2893();
    specparam_declaration2894 specparam_declaration_instance2894();
    specparam_declaration2895 specparam_declaration_instance2895();
    specparam_declaration2896 specparam_declaration_instance2896();
    specparam_declaration2897 specparam_declaration_instance2897();
    specparam_declaration2898 specparam_declaration_instance2898();
    specparam_declaration2899 specparam_declaration_instance2899();
    specparam_declaration2900 specparam_declaration_instance2900();
    specparam_declaration2901 specparam_declaration_instance2901();
    specparam_declaration2902 specparam_declaration_instance2902();
    specparam_declaration2903 specparam_declaration_instance2903();
    specparam_declaration2904 specparam_declaration_instance2904();
    specparam_declaration2905 specparam_declaration_instance2905();
    specparam_declaration2906 specparam_declaration_instance2906();
    specparam_declaration2907 specparam_declaration_instance2907();
    specparam_declaration2908 specparam_declaration_instance2908();
    specparam_declaration2909 specparam_declaration_instance2909();
    specparam_declaration2910 specparam_declaration_instance2910();
    specparam_declaration2911 specparam_declaration_instance2911();
    specparam_declaration2912 specparam_declaration_instance2912();
    specparam_declaration2913 specparam_declaration_instance2913();
    specparam_declaration2914 specparam_declaration_instance2914();
    specparam_declaration2915 specparam_declaration_instance2915();
    specparam_declaration2916 specparam_declaration_instance2916();
    specparam_declaration2917 specparam_declaration_instance2917();
    specparam_declaration2918 specparam_declaration_instance2918();
    specparam_declaration2919 specparam_declaration_instance2919();
    specparam_declaration2920 specparam_declaration_instance2920();
    specparam_declaration2921 specparam_declaration_instance2921();
    specparam_declaration2922 specparam_declaration_instance2922();
    specparam_declaration2923 specparam_declaration_instance2923();
    specparam_declaration2924 specparam_declaration_instance2924();
    specparam_declaration2925 specparam_declaration_instance2925();
    specparam_declaration2926 specparam_declaration_instance2926();
    specparam_declaration2927 specparam_declaration_instance2927();
    specparam_declaration2928 specparam_declaration_instance2928();
    specparam_declaration2929 specparam_declaration_instance2929();
    specparam_declaration2930 specparam_declaration_instance2930();
    specparam_declaration2931 specparam_declaration_instance2931();
    specparam_declaration2932 specparam_declaration_instance2932();
    specparam_declaration2933 specparam_declaration_instance2933();
    specparam_declaration2934 specparam_declaration_instance2934();
    specparam_declaration2935 specparam_declaration_instance2935();
    specparam_declaration2936 specparam_declaration_instance2936();
    specparam_declaration2937 specparam_declaration_instance2937();
    specparam_declaration2938 specparam_declaration_instance2938();
    specparam_declaration2939 specparam_declaration_instance2939();
    specparam_declaration2940 specparam_declaration_instance2940();
    specparam_declaration2941 specparam_declaration_instance2941();
    specparam_declaration2942 specparam_declaration_instance2942();
    specparam_declaration2943 specparam_declaration_instance2943();
    specparam_declaration2944 specparam_declaration_instance2944();
    specparam_declaration2945 specparam_declaration_instance2945();
    specparam_declaration2946 specparam_declaration_instance2946();
    specparam_declaration2947 specparam_declaration_instance2947();
    specparam_declaration2948 specparam_declaration_instance2948();
    specparam_declaration2949 specparam_declaration_instance2949();
    specparam_declaration2950 specparam_declaration_instance2950();
    specparam_declaration2951 specparam_declaration_instance2951();
    specparam_declaration2952 specparam_declaration_instance2952();
    specparam_declaration2953 specparam_declaration_instance2953();
    specparam_declaration2954 specparam_declaration_instance2954();
    specparam_declaration2955 specparam_declaration_instance2955();
    specparam_declaration2956 specparam_declaration_instance2956();
    specparam_declaration2957 specparam_declaration_instance2957();
    specparam_declaration2958 specparam_declaration_instance2958();
    specparam_declaration2959 specparam_declaration_instance2959();
    specparam_declaration2960 specparam_declaration_instance2960();
    specparam_declaration2961 specparam_declaration_instance2961();
    specparam_declaration2962 specparam_declaration_instance2962();
    specparam_declaration2963 specparam_declaration_instance2963();
    specparam_declaration2964 specparam_declaration_instance2964();
    specparam_declaration2965 specparam_declaration_instance2965();
    specparam_declaration2966 specparam_declaration_instance2966();
    specparam_declaration2967 specparam_declaration_instance2967();
    specparam_declaration2968 specparam_declaration_instance2968();
    specparam_declaration2969 specparam_declaration_instance2969();
    specparam_declaration2970 specparam_declaration_instance2970();
    specparam_declaration2971 specparam_declaration_instance2971();
    specparam_declaration2972 specparam_declaration_instance2972();
    specparam_declaration2973 specparam_declaration_instance2973();
    specparam_declaration2974 specparam_declaration_instance2974();
    specparam_declaration2975 specparam_declaration_instance2975();
    specparam_declaration2976 specparam_declaration_instance2976();
    specparam_declaration2977 specparam_declaration_instance2977();
    specparam_declaration2978 specparam_declaration_instance2978();
    specparam_declaration2979 specparam_declaration_instance2979();
    specparam_declaration2980 specparam_declaration_instance2980();
    specparam_declaration2981 specparam_declaration_instance2981();
    specparam_declaration2982 specparam_declaration_instance2982();
    specparam_declaration2983 specparam_declaration_instance2983();
    specparam_declaration2984 specparam_declaration_instance2984();
    specparam_declaration2985 specparam_declaration_instance2985();
    specparam_declaration2986 specparam_declaration_instance2986();
    specparam_declaration2987 specparam_declaration_instance2987();
    specparam_declaration2988 specparam_declaration_instance2988();
    specparam_declaration2989 specparam_declaration_instance2989();
    specparam_declaration2990 specparam_declaration_instance2990();
    specparam_declaration2991 specparam_declaration_instance2991();
    specparam_declaration2992 specparam_declaration_instance2992();
    specparam_declaration2993 specparam_declaration_instance2993();
    specparam_declaration2994 specparam_declaration_instance2994();
    specparam_declaration2995 specparam_declaration_instance2995();
    specparam_declaration2996 specparam_declaration_instance2996();
    specparam_declaration2997 specparam_declaration_instance2997();
    specparam_declaration2998 specparam_declaration_instance2998();
    specparam_declaration2999 specparam_declaration_instance2999();
    specparam_declaration3000 specparam_declaration_instance3000();
    specparam_declaration3001 specparam_declaration_instance3001();
    specparam_declaration3002 specparam_declaration_instance3002();
    specparam_declaration3003 specparam_declaration_instance3003();
    specparam_declaration3004 specparam_declaration_instance3004();
    specparam_declaration3005 specparam_declaration_instance3005();
    specparam_declaration3006 specparam_declaration_instance3006();
    specparam_declaration3007 specparam_declaration_instance3007();
    specparam_declaration3008 specparam_declaration_instance3008();
    specparam_declaration3009 specparam_declaration_instance3009();
    specparam_declaration3010 specparam_declaration_instance3010();
    specparam_declaration3011 specparam_declaration_instance3011();
    specparam_declaration3012 specparam_declaration_instance3012();
    specparam_declaration3013 specparam_declaration_instance3013();
    specparam_declaration3014 specparam_declaration_instance3014();
    specparam_declaration3015 specparam_declaration_instance3015();
    specparam_declaration3016 specparam_declaration_instance3016();
    specparam_declaration3017 specparam_declaration_instance3017();
    specparam_declaration3018 specparam_declaration_instance3018();
    specparam_declaration3019 specparam_declaration_instance3019();
    specparam_declaration3020 specparam_declaration_instance3020();
    specparam_declaration3021 specparam_declaration_instance3021();
    specparam_declaration3022 specparam_declaration_instance3022();
    specparam_declaration3023 specparam_declaration_instance3023();
    specparam_declaration3024 specparam_declaration_instance3024();
    specparam_declaration3025 specparam_declaration_instance3025();
    specparam_declaration3026 specparam_declaration_instance3026();
    specparam_declaration3027 specparam_declaration_instance3027();
    specparam_declaration3028 specparam_declaration_instance3028();
    specparam_declaration3029 specparam_declaration_instance3029();
    specparam_declaration3030 specparam_declaration_instance3030();
    specparam_declaration3031 specparam_declaration_instance3031();
    specparam_declaration3032 specparam_declaration_instance3032();
    specparam_declaration3033 specparam_declaration_instance3033();
    specparam_declaration3034 specparam_declaration_instance3034();
    specparam_declaration3035 specparam_declaration_instance3035();
    specparam_declaration3036 specparam_declaration_instance3036();
    specparam_declaration3037 specparam_declaration_instance3037();
    specparam_declaration3038 specparam_declaration_instance3038();
    specparam_declaration3039 specparam_declaration_instance3039();
    specparam_declaration3040 specparam_declaration_instance3040();
    specparam_declaration3041 specparam_declaration_instance3041();
    specparam_declaration3042 specparam_declaration_instance3042();
    specparam_declaration3043 specparam_declaration_instance3043();
    specparam_declaration3044 specparam_declaration_instance3044();
    specparam_declaration3045 specparam_declaration_instance3045();
    specparam_declaration3046 specparam_declaration_instance3046();
    specparam_declaration3047 specparam_declaration_instance3047();
    specparam_declaration3048 specparam_declaration_instance3048();
    specparam_declaration3049 specparam_declaration_instance3049();
    specparam_declaration3050 specparam_declaration_instance3050();
    specparam_declaration3051 specparam_declaration_instance3051();
    specparam_declaration3052 specparam_declaration_instance3052();
    specparam_declaration3053 specparam_declaration_instance3053();
    specparam_declaration3054 specparam_declaration_instance3054();
    specparam_declaration3055 specparam_declaration_instance3055();
    specparam_declaration3056 specparam_declaration_instance3056();
    specparam_declaration3057 specparam_declaration_instance3057();
    specparam_declaration3058 specparam_declaration_instance3058();
    specparam_declaration3059 specparam_declaration_instance3059();
    specparam_declaration3060 specparam_declaration_instance3060();
    specparam_declaration3061 specparam_declaration_instance3061();
    specparam_declaration3062 specparam_declaration_instance3062();
    specparam_declaration3063 specparam_declaration_instance3063();
    specparam_declaration3064 specparam_declaration_instance3064();
    specparam_declaration3065 specparam_declaration_instance3065();
    specparam_declaration3066 specparam_declaration_instance3066();
    specparam_declaration3067 specparam_declaration_instance3067();
    specparam_declaration3068 specparam_declaration_instance3068();
    specparam_declaration3069 specparam_declaration_instance3069();
    specparam_declaration3070 specparam_declaration_instance3070();
    specparam_declaration3071 specparam_declaration_instance3071();
    specparam_declaration3072 specparam_declaration_instance3072();
    specparam_declaration3073 specparam_declaration_instance3073();
    specparam_declaration3074 specparam_declaration_instance3074();
    specparam_declaration3075 specparam_declaration_instance3075();
    specparam_declaration3076 specparam_declaration_instance3076();
    specparam_declaration3077 specparam_declaration_instance3077();
    specparam_declaration3078 specparam_declaration_instance3078();
    specparam_declaration3079 specparam_declaration_instance3079();
    specparam_declaration3080 specparam_declaration_instance3080();
    specparam_declaration3081 specparam_declaration_instance3081();
    specparam_declaration3082 specparam_declaration_instance3082();
    specparam_declaration3083 specparam_declaration_instance3083();
    specparam_declaration3084 specparam_declaration_instance3084();
    specparam_declaration3085 specparam_declaration_instance3085();
    specparam_declaration3086 specparam_declaration_instance3086();
    specparam_declaration3087 specparam_declaration_instance3087();
    specparam_declaration3088 specparam_declaration_instance3088();
    specparam_declaration3089 specparam_declaration_instance3089();
    specparam_declaration3090 specparam_declaration_instance3090();
    specparam_declaration3091 specparam_declaration_instance3091();
    specparam_declaration3092 specparam_declaration_instance3092();
    specparam_declaration3093 specparam_declaration_instance3093();
    specparam_declaration3094 specparam_declaration_instance3094();
    specparam_declaration3095 specparam_declaration_instance3095();
    specparam_declaration3096 specparam_declaration_instance3096();
    specparam_declaration3097 specparam_declaration_instance3097();
    specparam_declaration3098 specparam_declaration_instance3098();
    specparam_declaration3099 specparam_declaration_instance3099();
    specparam_declaration3100 specparam_declaration_instance3100();
    specparam_declaration3101 specparam_declaration_instance3101();
    specparam_declaration3102 specparam_declaration_instance3102();
    specparam_declaration3103 specparam_declaration_instance3103();
    specparam_declaration3104 specparam_declaration_instance3104();
    specparam_declaration3105 specparam_declaration_instance3105();
    specparam_declaration3106 specparam_declaration_instance3106();
    specparam_declaration3107 specparam_declaration_instance3107();
    specparam_declaration3108 specparam_declaration_instance3108();
    specparam_declaration3109 specparam_declaration_instance3109();
    specparam_declaration3110 specparam_declaration_instance3110();
    specparam_declaration3111 specparam_declaration_instance3111();
    specparam_declaration3112 specparam_declaration_instance3112();
    specparam_declaration3113 specparam_declaration_instance3113();
    specparam_declaration3114 specparam_declaration_instance3114();
    specparam_declaration3115 specparam_declaration_instance3115();
    specparam_declaration3116 specparam_declaration_instance3116();
    specparam_declaration3117 specparam_declaration_instance3117();
    specparam_declaration3118 specparam_declaration_instance3118();
    specparam_declaration3119 specparam_declaration_instance3119();
    specparam_declaration3120 specparam_declaration_instance3120();
    specparam_declaration3121 specparam_declaration_instance3121();
    specparam_declaration3122 specparam_declaration_instance3122();
    specparam_declaration3123 specparam_declaration_instance3123();
    specparam_declaration3124 specparam_declaration_instance3124();
    specparam_declaration3125 specparam_declaration_instance3125();
    specparam_declaration3126 specparam_declaration_instance3126();
    specparam_declaration3127 specparam_declaration_instance3127();
    specparam_declaration3128 specparam_declaration_instance3128();
    specparam_declaration3129 specparam_declaration_instance3129();
    specparam_declaration3130 specparam_declaration_instance3130();
    specparam_declaration3131 specparam_declaration_instance3131();
    specparam_declaration3132 specparam_declaration_instance3132();
    specparam_declaration3133 specparam_declaration_instance3133();
    specparam_declaration3134 specparam_declaration_instance3134();
    specparam_declaration3135 specparam_declaration_instance3135();
    specparam_declaration3136 specparam_declaration_instance3136();
    specparam_declaration3137 specparam_declaration_instance3137();
    specparam_declaration3138 specparam_declaration_instance3138();
    specparam_declaration3139 specparam_declaration_instance3139();
    specparam_declaration3140 specparam_declaration_instance3140();
    specparam_declaration3141 specparam_declaration_instance3141();
    specparam_declaration3142 specparam_declaration_instance3142();
    specparam_declaration3143 specparam_declaration_instance3143();
    specparam_declaration3144 specparam_declaration_instance3144();
    specparam_declaration3145 specparam_declaration_instance3145();
    specparam_declaration3146 specparam_declaration_instance3146();
    specparam_declaration3147 specparam_declaration_instance3147();
    specparam_declaration3148 specparam_declaration_instance3148();
    specparam_declaration3149 specparam_declaration_instance3149();
    specparam_declaration3150 specparam_declaration_instance3150();
    specparam_declaration3151 specparam_declaration_instance3151();
    specparam_declaration3152 specparam_declaration_instance3152();
    specparam_declaration3153 specparam_declaration_instance3153();
    specparam_declaration3154 specparam_declaration_instance3154();
    specparam_declaration3155 specparam_declaration_instance3155();
    specparam_declaration3156 specparam_declaration_instance3156();
    specparam_declaration3157 specparam_declaration_instance3157();
    specparam_declaration3158 specparam_declaration_instance3158();
    specparam_declaration3159 specparam_declaration_instance3159();
    specparam_declaration3160 specparam_declaration_instance3160();
    specparam_declaration3161 specparam_declaration_instance3161();
    specparam_declaration3162 specparam_declaration_instance3162();
    specparam_declaration3163 specparam_declaration_instance3163();
    specparam_declaration3164 specparam_declaration_instance3164();
    specparam_declaration3165 specparam_declaration_instance3165();
    specparam_declaration3166 specparam_declaration_instance3166();
    specparam_declaration3167 specparam_declaration_instance3167();
    specparam_declaration3168 specparam_declaration_instance3168();
    specparam_declaration3169 specparam_declaration_instance3169();
    specparam_declaration3170 specparam_declaration_instance3170();
    specparam_declaration3171 specparam_declaration_instance3171();
    specparam_declaration3172 specparam_declaration_instance3172();
    specparam_declaration3173 specparam_declaration_instance3173();
    specparam_declaration3174 specparam_declaration_instance3174();
    specparam_declaration3175 specparam_declaration_instance3175();
    specparam_declaration3176 specparam_declaration_instance3176();
    specparam_declaration3177 specparam_declaration_instance3177();
    specparam_declaration3178 specparam_declaration_instance3178();
    specparam_declaration3179 specparam_declaration_instance3179();
    specparam_declaration3180 specparam_declaration_instance3180();
    specparam_declaration3181 specparam_declaration_instance3181();
    specparam_declaration3182 specparam_declaration_instance3182();
    specparam_declaration3183 specparam_declaration_instance3183();
    specparam_declaration3184 specparam_declaration_instance3184();
    specparam_declaration3185 specparam_declaration_instance3185();
    specparam_declaration3186 specparam_declaration_instance3186();
    specparam_declaration3187 specparam_declaration_instance3187();
    specparam_declaration3188 specparam_declaration_instance3188();
    specparam_declaration3189 specparam_declaration_instance3189();
    specparam_declaration3190 specparam_declaration_instance3190();
    specparam_declaration3191 specparam_declaration_instance3191();
    specparam_declaration3192 specparam_declaration_instance3192();
    specparam_declaration3193 specparam_declaration_instance3193();
    specparam_declaration3194 specparam_declaration_instance3194();
    specparam_declaration3195 specparam_declaration_instance3195();
    specparam_declaration3196 specparam_declaration_instance3196();
    specparam_declaration3197 specparam_declaration_instance3197();
    specparam_declaration3198 specparam_declaration_instance3198();
    specparam_declaration3199 specparam_declaration_instance3199();
    specparam_declaration3200 specparam_declaration_instance3200();
    specparam_declaration3201 specparam_declaration_instance3201();
    specparam_declaration3202 specparam_declaration_instance3202();
    specparam_declaration3203 specparam_declaration_instance3203();
    specparam_declaration3204 specparam_declaration_instance3204();
    specparam_declaration3205 specparam_declaration_instance3205();
    specparam_declaration3206 specparam_declaration_instance3206();
    specparam_declaration3207 specparam_declaration_instance3207();
    specparam_declaration3208 specparam_declaration_instance3208();
    specparam_declaration3209 specparam_declaration_instance3209();
    specparam_declaration3210 specparam_declaration_instance3210();
    specparam_declaration3211 specparam_declaration_instance3211();
    specparam_declaration3212 specparam_declaration_instance3212();
    specparam_declaration3213 specparam_declaration_instance3213();
    specparam_declaration3214 specparam_declaration_instance3214();
    specparam_declaration3215 specparam_declaration_instance3215();
    specparam_declaration3216 specparam_declaration_instance3216();
    specparam_declaration3217 specparam_declaration_instance3217();
    specparam_declaration3218 specparam_declaration_instance3218();
    specparam_declaration3219 specparam_declaration_instance3219();
    specparam_declaration3220 specparam_declaration_instance3220();
    specparam_declaration3221 specparam_declaration_instance3221();
    specparam_declaration3222 specparam_declaration_instance3222();
    specparam_declaration3223 specparam_declaration_instance3223();
    specparam_declaration3224 specparam_declaration_instance3224();
    specparam_declaration3225 specparam_declaration_instance3225();
    specparam_declaration3226 specparam_declaration_instance3226();
    specparam_declaration3227 specparam_declaration_instance3227();
    specparam_declaration3228 specparam_declaration_instance3228();
    specparam_declaration3229 specparam_declaration_instance3229();
    specparam_declaration3230 specparam_declaration_instance3230();
    specparam_declaration3231 specparam_declaration_instance3231();
    specparam_declaration3232 specparam_declaration_instance3232();
    specparam_declaration3233 specparam_declaration_instance3233();
    specparam_declaration3234 specparam_declaration_instance3234();
    specparam_declaration3235 specparam_declaration_instance3235();
    specparam_declaration3236 specparam_declaration_instance3236();
    specparam_declaration3237 specparam_declaration_instance3237();
    specparam_declaration3238 specparam_declaration_instance3238();
    specparam_declaration3239 specparam_declaration_instance3239();
    specparam_declaration3240 specparam_declaration_instance3240();
    specparam_declaration3241 specparam_declaration_instance3241();
    specparam_declaration3242 specparam_declaration_instance3242();
    specparam_declaration3243 specparam_declaration_instance3243();
    specparam_declaration3244 specparam_declaration_instance3244();
    specparam_declaration3245 specparam_declaration_instance3245();
    specparam_declaration3246 specparam_declaration_instance3246();
    specparam_declaration3247 specparam_declaration_instance3247();
    specparam_declaration3248 specparam_declaration_instance3248();
    specparam_declaration3249 specparam_declaration_instance3249();
    specparam_declaration3250 specparam_declaration_instance3250();
    specparam_declaration3251 specparam_declaration_instance3251();
    specparam_declaration3252 specparam_declaration_instance3252();
    specparam_declaration3253 specparam_declaration_instance3253();
    specparam_declaration3254 specparam_declaration_instance3254();
    specparam_declaration3255 specparam_declaration_instance3255();
    specparam_declaration3256 specparam_declaration_instance3256();
    specparam_declaration3257 specparam_declaration_instance3257();
    specparam_declaration3258 specparam_declaration_instance3258();
    specparam_declaration3259 specparam_declaration_instance3259();
    specparam_declaration3260 specparam_declaration_instance3260();
    specparam_declaration3261 specparam_declaration_instance3261();
    specparam_declaration3262 specparam_declaration_instance3262();
    specparam_declaration3263 specparam_declaration_instance3263();
    specparam_declaration3264 specparam_declaration_instance3264();
    specparam_declaration3265 specparam_declaration_instance3265();
    specparam_declaration3266 specparam_declaration_instance3266();
    specparam_declaration3267 specparam_declaration_instance3267();
    specparam_declaration3268 specparam_declaration_instance3268();
    specparam_declaration3269 specparam_declaration_instance3269();
    specparam_declaration3270 specparam_declaration_instance3270();
    specparam_declaration3271 specparam_declaration_instance3271();
    specparam_declaration3272 specparam_declaration_instance3272();
    specparam_declaration3273 specparam_declaration_instance3273();
    specparam_declaration3274 specparam_declaration_instance3274();
    specparam_declaration3275 specparam_declaration_instance3275();
    specparam_declaration3276 specparam_declaration_instance3276();
    specparam_declaration3277 specparam_declaration_instance3277();
    specparam_declaration3278 specparam_declaration_instance3278();
    specparam_declaration3279 specparam_declaration_instance3279();
    specparam_declaration3280 specparam_declaration_instance3280();
    specparam_declaration3281 specparam_declaration_instance3281();
    specparam_declaration3282 specparam_declaration_instance3282();
    specparam_declaration3283 specparam_declaration_instance3283();
    specparam_declaration3284 specparam_declaration_instance3284();
    specparam_declaration3285 specparam_declaration_instance3285();
    specparam_declaration3286 specparam_declaration_instance3286();
    specparam_declaration3287 specparam_declaration_instance3287();
    specparam_declaration3288 specparam_declaration_instance3288();
    specparam_declaration3289 specparam_declaration_instance3289();
    specparam_declaration3290 specparam_declaration_instance3290();
    specparam_declaration3291 specparam_declaration_instance3291();
    specparam_declaration3292 specparam_declaration_instance3292();
    specparam_declaration3293 specparam_declaration_instance3293();
    specparam_declaration3294 specparam_declaration_instance3294();
    specparam_declaration3295 specparam_declaration_instance3295();
    specparam_declaration3296 specparam_declaration_instance3296();
    specparam_declaration3297 specparam_declaration_instance3297();
    specparam_declaration3298 specparam_declaration_instance3298();
    specparam_declaration3299 specparam_declaration_instance3299();
    specparam_declaration3300 specparam_declaration_instance3300();
    specparam_declaration3301 specparam_declaration_instance3301();
    specparam_declaration3302 specparam_declaration_instance3302();
    specparam_declaration3303 specparam_declaration_instance3303();
    specparam_declaration3304 specparam_declaration_instance3304();
    specparam_declaration3305 specparam_declaration_instance3305();
    specparam_declaration3306 specparam_declaration_instance3306();
    specparam_declaration3307 specparam_declaration_instance3307();
    specparam_declaration3308 specparam_declaration_instance3308();
    specparam_declaration3309 specparam_declaration_instance3309();
    specparam_declaration3310 specparam_declaration_instance3310();
    specparam_declaration3311 specparam_declaration_instance3311();
    specparam_declaration3312 specparam_declaration_instance3312();
    specparam_declaration3313 specparam_declaration_instance3313();
    specparam_declaration3314 specparam_declaration_instance3314();
    specparam_declaration3315 specparam_declaration_instance3315();
    specparam_declaration3316 specparam_declaration_instance3316();
    specparam_declaration3317 specparam_declaration_instance3317();
    specparam_declaration3318 specparam_declaration_instance3318();
    specparam_declaration3319 specparam_declaration_instance3319();
    specparam_declaration3320 specparam_declaration_instance3320();
    specparam_declaration3321 specparam_declaration_instance3321();
    specparam_declaration3322 specparam_declaration_instance3322();
    specparam_declaration3323 specparam_declaration_instance3323();
    specparam_declaration3324 specparam_declaration_instance3324();
    specparam_declaration3325 specparam_declaration_instance3325();
    specparam_declaration3326 specparam_declaration_instance3326();
    specparam_declaration3327 specparam_declaration_instance3327();
    specparam_declaration3328 specparam_declaration_instance3328();
    specparam_declaration3329 specparam_declaration_instance3329();
    specparam_declaration3330 specparam_declaration_instance3330();
    specparam_declaration3331 specparam_declaration_instance3331();
    specparam_declaration3332 specparam_declaration_instance3332();
    specparam_declaration3333 specparam_declaration_instance3333();
    specparam_declaration3334 specparam_declaration_instance3334();
    specparam_declaration3335 specparam_declaration_instance3335();
    specparam_declaration3336 specparam_declaration_instance3336();
    specparam_declaration3337 specparam_declaration_instance3337();
    specparam_declaration3338 specparam_declaration_instance3338();
    specparam_declaration3339 specparam_declaration_instance3339();
    specparam_declaration3340 specparam_declaration_instance3340();
    specparam_declaration3341 specparam_declaration_instance3341();
    specparam_declaration3342 specparam_declaration_instance3342();
    specparam_declaration3343 specparam_declaration_instance3343();
    specparam_declaration3344 specparam_declaration_instance3344();
    specparam_declaration3345 specparam_declaration_instance3345();
    specparam_declaration3346 specparam_declaration_instance3346();
    specparam_declaration3347 specparam_declaration_instance3347();
    specparam_declaration3348 specparam_declaration_instance3348();
    specparam_declaration3349 specparam_declaration_instance3349();
    specparam_declaration3350 specparam_declaration_instance3350();
    specparam_declaration3351 specparam_declaration_instance3351();
    specparam_declaration3352 specparam_declaration_instance3352();
    specparam_declaration3353 specparam_declaration_instance3353();
    specparam_declaration3354 specparam_declaration_instance3354();
    specparam_declaration3355 specparam_declaration_instance3355();
    specparam_declaration3356 specparam_declaration_instance3356();
    specparam_declaration3357 specparam_declaration_instance3357();
    specparam_declaration3358 specparam_declaration_instance3358();
    specparam_declaration3359 specparam_declaration_instance3359();
    specparam_declaration3360 specparam_declaration_instance3360();
    specparam_declaration3361 specparam_declaration_instance3361();
    specparam_declaration3362 specparam_declaration_instance3362();
    specparam_declaration3363 specparam_declaration_instance3363();
    specparam_declaration3364 specparam_declaration_instance3364();
    specparam_declaration3365 specparam_declaration_instance3365();
    specparam_declaration3366 specparam_declaration_instance3366();
    specparam_declaration3367 specparam_declaration_instance3367();
    specparam_declaration3368 specparam_declaration_instance3368();
    specparam_declaration3369 specparam_declaration_instance3369();
    specparam_declaration3370 specparam_declaration_instance3370();
    specparam_declaration3371 specparam_declaration_instance3371();
    specparam_declaration3372 specparam_declaration_instance3372();
    specparam_declaration3373 specparam_declaration_instance3373();
    specparam_declaration3374 specparam_declaration_instance3374();
    specparam_declaration3375 specparam_declaration_instance3375();
    specparam_declaration3376 specparam_declaration_instance3376();
    specparam_declaration3377 specparam_declaration_instance3377();
    specparam_declaration3378 specparam_declaration_instance3378();
    specparam_declaration3379 specparam_declaration_instance3379();
    specparam_declaration3380 specparam_declaration_instance3380();
    specparam_declaration3381 specparam_declaration_instance3381();
    specparam_declaration3382 specparam_declaration_instance3382();
    specparam_declaration3383 specparam_declaration_instance3383();
    specparam_declaration3384 specparam_declaration_instance3384();
    specparam_declaration3385 specparam_declaration_instance3385();
    specparam_declaration3386 specparam_declaration_instance3386();
    specparam_declaration3387 specparam_declaration_instance3387();
    specparam_declaration3388 specparam_declaration_instance3388();
    specparam_declaration3389 specparam_declaration_instance3389();
    specparam_declaration3390 specparam_declaration_instance3390();
    specparam_declaration3391 specparam_declaration_instance3391();
    specparam_declaration3392 specparam_declaration_instance3392();
    specparam_declaration3393 specparam_declaration_instance3393();
    specparam_declaration3394 specparam_declaration_instance3394();
    specparam_declaration3395 specparam_declaration_instance3395();
    specparam_declaration3396 specparam_declaration_instance3396();
    specparam_declaration3397 specparam_declaration_instance3397();
    specparam_declaration3398 specparam_declaration_instance3398();
    specparam_declaration3399 specparam_declaration_instance3399();
    specparam_declaration3400 specparam_declaration_instance3400();
    specparam_declaration3401 specparam_declaration_instance3401();
    specparam_declaration3402 specparam_declaration_instance3402();
    specparam_declaration3403 specparam_declaration_instance3403();
    specparam_declaration3404 specparam_declaration_instance3404();
    specparam_declaration3405 specparam_declaration_instance3405();
    specparam_declaration3406 specparam_declaration_instance3406();
    specparam_declaration3407 specparam_declaration_instance3407();
    specparam_declaration3408 specparam_declaration_instance3408();
    specparam_declaration3409 specparam_declaration_instance3409();
    specparam_declaration3410 specparam_declaration_instance3410();
    specparam_declaration3411 specparam_declaration_instance3411();
    specparam_declaration3412 specparam_declaration_instance3412();
    specparam_declaration3413 specparam_declaration_instance3413();
    specparam_declaration3414 specparam_declaration_instance3414();
    specparam_declaration3415 specparam_declaration_instance3415();
    specparam_declaration3416 specparam_declaration_instance3416();
    specparam_declaration3417 specparam_declaration_instance3417();
    specparam_declaration3418 specparam_declaration_instance3418();
    specparam_declaration3419 specparam_declaration_instance3419();
    specparam_declaration3420 specparam_declaration_instance3420();
    specparam_declaration3421 specparam_declaration_instance3421();
    specparam_declaration3422 specparam_declaration_instance3422();
    specparam_declaration3423 specparam_declaration_instance3423();
    specparam_declaration3424 specparam_declaration_instance3424();
    specparam_declaration3425 specparam_declaration_instance3425();
    specparam_declaration3426 specparam_declaration_instance3426();
    specparam_declaration3427 specparam_declaration_instance3427();
    specparam_declaration3428 specparam_declaration_instance3428();
    specparam_declaration3429 specparam_declaration_instance3429();
    specparam_declaration3430 specparam_declaration_instance3430();
    specparam_declaration3431 specparam_declaration_instance3431();
    specparam_declaration3432 specparam_declaration_instance3432();
    specparam_declaration3433 specparam_declaration_instance3433();
    specparam_declaration3434 specparam_declaration_instance3434();
    specparam_declaration3435 specparam_declaration_instance3435();
    specparam_declaration3436 specparam_declaration_instance3436();
    specparam_declaration3437 specparam_declaration_instance3437();
    specparam_declaration3438 specparam_declaration_instance3438();
    specparam_declaration3439 specparam_declaration_instance3439();
    specparam_declaration3440 specparam_declaration_instance3440();
    specparam_declaration3441 specparam_declaration_instance3441();
    specparam_declaration3442 specparam_declaration_instance3442();
    specparam_declaration3443 specparam_declaration_instance3443();
    specparam_declaration3444 specparam_declaration_instance3444();
    specparam_declaration3445 specparam_declaration_instance3445();
    specparam_declaration3446 specparam_declaration_instance3446();
    specparam_declaration3447 specparam_declaration_instance3447();
    specparam_declaration3448 specparam_declaration_instance3448();
    specparam_declaration3449 specparam_declaration_instance3449();
    specparam_declaration3450 specparam_declaration_instance3450();
    specparam_declaration3451 specparam_declaration_instance3451();
    specparam_declaration3452 specparam_declaration_instance3452();
    specparam_declaration3453 specparam_declaration_instance3453();
    specparam_declaration3454 specparam_declaration_instance3454();
    specparam_declaration3455 specparam_declaration_instance3455();
    specparam_declaration3456 specparam_declaration_instance3456();
    specparam_declaration3457 specparam_declaration_instance3457();
    specparam_declaration3458 specparam_declaration_instance3458();
    specparam_declaration3459 specparam_declaration_instance3459();
    specparam_declaration3460 specparam_declaration_instance3460();
    specparam_declaration3461 specparam_declaration_instance3461();
    specparam_declaration3462 specparam_declaration_instance3462();
    specparam_declaration3463 specparam_declaration_instance3463();
    specparam_declaration3464 specparam_declaration_instance3464();
    specparam_declaration3465 specparam_declaration_instance3465();
    specparam_declaration3466 specparam_declaration_instance3466();
    specparam_declaration3467 specparam_declaration_instance3467();
    specparam_declaration3468 specparam_declaration_instance3468();
    specparam_declaration3469 specparam_declaration_instance3469();
    specparam_declaration3470 specparam_declaration_instance3470();
    specparam_declaration3471 specparam_declaration_instance3471();
    specparam_declaration3472 specparam_declaration_instance3472();
    specparam_declaration3473 specparam_declaration_instance3473();
    specparam_declaration3474 specparam_declaration_instance3474();
    specparam_declaration3475 specparam_declaration_instance3475();
    specparam_declaration3476 specparam_declaration_instance3476();
    specparam_declaration3477 specparam_declaration_instance3477();
    specparam_declaration3478 specparam_declaration_instance3478();
    specparam_declaration3479 specparam_declaration_instance3479();
    specparam_declaration3480 specparam_declaration_instance3480();
    specparam_declaration3481 specparam_declaration_instance3481();
    specparam_declaration3482 specparam_declaration_instance3482();
    specparam_declaration3483 specparam_declaration_instance3483();
    specparam_declaration3484 specparam_declaration_instance3484();
    specparam_declaration3485 specparam_declaration_instance3485();
    specparam_declaration3486 specparam_declaration_instance3486();
    specparam_declaration3487 specparam_declaration_instance3487();
    specparam_declaration3488 specparam_declaration_instance3488();
    specparam_declaration3489 specparam_declaration_instance3489();
    specparam_declaration3490 specparam_declaration_instance3490();
    specparam_declaration3491 specparam_declaration_instance3491();
    specparam_declaration3492 specparam_declaration_instance3492();
    specparam_declaration3493 specparam_declaration_instance3493();
    specparam_declaration3494 specparam_declaration_instance3494();
    specparam_declaration3495 specparam_declaration_instance3495();
    specparam_declaration3496 specparam_declaration_instance3496();
    specparam_declaration3497 specparam_declaration_instance3497();
    specparam_declaration3498 specparam_declaration_instance3498();
    specparam_declaration3499 specparam_declaration_instance3499();
    specparam_declaration3500 specparam_declaration_instance3500();
    specparam_declaration3501 specparam_declaration_instance3501();
    specparam_declaration3502 specparam_declaration_instance3502();
    specparam_declaration3503 specparam_declaration_instance3503();
    specparam_declaration3504 specparam_declaration_instance3504();
    specparam_declaration3505 specparam_declaration_instance3505();
    specparam_declaration3506 specparam_declaration_instance3506();
    specparam_declaration3507 specparam_declaration_instance3507();
    specparam_declaration3508 specparam_declaration_instance3508();
    specparam_declaration3509 specparam_declaration_instance3509();
    specparam_declaration3510 specparam_declaration_instance3510();
    specparam_declaration3511 specparam_declaration_instance3511();
    specparam_declaration3512 specparam_declaration_instance3512();
    specparam_declaration3513 specparam_declaration_instance3513();
    specparam_declaration3514 specparam_declaration_instance3514();
    specparam_declaration3515 specparam_declaration_instance3515();
    specparam_declaration3516 specparam_declaration_instance3516();
    specparam_declaration3517 specparam_declaration_instance3517();
    specparam_declaration3518 specparam_declaration_instance3518();
    specparam_declaration3519 specparam_declaration_instance3519();
    specparam_declaration3520 specparam_declaration_instance3520();
    specparam_declaration3521 specparam_declaration_instance3521();
    specparam_declaration3522 specparam_declaration_instance3522();
    specparam_declaration3523 specparam_declaration_instance3523();
    specparam_declaration3524 specparam_declaration_instance3524();
    specparam_declaration3525 specparam_declaration_instance3525();
    specparam_declaration3526 specparam_declaration_instance3526();
    specparam_declaration3527 specparam_declaration_instance3527();
    specparam_declaration3528 specparam_declaration_instance3528();
    specparam_declaration3529 specparam_declaration_instance3529();
    specparam_declaration3530 specparam_declaration_instance3530();
    specparam_declaration3531 specparam_declaration_instance3531();
    specparam_declaration3532 specparam_declaration_instance3532();
    specparam_declaration3533 specparam_declaration_instance3533();
    specparam_declaration3534 specparam_declaration_instance3534();
    specparam_declaration3535 specparam_declaration_instance3535();
    specparam_declaration3536 specparam_declaration_instance3536();
    specparam_declaration3537 specparam_declaration_instance3537();
    specparam_declaration3538 specparam_declaration_instance3538();
    specparam_declaration3539 specparam_declaration_instance3539();
    specparam_declaration3540 specparam_declaration_instance3540();
    specparam_declaration3541 specparam_declaration_instance3541();
    specparam_declaration3542 specparam_declaration_instance3542();
    specparam_declaration3543 specparam_declaration_instance3543();
    specparam_declaration3544 specparam_declaration_instance3544();
    specparam_declaration3545 specparam_declaration_instance3545();
    specparam_declaration3546 specparam_declaration_instance3546();
    specparam_declaration3547 specparam_declaration_instance3547();
    specparam_declaration3548 specparam_declaration_instance3548();
    specparam_declaration3549 specparam_declaration_instance3549();
    specparam_declaration3550 specparam_declaration_instance3550();
    specparam_declaration3551 specparam_declaration_instance3551();
    specparam_declaration3552 specparam_declaration_instance3552();
    specparam_declaration3553 specparam_declaration_instance3553();
    specparam_declaration3554 specparam_declaration_instance3554();
    specparam_declaration3555 specparam_declaration_instance3555();
    specparam_declaration3556 specparam_declaration_instance3556();
    specparam_declaration3557 specparam_declaration_instance3557();
    specparam_declaration3558 specparam_declaration_instance3558();
    specparam_declaration3559 specparam_declaration_instance3559();
    specparam_declaration3560 specparam_declaration_instance3560();
    specparam_declaration3561 specparam_declaration_instance3561();
    specparam_declaration3562 specparam_declaration_instance3562();
    specparam_declaration3563 specparam_declaration_instance3563();
    specparam_declaration3564 specparam_declaration_instance3564();
    specparam_declaration3565 specparam_declaration_instance3565();
    specparam_declaration3566 specparam_declaration_instance3566();
    specparam_declaration3567 specparam_declaration_instance3567();
    specparam_declaration3568 specparam_declaration_instance3568();
    specparam_declaration3569 specparam_declaration_instance3569();
    specparam_declaration3570 specparam_declaration_instance3570();
    specparam_declaration3571 specparam_declaration_instance3571();
    specparam_declaration3572 specparam_declaration_instance3572();
    specparam_declaration3573 specparam_declaration_instance3573();
    specparam_declaration3574 specparam_declaration_instance3574();
    specparam_declaration3575 specparam_declaration_instance3575();
    specparam_declaration3576 specparam_declaration_instance3576();
    specparam_declaration3577 specparam_declaration_instance3577();
    specparam_declaration3578 specparam_declaration_instance3578();
    specparam_declaration3579 specparam_declaration_instance3579();
    specparam_declaration3580 specparam_declaration_instance3580();
    specparam_declaration3581 specparam_declaration_instance3581();
    specparam_declaration3582 specparam_declaration_instance3582();
    specparam_declaration3583 specparam_declaration_instance3583();
    specparam_declaration3584 specparam_declaration_instance3584();
    specparam_declaration3585 specparam_declaration_instance3585();
    specparam_declaration3586 specparam_declaration_instance3586();
    specparam_declaration3587 specparam_declaration_instance3587();
    specparam_declaration3588 specparam_declaration_instance3588();
    specparam_declaration3589 specparam_declaration_instance3589();
    specparam_declaration3590 specparam_declaration_instance3590();
    specparam_declaration3591 specparam_declaration_instance3591();
    specparam_declaration3592 specparam_declaration_instance3592();
    specparam_declaration3593 specparam_declaration_instance3593();
    specparam_declaration3594 specparam_declaration_instance3594();
    specparam_declaration3595 specparam_declaration_instance3595();
    specparam_declaration3596 specparam_declaration_instance3596();
    specparam_declaration3597 specparam_declaration_instance3597();
    specparam_declaration3598 specparam_declaration_instance3598();
    specparam_declaration3599 specparam_declaration_instance3599();
    specparam_declaration3600 specparam_declaration_instance3600();
    specparam_declaration3601 specparam_declaration_instance3601();
    specparam_declaration3602 specparam_declaration_instance3602();
    specparam_declaration3603 specparam_declaration_instance3603();
    specparam_declaration3604 specparam_declaration_instance3604();
    specparam_declaration3605 specparam_declaration_instance3605();
    specparam_declaration3606 specparam_declaration_instance3606();
    specparam_declaration3607 specparam_declaration_instance3607();
    specparam_declaration3608 specparam_declaration_instance3608();
    specparam_declaration3609 specparam_declaration_instance3609();
    specparam_declaration3610 specparam_declaration_instance3610();
    specparam_declaration3611 specparam_declaration_instance3611();
    specparam_declaration3612 specparam_declaration_instance3612();
    specparam_declaration3613 specparam_declaration_instance3613();
    specparam_declaration3614 specparam_declaration_instance3614();
    specparam_declaration3615 specparam_declaration_instance3615();
    specparam_declaration3616 specparam_declaration_instance3616();
    specparam_declaration3617 specparam_declaration_instance3617();
    specparam_declaration3618 specparam_declaration_instance3618();
    specparam_declaration3619 specparam_declaration_instance3619();
    specparam_declaration3620 specparam_declaration_instance3620();
    specparam_declaration3621 specparam_declaration_instance3621();
    specparam_declaration3622 specparam_declaration_instance3622();
    specparam_declaration3623 specparam_declaration_instance3623();
    specparam_declaration3624 specparam_declaration_instance3624();
    specparam_declaration3625 specparam_declaration_instance3625();
    specparam_declaration3626 specparam_declaration_instance3626();
    specparam_declaration3627 specparam_declaration_instance3627();
    specparam_declaration3628 specparam_declaration_instance3628();
    specparam_declaration3629 specparam_declaration_instance3629();
    specparam_declaration3630 specparam_declaration_instance3630();
    specparam_declaration3631 specparam_declaration_instance3631();
    specparam_declaration3632 specparam_declaration_instance3632();
    specparam_declaration3633 specparam_declaration_instance3633();
    specparam_declaration3634 specparam_declaration_instance3634();
    specparam_declaration3635 specparam_declaration_instance3635();
    specparam_declaration3636 specparam_declaration_instance3636();
    specparam_declaration3637 specparam_declaration_instance3637();
    specparam_declaration3638 specparam_declaration_instance3638();
    specparam_declaration3639 specparam_declaration_instance3639();
    specparam_declaration3640 specparam_declaration_instance3640();
    specparam_declaration3641 specparam_declaration_instance3641();
    specparam_declaration3642 specparam_declaration_instance3642();
    specparam_declaration3643 specparam_declaration_instance3643();
    specparam_declaration3644 specparam_declaration_instance3644();
    specparam_declaration3645 specparam_declaration_instance3645();
    specparam_declaration3646 specparam_declaration_instance3646();
    specparam_declaration3647 specparam_declaration_instance3647();
    specparam_declaration3648 specparam_declaration_instance3648();
    specparam_declaration3649 specparam_declaration_instance3649();
    specparam_declaration3650 specparam_declaration_instance3650();
    specparam_declaration3651 specparam_declaration_instance3651();
    specparam_declaration3652 specparam_declaration_instance3652();
    specparam_declaration3653 specparam_declaration_instance3653();
    specparam_declaration3654 specparam_declaration_instance3654();
    specparam_declaration3655 specparam_declaration_instance3655();
    specparam_declaration3656 specparam_declaration_instance3656();
    specparam_declaration3657 specparam_declaration_instance3657();
    specparam_declaration3658 specparam_declaration_instance3658();
    specparam_declaration3659 specparam_declaration_instance3659();
    specparam_declaration3660 specparam_declaration_instance3660();
    specparam_declaration3661 specparam_declaration_instance3661();
    specparam_declaration3662 specparam_declaration_instance3662();
    specparam_declaration3663 specparam_declaration_instance3663();
    specparam_declaration3664 specparam_declaration_instance3664();
    specparam_declaration3665 specparam_declaration_instance3665();
    specparam_declaration3666 specparam_declaration_instance3666();
    specparam_declaration3667 specparam_declaration_instance3667();
    specparam_declaration3668 specparam_declaration_instance3668();
    specparam_declaration3669 specparam_declaration_instance3669();
    specparam_declaration3670 specparam_declaration_instance3670();
    specparam_declaration3671 specparam_declaration_instance3671();
    specparam_declaration3672 specparam_declaration_instance3672();
    specparam_declaration3673 specparam_declaration_instance3673();
    specparam_declaration3674 specparam_declaration_instance3674();
    specparam_declaration3675 specparam_declaration_instance3675();
    specparam_declaration3676 specparam_declaration_instance3676();
    specparam_declaration3677 specparam_declaration_instance3677();
    specparam_declaration3678 specparam_declaration_instance3678();
    specparam_declaration3679 specparam_declaration_instance3679();
    specparam_declaration3680 specparam_declaration_instance3680();
    specparam_declaration3681 specparam_declaration_instance3681();
    specparam_declaration3682 specparam_declaration_instance3682();
    specparam_declaration3683 specparam_declaration_instance3683();
    specparam_declaration3684 specparam_declaration_instance3684();
    specparam_declaration3685 specparam_declaration_instance3685();
    specparam_declaration3686 specparam_declaration_instance3686();
    specparam_declaration3687 specparam_declaration_instance3687();
    specparam_declaration3688 specparam_declaration_instance3688();
    specparam_declaration3689 specparam_declaration_instance3689();
    specparam_declaration3690 specparam_declaration_instance3690();
    specparam_declaration3691 specparam_declaration_instance3691();
    specparam_declaration3692 specparam_declaration_instance3692();
    specparam_declaration3693 specparam_declaration_instance3693();
    specparam_declaration3694 specparam_declaration_instance3694();
    specparam_declaration3695 specparam_declaration_instance3695();
    specparam_declaration3696 specparam_declaration_instance3696();
    specparam_declaration3697 specparam_declaration_instance3697();
    specparam_declaration3698 specparam_declaration_instance3698();
    specparam_declaration3699 specparam_declaration_instance3699();
    specparam_declaration3700 specparam_declaration_instance3700();
    specparam_declaration3701 specparam_declaration_instance3701();
    specparam_declaration3702 specparam_declaration_instance3702();
    specparam_declaration3703 specparam_declaration_instance3703();
    specparam_declaration3704 specparam_declaration_instance3704();
    specparam_declaration3705 specparam_declaration_instance3705();
    specparam_declaration3706 specparam_declaration_instance3706();
    specparam_declaration3707 specparam_declaration_instance3707();
    specparam_declaration3708 specparam_declaration_instance3708();
    specparam_declaration3709 specparam_declaration_instance3709();
    specparam_declaration3710 specparam_declaration_instance3710();
    specparam_declaration3711 specparam_declaration_instance3711();
    specparam_declaration3712 specparam_declaration_instance3712();
    specparam_declaration3713 specparam_declaration_instance3713();
    specparam_declaration3714 specparam_declaration_instance3714();
    specparam_declaration3715 specparam_declaration_instance3715();
    specparam_declaration3716 specparam_declaration_instance3716();
    specparam_declaration3717 specparam_declaration_instance3717();
    specparam_declaration3718 specparam_declaration_instance3718();
    specparam_declaration3719 specparam_declaration_instance3719();
    specparam_declaration3720 specparam_declaration_instance3720();
    specparam_declaration3721 specparam_declaration_instance3721();
    specparam_declaration3722 specparam_declaration_instance3722();
    specparam_declaration3723 specparam_declaration_instance3723();
    specparam_declaration3724 specparam_declaration_instance3724();
    specparam_declaration3725 specparam_declaration_instance3725();
    specparam_declaration3726 specparam_declaration_instance3726();
    specparam_declaration3727 specparam_declaration_instance3727();
    specparam_declaration3728 specparam_declaration_instance3728();
    specparam_declaration3729 specparam_declaration_instance3729();
    specparam_declaration3730 specparam_declaration_instance3730();
    specparam_declaration3731 specparam_declaration_instance3731();
    specparam_declaration3732 specparam_declaration_instance3732();
    specparam_declaration3733 specparam_declaration_instance3733();
    specparam_declaration3734 specparam_declaration_instance3734();
    specparam_declaration3735 specparam_declaration_instance3735();
    specparam_declaration3736 specparam_declaration_instance3736();
    specparam_declaration3737 specparam_declaration_instance3737();
    specparam_declaration3738 specparam_declaration_instance3738();
    specparam_declaration3739 specparam_declaration_instance3739();
    specparam_declaration3740 specparam_declaration_instance3740();
    specparam_declaration3741 specparam_declaration_instance3741();
    specparam_declaration3742 specparam_declaration_instance3742();
    specparam_declaration3743 specparam_declaration_instance3743();
    specparam_declaration3744 specparam_declaration_instance3744();
    specparam_declaration3745 specparam_declaration_instance3745();
    specparam_declaration3746 specparam_declaration_instance3746();
    specparam_declaration3747 specparam_declaration_instance3747();
    specparam_declaration3748 specparam_declaration_instance3748();
    specparam_declaration3749 specparam_declaration_instance3749();
    specparam_declaration3750 specparam_declaration_instance3750();
    specparam_declaration3751 specparam_declaration_instance3751();
    specparam_declaration3752 specparam_declaration_instance3752();
    specparam_declaration3753 specparam_declaration_instance3753();
    specparam_declaration3754 specparam_declaration_instance3754();
    specparam_declaration3755 specparam_declaration_instance3755();
    specparam_declaration3756 specparam_declaration_instance3756();
    specparam_declaration3757 specparam_declaration_instance3757();
    specparam_declaration3758 specparam_declaration_instance3758();
    specparam_declaration3759 specparam_declaration_instance3759();
    specparam_declaration3760 specparam_declaration_instance3760();
    specparam_declaration3761 specparam_declaration_instance3761();
    specparam_declaration3762 specparam_declaration_instance3762();
    specparam_declaration3763 specparam_declaration_instance3763();
    specparam_declaration3764 specparam_declaration_instance3764();
    specparam_declaration3765 specparam_declaration_instance3765();
    specparam_declaration3766 specparam_declaration_instance3766();
    specparam_declaration3767 specparam_declaration_instance3767();
    specparam_declaration3768 specparam_declaration_instance3768();
    specparam_declaration3769 specparam_declaration_instance3769();
    specparam_declaration3770 specparam_declaration_instance3770();
    specparam_declaration3771 specparam_declaration_instance3771();
    specparam_declaration3772 specparam_declaration_instance3772();
    specparam_declaration3773 specparam_declaration_instance3773();
    specparam_declaration3774 specparam_declaration_instance3774();
    specparam_declaration3775 specparam_declaration_instance3775();
    specparam_declaration3776 specparam_declaration_instance3776();
    specparam_declaration3777 specparam_declaration_instance3777();
    specparam_declaration3778 specparam_declaration_instance3778();
    specparam_declaration3779 specparam_declaration_instance3779();
    specparam_declaration3780 specparam_declaration_instance3780();
    specparam_declaration3781 specparam_declaration_instance3781();
    specparam_declaration3782 specparam_declaration_instance3782();
    specparam_declaration3783 specparam_declaration_instance3783();
    specparam_declaration3784 specparam_declaration_instance3784();
    specparam_declaration3785 specparam_declaration_instance3785();
    specparam_declaration3786 specparam_declaration_instance3786();
    specparam_declaration3787 specparam_declaration_instance3787();
    specparam_declaration3788 specparam_declaration_instance3788();
    specparam_declaration3789 specparam_declaration_instance3789();
    specparam_declaration3790 specparam_declaration_instance3790();
    specparam_declaration3791 specparam_declaration_instance3791();
    specparam_declaration3792 specparam_declaration_instance3792();
    specparam_declaration3793 specparam_declaration_instance3793();
    specparam_declaration3794 specparam_declaration_instance3794();
    specparam_declaration3795 specparam_declaration_instance3795();
    specparam_declaration3796 specparam_declaration_instance3796();
    specparam_declaration3797 specparam_declaration_instance3797();
    specparam_declaration3798 specparam_declaration_instance3798();
    specparam_declaration3799 specparam_declaration_instance3799();
    specparam_declaration3800 specparam_declaration_instance3800();
    specparam_declaration3801 specparam_declaration_instance3801();
    specparam_declaration3802 specparam_declaration_instance3802();
    specparam_declaration3803 specparam_declaration_instance3803();
    specparam_declaration3804 specparam_declaration_instance3804();
    specparam_declaration3805 specparam_declaration_instance3805();
    specparam_declaration3806 specparam_declaration_instance3806();
    specparam_declaration3807 specparam_declaration_instance3807();
    specparam_declaration3808 specparam_declaration_instance3808();
    specparam_declaration3809 specparam_declaration_instance3809();
    specparam_declaration3810 specparam_declaration_instance3810();
    specparam_declaration3811 specparam_declaration_instance3811();
    specparam_declaration3812 specparam_declaration_instance3812();
    specparam_declaration3813 specparam_declaration_instance3813();
    specparam_declaration3814 specparam_declaration_instance3814();
    specparam_declaration3815 specparam_declaration_instance3815();
    specparam_declaration3816 specparam_declaration_instance3816();
    specparam_declaration3817 specparam_declaration_instance3817();
    specparam_declaration3818 specparam_declaration_instance3818();
    specparam_declaration3819 specparam_declaration_instance3819();
    specparam_declaration3820 specparam_declaration_instance3820();
    specparam_declaration3821 specparam_declaration_instance3821();
    specparam_declaration3822 specparam_declaration_instance3822();
    specparam_declaration3823 specparam_declaration_instance3823();
    specparam_declaration3824 specparam_declaration_instance3824();
    specparam_declaration3825 specparam_declaration_instance3825();
    specparam_declaration3826 specparam_declaration_instance3826();
    specparam_declaration3827 specparam_declaration_instance3827();
    specparam_declaration3828 specparam_declaration_instance3828();
    specparam_declaration3829 specparam_declaration_instance3829();
    specparam_declaration3830 specparam_declaration_instance3830();
    specparam_declaration3831 specparam_declaration_instance3831();
    specparam_declaration3832 specparam_declaration_instance3832();
    specparam_declaration3833 specparam_declaration_instance3833();
    specparam_declaration3834 specparam_declaration_instance3834();
    specparam_declaration3835 specparam_declaration_instance3835();
    specparam_declaration3836 specparam_declaration_instance3836();
    specparam_declaration3837 specparam_declaration_instance3837();
    specparam_declaration3838 specparam_declaration_instance3838();
    specparam_declaration3839 specparam_declaration_instance3839();
    specparam_declaration3840 specparam_declaration_instance3840();
    specparam_declaration3841 specparam_declaration_instance3841();
    specparam_declaration3842 specparam_declaration_instance3842();
    specparam_declaration3843 specparam_declaration_instance3843();
    specparam_declaration3844 specparam_declaration_instance3844();
    specparam_declaration3845 specparam_declaration_instance3845();
    specparam_declaration3846 specparam_declaration_instance3846();
    specparam_declaration3847 specparam_declaration_instance3847();
    specparam_declaration3848 specparam_declaration_instance3848();
    specparam_declaration3849 specparam_declaration_instance3849();
    specparam_declaration3850 specparam_declaration_instance3850();
    specparam_declaration3851 specparam_declaration_instance3851();
    specparam_declaration3852 specparam_declaration_instance3852();
    specparam_declaration3853 specparam_declaration_instance3853();
    specparam_declaration3854 specparam_declaration_instance3854();
    specparam_declaration3855 specparam_declaration_instance3855();
    specparam_declaration3856 specparam_declaration_instance3856();
    specparam_declaration3857 specparam_declaration_instance3857();
    specparam_declaration3858 specparam_declaration_instance3858();
    specparam_declaration3859 specparam_declaration_instance3859();
    specparam_declaration3860 specparam_declaration_instance3860();
    specparam_declaration3861 specparam_declaration_instance3861();
    specparam_declaration3862 specparam_declaration_instance3862();
    specparam_declaration3863 specparam_declaration_instance3863();
    specparam_declaration3864 specparam_declaration_instance3864();
    specparam_declaration3865 specparam_declaration_instance3865();
    specparam_declaration3866 specparam_declaration_instance3866();
    specparam_declaration3867 specparam_declaration_instance3867();
    specparam_declaration3868 specparam_declaration_instance3868();
    specparam_declaration3869 specparam_declaration_instance3869();
    specparam_declaration3870 specparam_declaration_instance3870();
    specparam_declaration3871 specparam_declaration_instance3871();
    specparam_declaration3872 specparam_declaration_instance3872();
    specparam_declaration3873 specparam_declaration_instance3873();
    specparam_declaration3874 specparam_declaration_instance3874();
    specparam_declaration3875 specparam_declaration_instance3875();
    specparam_declaration3876 specparam_declaration_instance3876();
    specparam_declaration3877 specparam_declaration_instance3877();
    specparam_declaration3878 specparam_declaration_instance3878();
    specparam_declaration3879 specparam_declaration_instance3879();
    specparam_declaration3880 specparam_declaration_instance3880();
    specparam_declaration3881 specparam_declaration_instance3881();
    specparam_declaration3882 specparam_declaration_instance3882();
    specparam_declaration3883 specparam_declaration_instance3883();
    specparam_declaration3884 specparam_declaration_instance3884();
    specparam_declaration3885 specparam_declaration_instance3885();
    specparam_declaration3886 specparam_declaration_instance3886();
    specparam_declaration3887 specparam_declaration_instance3887();
    specparam_declaration3888 specparam_declaration_instance3888();
    specparam_declaration3889 specparam_declaration_instance3889();
    specparam_declaration3890 specparam_declaration_instance3890();
    specparam_declaration3891 specparam_declaration_instance3891();
    specparam_declaration3892 specparam_declaration_instance3892();
    specparam_declaration3893 specparam_declaration_instance3893();
    specparam_declaration3894 specparam_declaration_instance3894();
    specparam_declaration3895 specparam_declaration_instance3895();
    specparam_declaration3896 specparam_declaration_instance3896();
    specparam_declaration3897 specparam_declaration_instance3897();
    specparam_declaration3898 specparam_declaration_instance3898();
    specparam_declaration3899 specparam_declaration_instance3899();
    specparam_declaration3900 specparam_declaration_instance3900();
    specparam_declaration3901 specparam_declaration_instance3901();
    specparam_declaration3902 specparam_declaration_instance3902();
    specparam_declaration3903 specparam_declaration_instance3903();
    specparam_declaration3904 specparam_declaration_instance3904();
    specparam_declaration3905 specparam_declaration_instance3905();
    specparam_declaration3906 specparam_declaration_instance3906();
    specparam_declaration3907 specparam_declaration_instance3907();
    specparam_declaration3908 specparam_declaration_instance3908();
    specparam_declaration3909 specparam_declaration_instance3909();
    specparam_declaration3910 specparam_declaration_instance3910();
    specparam_declaration3911 specparam_declaration_instance3911();
    specparam_declaration3912 specparam_declaration_instance3912();
    specparam_declaration3913 specparam_declaration_instance3913();
    specparam_declaration3914 specparam_declaration_instance3914();
    specparam_declaration3915 specparam_declaration_instance3915();
    specparam_declaration3916 specparam_declaration_instance3916();
    specparam_declaration3917 specparam_declaration_instance3917();
    specparam_declaration3918 specparam_declaration_instance3918();
    specparam_declaration3919 specparam_declaration_instance3919();
    specparam_declaration3920 specparam_declaration_instance3920();
    specparam_declaration3921 specparam_declaration_instance3921();
    specparam_declaration3922 specparam_declaration_instance3922();
    specparam_declaration3923 specparam_declaration_instance3923();
    specparam_declaration3924 specparam_declaration_instance3924();
    specparam_declaration3925 specparam_declaration_instance3925();
    specparam_declaration3926 specparam_declaration_instance3926();
    specparam_declaration3927 specparam_declaration_instance3927();
    specparam_declaration3928 specparam_declaration_instance3928();
    specparam_declaration3929 specparam_declaration_instance3929();
    specparam_declaration3930 specparam_declaration_instance3930();
    specparam_declaration3931 specparam_declaration_instance3931();
    specparam_declaration3932 specparam_declaration_instance3932();
    specparam_declaration3933 specparam_declaration_instance3933();
    specparam_declaration3934 specparam_declaration_instance3934();
    specparam_declaration3935 specparam_declaration_instance3935();
    specparam_declaration3936 specparam_declaration_instance3936();
    specparam_declaration3937 specparam_declaration_instance3937();
    specparam_declaration3938 specparam_declaration_instance3938();
    specparam_declaration3939 specparam_declaration_instance3939();
    specparam_declaration3940 specparam_declaration_instance3940();
    specparam_declaration3941 specparam_declaration_instance3941();
    specparam_declaration3942 specparam_declaration_instance3942();
    specparam_declaration3943 specparam_declaration_instance3943();
    specparam_declaration3944 specparam_declaration_instance3944();
    specparam_declaration3945 specparam_declaration_instance3945();
    specparam_declaration3946 specparam_declaration_instance3946();
    specparam_declaration3947 specparam_declaration_instance3947();
    specparam_declaration3948 specparam_declaration_instance3948();
    specparam_declaration3949 specparam_declaration_instance3949();
    specparam_declaration3950 specparam_declaration_instance3950();
    specparam_declaration3951 specparam_declaration_instance3951();
    specparam_declaration3952 specparam_declaration_instance3952();
    specparam_declaration3953 specparam_declaration_instance3953();
    specparam_declaration3954 specparam_declaration_instance3954();
    specparam_declaration3955 specparam_declaration_instance3955();
    specparam_declaration3956 specparam_declaration_instance3956();
    specparam_declaration3957 specparam_declaration_instance3957();
    specparam_declaration3958 specparam_declaration_instance3958();
    specparam_declaration3959 specparam_declaration_instance3959();
    specparam_declaration3960 specparam_declaration_instance3960();
    specparam_declaration3961 specparam_declaration_instance3961();
    specparam_declaration3962 specparam_declaration_instance3962();
    specparam_declaration3963 specparam_declaration_instance3963();
    specparam_declaration3964 specparam_declaration_instance3964();
    specparam_declaration3965 specparam_declaration_instance3965();
    specparam_declaration3966 specparam_declaration_instance3966();
    specparam_declaration3967 specparam_declaration_instance3967();
    specparam_declaration3968 specparam_declaration_instance3968();
    specparam_declaration3969 specparam_declaration_instance3969();
    specparam_declaration3970 specparam_declaration_instance3970();
    specparam_declaration3971 specparam_declaration_instance3971();
    specparam_declaration3972 specparam_declaration_instance3972();
    specparam_declaration3973 specparam_declaration_instance3973();
    specparam_declaration3974 specparam_declaration_instance3974();
    specparam_declaration3975 specparam_declaration_instance3975();
    specparam_declaration3976 specparam_declaration_instance3976();
    specparam_declaration3977 specparam_declaration_instance3977();
    specparam_declaration3978 specparam_declaration_instance3978();
    specparam_declaration3979 specparam_declaration_instance3979();
    specparam_declaration3980 specparam_declaration_instance3980();
    specparam_declaration3981 specparam_declaration_instance3981();
    specparam_declaration3982 specparam_declaration_instance3982();
    specparam_declaration3983 specparam_declaration_instance3983();
    specparam_declaration3984 specparam_declaration_instance3984();
    specparam_declaration3985 specparam_declaration_instance3985();
    specparam_declaration3986 specparam_declaration_instance3986();
    specparam_declaration3987 specparam_declaration_instance3987();
    specparam_declaration3988 specparam_declaration_instance3988();
    specparam_declaration3989 specparam_declaration_instance3989();
    specparam_declaration3990 specparam_declaration_instance3990();
    specparam_declaration3991 specparam_declaration_instance3991();
    specparam_declaration3992 specparam_declaration_instance3992();
    specparam_declaration3993 specparam_declaration_instance3993();
    specparam_declaration3994 specparam_declaration_instance3994();
    specparam_declaration3995 specparam_declaration_instance3995();
    specparam_declaration3996 specparam_declaration_instance3996();
    specparam_declaration3997 specparam_declaration_instance3997();
    specparam_declaration3998 specparam_declaration_instance3998();
    specparam_declaration3999 specparam_declaration_instance3999();
    specparam_declaration4000 specparam_declaration_instance4000();
    specparam_declaration4001 specparam_declaration_instance4001();
    specparam_declaration4002 specparam_declaration_instance4002();
    specparam_declaration4003 specparam_declaration_instance4003();
    specparam_declaration4004 specparam_declaration_instance4004();
    specparam_declaration4005 specparam_declaration_instance4005();
    specparam_declaration4006 specparam_declaration_instance4006();
    specparam_declaration4007 specparam_declaration_instance4007();
    specparam_declaration4008 specparam_declaration_instance4008();
    specparam_declaration4009 specparam_declaration_instance4009();
    specparam_declaration4010 specparam_declaration_instance4010();
    specparam_declaration4011 specparam_declaration_instance4011();
    specparam_declaration4012 specparam_declaration_instance4012();
    specparam_declaration4013 specparam_declaration_instance4013();
    specparam_declaration4014 specparam_declaration_instance4014();
    specparam_declaration4015 specparam_declaration_instance4015();
    specparam_declaration4016 specparam_declaration_instance4016();
    specparam_declaration4017 specparam_declaration_instance4017();
    specparam_declaration4018 specparam_declaration_instance4018();
    specparam_declaration4019 specparam_declaration_instance4019();
    specparam_declaration4020 specparam_declaration_instance4020();
    specparam_declaration4021 specparam_declaration_instance4021();
    specparam_declaration4022 specparam_declaration_instance4022();
    specparam_declaration4023 specparam_declaration_instance4023();
    specparam_declaration4024 specparam_declaration_instance4024();
    specparam_declaration4025 specparam_declaration_instance4025();
    specparam_declaration4026 specparam_declaration_instance4026();
    specparam_declaration4027 specparam_declaration_instance4027();
    specparam_declaration4028 specparam_declaration_instance4028();
    specparam_declaration4029 specparam_declaration_instance4029();
    specparam_declaration4030 specparam_declaration_instance4030();
    specparam_declaration4031 specparam_declaration_instance4031();
    specparam_declaration4032 specparam_declaration_instance4032();
    specparam_declaration4033 specparam_declaration_instance4033();
    specparam_declaration4034 specparam_declaration_instance4034();
    specparam_declaration4035 specparam_declaration_instance4035();
    specparam_declaration4036 specparam_declaration_instance4036();
    specparam_declaration4037 specparam_declaration_instance4037();
    specparam_declaration4038 specparam_declaration_instance4038();
    specparam_declaration4039 specparam_declaration_instance4039();
    specparam_declaration4040 specparam_declaration_instance4040();
    specparam_declaration4041 specparam_declaration_instance4041();
    specparam_declaration4042 specparam_declaration_instance4042();
    specparam_declaration4043 specparam_declaration_instance4043();
    specparam_declaration4044 specparam_declaration_instance4044();
    specparam_declaration4045 specparam_declaration_instance4045();
    specparam_declaration4046 specparam_declaration_instance4046();
    specparam_declaration4047 specparam_declaration_instance4047();
    specparam_declaration4048 specparam_declaration_instance4048();
    specparam_declaration4049 specparam_declaration_instance4049();
    specparam_declaration4050 specparam_declaration_instance4050();
    specparam_declaration4051 specparam_declaration_instance4051();
    specparam_declaration4052 specparam_declaration_instance4052();
    specparam_declaration4053 specparam_declaration_instance4053();
    specparam_declaration4054 specparam_declaration_instance4054();
    specparam_declaration4055 specparam_declaration_instance4055();
    specparam_declaration4056 specparam_declaration_instance4056();
    specparam_declaration4057 specparam_declaration_instance4057();
    specparam_declaration4058 specparam_declaration_instance4058();
    specparam_declaration4059 specparam_declaration_instance4059();
    specparam_declaration4060 specparam_declaration_instance4060();
    specparam_declaration4061 specparam_declaration_instance4061();
    specparam_declaration4062 specparam_declaration_instance4062();
    specparam_declaration4063 specparam_declaration_instance4063();
    specparam_declaration4064 specparam_declaration_instance4064();
    specparam_declaration4065 specparam_declaration_instance4065();
    specparam_declaration4066 specparam_declaration_instance4066();
    specparam_declaration4067 specparam_declaration_instance4067();
    specparam_declaration4068 specparam_declaration_instance4068();
    specparam_declaration4069 specparam_declaration_instance4069();
    specparam_declaration4070 specparam_declaration_instance4070();
    specparam_declaration4071 specparam_declaration_instance4071();
    specparam_declaration4072 specparam_declaration_instance4072();
    specparam_declaration4073 specparam_declaration_instance4073();
    specparam_declaration4074 specparam_declaration_instance4074();
    specparam_declaration4075 specparam_declaration_instance4075();
    specparam_declaration4076 specparam_declaration_instance4076();
    specparam_declaration4077 specparam_declaration_instance4077();
    specparam_declaration4078 specparam_declaration_instance4078();
    specparam_declaration4079 specparam_declaration_instance4079();
    specparam_declaration4080 specparam_declaration_instance4080();
    specparam_declaration4081 specparam_declaration_instance4081();
    specparam_declaration4082 specparam_declaration_instance4082();
    specparam_declaration4083 specparam_declaration_instance4083();
    specparam_declaration4084 specparam_declaration_instance4084();
    specparam_declaration4085 specparam_declaration_instance4085();
    specparam_declaration4086 specparam_declaration_instance4086();
    specparam_declaration4087 specparam_declaration_instance4087();
    specparam_declaration4088 specparam_declaration_instance4088();
    specparam_declaration4089 specparam_declaration_instance4089();
    specparam_declaration4090 specparam_declaration_instance4090();
    specparam_declaration4091 specparam_declaration_instance4091();
    specparam_declaration4092 specparam_declaration_instance4092();
    specparam_declaration4093 specparam_declaration_instance4093();
    specparam_declaration4094 specparam_declaration_instance4094();
    specparam_declaration4095 specparam_declaration_instance4095();
    specparam_declaration4096 specparam_declaration_instance4096();
    specparam_declaration4097 specparam_declaration_instance4097();
    specparam_declaration4098 specparam_declaration_instance4098();
    specparam_declaration4099 specparam_declaration_instance4099();
    specparam_declaration4100 specparam_declaration_instance4100();
    specparam_declaration4101 specparam_declaration_instance4101();
    specparam_declaration4102 specparam_declaration_instance4102();
    specparam_declaration4103 specparam_declaration_instance4103();
    specparam_declaration4104 specparam_declaration_instance4104();
    specparam_declaration4105 specparam_declaration_instance4105();
    specparam_declaration4106 specparam_declaration_instance4106();
    specparam_declaration4107 specparam_declaration_instance4107();
    specparam_declaration4108 specparam_declaration_instance4108();
    specparam_declaration4109 specparam_declaration_instance4109();
    specparam_declaration4110 specparam_declaration_instance4110();
    specparam_declaration4111 specparam_declaration_instance4111();
    specparam_declaration4112 specparam_declaration_instance4112();
    specparam_declaration4113 specparam_declaration_instance4113();
    specparam_declaration4114 specparam_declaration_instance4114();
    specparam_declaration4115 specparam_declaration_instance4115();
    specparam_declaration4116 specparam_declaration_instance4116();
    specparam_declaration4117 specparam_declaration_instance4117();
    specparam_declaration4118 specparam_declaration_instance4118();
    specparam_declaration4119 specparam_declaration_instance4119();
    specparam_declaration4120 specparam_declaration_instance4120();
    specparam_declaration4121 specparam_declaration_instance4121();
    specparam_declaration4122 specparam_declaration_instance4122();
    specparam_declaration4123 specparam_declaration_instance4123();
    specparam_declaration4124 specparam_declaration_instance4124();
    specparam_declaration4125 specparam_declaration_instance4125();
    specparam_declaration4126 specparam_declaration_instance4126();
    specparam_declaration4127 specparam_declaration_instance4127();
    specparam_declaration4128 specparam_declaration_instance4128();
    specparam_declaration4129 specparam_declaration_instance4129();
    specparam_declaration4130 specparam_declaration_instance4130();
    specparam_declaration4131 specparam_declaration_instance4131();
    specparam_declaration4132 specparam_declaration_instance4132();
    specparam_declaration4133 specparam_declaration_instance4133();
    specparam_declaration4134 specparam_declaration_instance4134();
    specparam_declaration4135 specparam_declaration_instance4135();
    specparam_declaration4136 specparam_declaration_instance4136();
    specparam_declaration4137 specparam_declaration_instance4137();
    specparam_declaration4138 specparam_declaration_instance4138();
    specparam_declaration4139 specparam_declaration_instance4139();
    specparam_declaration4140 specparam_declaration_instance4140();
    specparam_declaration4141 specparam_declaration_instance4141();
    specparam_declaration4142 specparam_declaration_instance4142();
    specparam_declaration4143 specparam_declaration_instance4143();
    specparam_declaration4144 specparam_declaration_instance4144();
    specparam_declaration4145 specparam_declaration_instance4145();
    specparam_declaration4146 specparam_declaration_instance4146();
    specparam_declaration4147 specparam_declaration_instance4147();
    specparam_declaration4148 specparam_declaration_instance4148();
    specparam_declaration4149 specparam_declaration_instance4149();
    specparam_declaration4150 specparam_declaration_instance4150();
    specparam_declaration4151 specparam_declaration_instance4151();
    specparam_declaration4152 specparam_declaration_instance4152();
    specparam_declaration4153 specparam_declaration_instance4153();
    specparam_declaration4154 specparam_declaration_instance4154();
    specparam_declaration4155 specparam_declaration_instance4155();
    specparam_declaration4156 specparam_declaration_instance4156();
    specparam_declaration4157 specparam_declaration_instance4157();
    specparam_declaration4158 specparam_declaration_instance4158();
    specparam_declaration4159 specparam_declaration_instance4159();
    specparam_declaration4160 specparam_declaration_instance4160();
    specparam_declaration4161 specparam_declaration_instance4161();
    specparam_declaration4162 specparam_declaration_instance4162();
    specparam_declaration4163 specparam_declaration_instance4163();
    specparam_declaration4164 specparam_declaration_instance4164();
    specparam_declaration4165 specparam_declaration_instance4165();
    specparam_declaration4166 specparam_declaration_instance4166();
    specparam_declaration4167 specparam_declaration_instance4167();
    specparam_declaration4168 specparam_declaration_instance4168();
    specparam_declaration4169 specparam_declaration_instance4169();
    specparam_declaration4170 specparam_declaration_instance4170();
    specparam_declaration4171 specparam_declaration_instance4171();
    specparam_declaration4172 specparam_declaration_instance4172();
    specparam_declaration4173 specparam_declaration_instance4173();
    specparam_declaration4174 specparam_declaration_instance4174();
    specparam_declaration4175 specparam_declaration_instance4175();
    specparam_declaration4176 specparam_declaration_instance4176();
    specparam_declaration4177 specparam_declaration_instance4177();
    specparam_declaration4178 specparam_declaration_instance4178();
    specparam_declaration4179 specparam_declaration_instance4179();
    specparam_declaration4180 specparam_declaration_instance4180();
    specparam_declaration4181 specparam_declaration_instance4181();
    specparam_declaration4182 specparam_declaration_instance4182();
    specparam_declaration4183 specparam_declaration_instance4183();
    specparam_declaration4184 specparam_declaration_instance4184();
    specparam_declaration4185 specparam_declaration_instance4185();
    specparam_declaration4186 specparam_declaration_instance4186();
    specparam_declaration4187 specparam_declaration_instance4187();
    specparam_declaration4188 specparam_declaration_instance4188();
    specparam_declaration4189 specparam_declaration_instance4189();
    specparam_declaration4190 specparam_declaration_instance4190();
    specparam_declaration4191 specparam_declaration_instance4191();
    specparam_declaration4192 specparam_declaration_instance4192();
    specparam_declaration4193 specparam_declaration_instance4193();
    specparam_declaration4194 specparam_declaration_instance4194();
    specparam_declaration4195 specparam_declaration_instance4195();
    specparam_declaration4196 specparam_declaration_instance4196();
    specparam_declaration4197 specparam_declaration_instance4197();
    specparam_declaration4198 specparam_declaration_instance4198();
    specparam_declaration4199 specparam_declaration_instance4199();
    specparam_declaration4200 specparam_declaration_instance4200();
    specparam_declaration4201 specparam_declaration_instance4201();
    specparam_declaration4202 specparam_declaration_instance4202();
    specparam_declaration4203 specparam_declaration_instance4203();
    specparam_declaration4204 specparam_declaration_instance4204();
    specparam_declaration4205 specparam_declaration_instance4205();
    specparam_declaration4206 specparam_declaration_instance4206();
    specparam_declaration4207 specparam_declaration_instance4207();
    specparam_declaration4208 specparam_declaration_instance4208();
    specparam_declaration4209 specparam_declaration_instance4209();
    specparam_declaration4210 specparam_declaration_instance4210();
    specparam_declaration4211 specparam_declaration_instance4211();
    specparam_declaration4212 specparam_declaration_instance4212();
    specparam_declaration4213 specparam_declaration_instance4213();
    specparam_declaration4214 specparam_declaration_instance4214();
    specparam_declaration4215 specparam_declaration_instance4215();
    specparam_declaration4216 specparam_declaration_instance4216();
    specparam_declaration4217 specparam_declaration_instance4217();
    specparam_declaration4218 specparam_declaration_instance4218();
    specparam_declaration4219 specparam_declaration_instance4219();
    specparam_declaration4220 specparam_declaration_instance4220();
    specparam_declaration4221 specparam_declaration_instance4221();
    specparam_declaration4222 specparam_declaration_instance4222();
    specparam_declaration4223 specparam_declaration_instance4223();
    specparam_declaration4224 specparam_declaration_instance4224();
    specparam_declaration4225 specparam_declaration_instance4225();
    specparam_declaration4226 specparam_declaration_instance4226();
    specparam_declaration4227 specparam_declaration_instance4227();
    specparam_declaration4228 specparam_declaration_instance4228();
    specparam_declaration4229 specparam_declaration_instance4229();
    specparam_declaration4230 specparam_declaration_instance4230();
    specparam_declaration4231 specparam_declaration_instance4231();
    specparam_declaration4232 specparam_declaration_instance4232();
    specparam_declaration4233 specparam_declaration_instance4233();
    specparam_declaration4234 specparam_declaration_instance4234();
    specparam_declaration4235 specparam_declaration_instance4235();
    specparam_declaration4236 specparam_declaration_instance4236();
    specparam_declaration4237 specparam_declaration_instance4237();
    specparam_declaration4238 specparam_declaration_instance4238();
    specparam_declaration4239 specparam_declaration_instance4239();
    specparam_declaration4240 specparam_declaration_instance4240();
    specparam_declaration4241 specparam_declaration_instance4241();
    specparam_declaration4242 specparam_declaration_instance4242();
    specparam_declaration4243 specparam_declaration_instance4243();
    specparam_declaration4244 specparam_declaration_instance4244();
    specparam_declaration4245 specparam_declaration_instance4245();
    specparam_declaration4246 specparam_declaration_instance4246();
    specparam_declaration4247 specparam_declaration_instance4247();
    specparam_declaration4248 specparam_declaration_instance4248();
    specparam_declaration4249 specparam_declaration_instance4249();
    specparam_declaration4250 specparam_declaration_instance4250();
    specparam_declaration4251 specparam_declaration_instance4251();
    specparam_declaration4252 specparam_declaration_instance4252();
    specparam_declaration4253 specparam_declaration_instance4253();
    specparam_declaration4254 specparam_declaration_instance4254();
    specparam_declaration4255 specparam_declaration_instance4255();
    specparam_declaration4256 specparam_declaration_instance4256();
    specparam_declaration4257 specparam_declaration_instance4257();
    specparam_declaration4258 specparam_declaration_instance4258();
    specparam_declaration4259 specparam_declaration_instance4259();
    specparam_declaration4260 specparam_declaration_instance4260();
    specparam_declaration4261 specparam_declaration_instance4261();
    specparam_declaration4262 specparam_declaration_instance4262();
    specparam_declaration4263 specparam_declaration_instance4263();
    specparam_declaration4264 specparam_declaration_instance4264();
    specparam_declaration4265 specparam_declaration_instance4265();
    specparam_declaration4266 specparam_declaration_instance4266();
    specparam_declaration4267 specparam_declaration_instance4267();
    specparam_declaration4268 specparam_declaration_instance4268();
    specparam_declaration4269 specparam_declaration_instance4269();
    specparam_declaration4270 specparam_declaration_instance4270();
    specparam_declaration4271 specparam_declaration_instance4271();
    specparam_declaration4272 specparam_declaration_instance4272();
    specparam_declaration4273 specparam_declaration_instance4273();
    specparam_declaration4274 specparam_declaration_instance4274();
    specparam_declaration4275 specparam_declaration_instance4275();
    specparam_declaration4276 specparam_declaration_instance4276();
    specparam_declaration4277 specparam_declaration_instance4277();
    specparam_declaration4278 specparam_declaration_instance4278();
    specparam_declaration4279 specparam_declaration_instance4279();
    specparam_declaration4280 specparam_declaration_instance4280();
    specparam_declaration4281 specparam_declaration_instance4281();
    specparam_declaration4282 specparam_declaration_instance4282();
    specparam_declaration4283 specparam_declaration_instance4283();
    specparam_declaration4284 specparam_declaration_instance4284();
    specparam_declaration4285 specparam_declaration_instance4285();
    specparam_declaration4286 specparam_declaration_instance4286();
    specparam_declaration4287 specparam_declaration_instance4287();
    specparam_declaration4288 specparam_declaration_instance4288();
    specparam_declaration4289 specparam_declaration_instance4289();
    specparam_declaration4290 specparam_declaration_instance4290();
    specparam_declaration4291 specparam_declaration_instance4291();
    specparam_declaration4292 specparam_declaration_instance4292();
    specparam_declaration4293 specparam_declaration_instance4293();
    specparam_declaration4294 specparam_declaration_instance4294();
    specparam_declaration4295 specparam_declaration_instance4295();
    specparam_declaration4296 specparam_declaration_instance4296();
    specparam_declaration4297 specparam_declaration_instance4297();
    specparam_declaration4298 specparam_declaration_instance4298();
    specparam_declaration4299 specparam_declaration_instance4299();
    specparam_declaration4300 specparam_declaration_instance4300();
    specparam_declaration4301 specparam_declaration_instance4301();
    specparam_declaration4302 specparam_declaration_instance4302();
    specparam_declaration4303 specparam_declaration_instance4303();
    specparam_declaration4304 specparam_declaration_instance4304();
    specparam_declaration4305 specparam_declaration_instance4305();
    specparam_declaration4306 specparam_declaration_instance4306();
    specparam_declaration4307 specparam_declaration_instance4307();
    specparam_declaration4308 specparam_declaration_instance4308();
    specparam_declaration4309 specparam_declaration_instance4309();
    specparam_declaration4310 specparam_declaration_instance4310();
    specparam_declaration4311 specparam_declaration_instance4311();
    specparam_declaration4312 specparam_declaration_instance4312();
    specparam_declaration4313 specparam_declaration_instance4313();
    specparam_declaration4314 specparam_declaration_instance4314();
    specparam_declaration4315 specparam_declaration_instance4315();
    specparam_declaration4316 specparam_declaration_instance4316();
    specparam_declaration4317 specparam_declaration_instance4317();
    specparam_declaration4318 specparam_declaration_instance4318();
    specparam_declaration4319 specparam_declaration_instance4319();
    specparam_declaration4320 specparam_declaration_instance4320();
    specparam_declaration4321 specparam_declaration_instance4321();
    specparam_declaration4322 specparam_declaration_instance4322();
    specparam_declaration4323 specparam_declaration_instance4323();
    specparam_declaration4324 specparam_declaration_instance4324();
    specparam_declaration4325 specparam_declaration_instance4325();
    specparam_declaration4326 specparam_declaration_instance4326();
    specparam_declaration4327 specparam_declaration_instance4327();
    specparam_declaration4328 specparam_declaration_instance4328();
    specparam_declaration4329 specparam_declaration_instance4329();
    specparam_declaration4330 specparam_declaration_instance4330();
    specparam_declaration4331 specparam_declaration_instance4331();
    specparam_declaration4332 specparam_declaration_instance4332();
    specparam_declaration4333 specparam_declaration_instance4333();
    specparam_declaration4334 specparam_declaration_instance4334();
    specparam_declaration4335 specparam_declaration_instance4335();
    specparam_declaration4336 specparam_declaration_instance4336();
    specparam_declaration4337 specparam_declaration_instance4337();
    specparam_declaration4338 specparam_declaration_instance4338();
    specparam_declaration4339 specparam_declaration_instance4339();
    specparam_declaration4340 specparam_declaration_instance4340();
    specparam_declaration4341 specparam_declaration_instance4341();
    specparam_declaration4342 specparam_declaration_instance4342();
    specparam_declaration4343 specparam_declaration_instance4343();
    specparam_declaration4344 specparam_declaration_instance4344();
    specparam_declaration4345 specparam_declaration_instance4345();
    specparam_declaration4346 specparam_declaration_instance4346();
    specparam_declaration4347 specparam_declaration_instance4347();
    specparam_declaration4348 specparam_declaration_instance4348();
    specparam_declaration4349 specparam_declaration_instance4349();
    specparam_declaration4350 specparam_declaration_instance4350();
    specparam_declaration4351 specparam_declaration_instance4351();
    specparam_declaration4352 specparam_declaration_instance4352();
    specparam_declaration4353 specparam_declaration_instance4353();
    specparam_declaration4354 specparam_declaration_instance4354();
    specparam_declaration4355 specparam_declaration_instance4355();
    specparam_declaration4356 specparam_declaration_instance4356();
    specparam_declaration4357 specparam_declaration_instance4357();
    specparam_declaration4358 specparam_declaration_instance4358();
    specparam_declaration4359 specparam_declaration_instance4359();
    specparam_declaration4360 specparam_declaration_instance4360();
    specparam_declaration4361 specparam_declaration_instance4361();
    specparam_declaration4362 specparam_declaration_instance4362();
    specparam_declaration4363 specparam_declaration_instance4363();
    specparam_declaration4364 specparam_declaration_instance4364();
    specparam_declaration4365 specparam_declaration_instance4365();
    specparam_declaration4366 specparam_declaration_instance4366();
    specparam_declaration4367 specparam_declaration_instance4367();
    specparam_declaration4368 specparam_declaration_instance4368();
    specparam_declaration4369 specparam_declaration_instance4369();
    specparam_declaration4370 specparam_declaration_instance4370();
    specparam_declaration4371 specparam_declaration_instance4371();
    specparam_declaration4372 specparam_declaration_instance4372();
    specparam_declaration4373 specparam_declaration_instance4373();
    specparam_declaration4374 specparam_declaration_instance4374();
    specparam_declaration4375 specparam_declaration_instance4375();
    specparam_declaration4376 specparam_declaration_instance4376();
    specparam_declaration4377 specparam_declaration_instance4377();
    specparam_declaration4378 specparam_declaration_instance4378();
    specparam_declaration4379 specparam_declaration_instance4379();
    specparam_declaration4380 specparam_declaration_instance4380();
    specparam_declaration4381 specparam_declaration_instance4381();
    specparam_declaration4382 specparam_declaration_instance4382();
    specparam_declaration4383 specparam_declaration_instance4383();
    specparam_declaration4384 specparam_declaration_instance4384();
    specparam_declaration4385 specparam_declaration_instance4385();
    specparam_declaration4386 specparam_declaration_instance4386();
    specparam_declaration4387 specparam_declaration_instance4387();
    specparam_declaration4388 specparam_declaration_instance4388();
    specparam_declaration4389 specparam_declaration_instance4389();
    specparam_declaration4390 specparam_declaration_instance4390();
    specparam_declaration4391 specparam_declaration_instance4391();
    specparam_declaration4392 specparam_declaration_instance4392();
    specparam_declaration4393 specparam_declaration_instance4393();
    specparam_declaration4394 specparam_declaration_instance4394();
    specparam_declaration4395 specparam_declaration_instance4395();
    specparam_declaration4396 specparam_declaration_instance4396();
    specparam_declaration4397 specparam_declaration_instance4397();
    specparam_declaration4398 specparam_declaration_instance4398();
    specparam_declaration4399 specparam_declaration_instance4399();
    specparam_declaration4400 specparam_declaration_instance4400();
    specparam_declaration4401 specparam_declaration_instance4401();
    specparam_declaration4402 specparam_declaration_instance4402();
    specparam_declaration4403 specparam_declaration_instance4403();
    specparam_declaration4404 specparam_declaration_instance4404();
    specparam_declaration4405 specparam_declaration_instance4405();
    specparam_declaration4406 specparam_declaration_instance4406();
    specparam_declaration4407 specparam_declaration_instance4407();
    specparam_declaration4408 specparam_declaration_instance4408();
    specparam_declaration4409 specparam_declaration_instance4409();
    specparam_declaration4410 specparam_declaration_instance4410();
    specparam_declaration4411 specparam_declaration_instance4411();
    specparam_declaration4412 specparam_declaration_instance4412();
    specparam_declaration4413 specparam_declaration_instance4413();
    specparam_declaration4414 specparam_declaration_instance4414();
    specparam_declaration4415 specparam_declaration_instance4415();
    specparam_declaration4416 specparam_declaration_instance4416();
    specparam_declaration4417 specparam_declaration_instance4417();
    specparam_declaration4418 specparam_declaration_instance4418();
    specparam_declaration4419 specparam_declaration_instance4419();
    specparam_declaration4420 specparam_declaration_instance4420();
    specparam_declaration4421 specparam_declaration_instance4421();
    specparam_declaration4422 specparam_declaration_instance4422();
    specparam_declaration4423 specparam_declaration_instance4423();
    specparam_declaration4424 specparam_declaration_instance4424();
    specparam_declaration4425 specparam_declaration_instance4425();
    specparam_declaration4426 specparam_declaration_instance4426();
    specparam_declaration4427 specparam_declaration_instance4427();
    specparam_declaration4428 specparam_declaration_instance4428();
    specparam_declaration4429 specparam_declaration_instance4429();
    specparam_declaration4430 specparam_declaration_instance4430();
    specparam_declaration4431 specparam_declaration_instance4431();
    specparam_declaration4432 specparam_declaration_instance4432();
    specparam_declaration4433 specparam_declaration_instance4433();
    specparam_declaration4434 specparam_declaration_instance4434();
    specparam_declaration4435 specparam_declaration_instance4435();
    specparam_declaration4436 specparam_declaration_instance4436();
    specparam_declaration4437 specparam_declaration_instance4437();
    specparam_declaration4438 specparam_declaration_instance4438();
    specparam_declaration4439 specparam_declaration_instance4439();
    specparam_declaration4440 specparam_declaration_instance4440();
    specparam_declaration4441 specparam_declaration_instance4441();
    specparam_declaration4442 specparam_declaration_instance4442();
    specparam_declaration4443 specparam_declaration_instance4443();
    specparam_declaration4444 specparam_declaration_instance4444();
    specparam_declaration4445 specparam_declaration_instance4445();
    specparam_declaration4446 specparam_declaration_instance4446();
    specparam_declaration4447 specparam_declaration_instance4447();
    specparam_declaration4448 specparam_declaration_instance4448();
    specparam_declaration4449 specparam_declaration_instance4449();
    specparam_declaration4450 specparam_declaration_instance4450();
    specparam_declaration4451 specparam_declaration_instance4451();
    specparam_declaration4452 specparam_declaration_instance4452();
    specparam_declaration4453 specparam_declaration_instance4453();
    specparam_declaration4454 specparam_declaration_instance4454();
    specparam_declaration4455 specparam_declaration_instance4455();
    specparam_declaration4456 specparam_declaration_instance4456();
    specparam_declaration4457 specparam_declaration_instance4457();
    specparam_declaration4458 specparam_declaration_instance4458();
    specparam_declaration4459 specparam_declaration_instance4459();
    specparam_declaration4460 specparam_declaration_instance4460();
    specparam_declaration4461 specparam_declaration_instance4461();
    specparam_declaration4462 specparam_declaration_instance4462();
    specparam_declaration4463 specparam_declaration_instance4463();
    specparam_declaration4464 specparam_declaration_instance4464();
    specparam_declaration4465 specparam_declaration_instance4465();
    specparam_declaration4466 specparam_declaration_instance4466();
    specparam_declaration4467 specparam_declaration_instance4467();
    specparam_declaration4468 specparam_declaration_instance4468();
    specparam_declaration4469 specparam_declaration_instance4469();
    specparam_declaration4470 specparam_declaration_instance4470();
    specparam_declaration4471 specparam_declaration_instance4471();
    specparam_declaration4472 specparam_declaration_instance4472();
    specparam_declaration4473 specparam_declaration_instance4473();
    specparam_declaration4474 specparam_declaration_instance4474();
    specparam_declaration4475 specparam_declaration_instance4475();
    specparam_declaration4476 specparam_declaration_instance4476();
    specparam_declaration4477 specparam_declaration_instance4477();
    specparam_declaration4478 specparam_declaration_instance4478();
    specparam_declaration4479 specparam_declaration_instance4479();
    specparam_declaration4480 specparam_declaration_instance4480();
    specparam_declaration4481 specparam_declaration_instance4481();
    specparam_declaration4482 specparam_declaration_instance4482();
    specparam_declaration4483 specparam_declaration_instance4483();
    specparam_declaration4484 specparam_declaration_instance4484();
    specparam_declaration4485 specparam_declaration_instance4485();
    specparam_declaration4486 specparam_declaration_instance4486();
    specparam_declaration4487 specparam_declaration_instance4487();
    specparam_declaration4488 specparam_declaration_instance4488();
    specparam_declaration4489 specparam_declaration_instance4489();
    specparam_declaration4490 specparam_declaration_instance4490();
    specparam_declaration4491 specparam_declaration_instance4491();
    specparam_declaration4492 specparam_declaration_instance4492();
    specparam_declaration4493 specparam_declaration_instance4493();
    specparam_declaration4494 specparam_declaration_instance4494();
    specparam_declaration4495 specparam_declaration_instance4495();
    specparam_declaration4496 specparam_declaration_instance4496();
    specparam_declaration4497 specparam_declaration_instance4497();
    specparam_declaration4498 specparam_declaration_instance4498();
    specparam_declaration4499 specparam_declaration_instance4499();
    specparam_declaration4500 specparam_declaration_instance4500();
    specparam_declaration4501 specparam_declaration_instance4501();
    specparam_declaration4502 specparam_declaration_instance4502();
    specparam_declaration4503 specparam_declaration_instance4503();
    specparam_declaration4504 specparam_declaration_instance4504();
    specparam_declaration4505 specparam_declaration_instance4505();
    specparam_declaration4506 specparam_declaration_instance4506();
    specparam_declaration4507 specparam_declaration_instance4507();
    specparam_declaration4508 specparam_declaration_instance4508();
    specparam_declaration4509 specparam_declaration_instance4509();
    specparam_declaration4510 specparam_declaration_instance4510();
    specparam_declaration4511 specparam_declaration_instance4511();
    specparam_declaration4512 specparam_declaration_instance4512();
    specparam_declaration4513 specparam_declaration_instance4513();
    specparam_declaration4514 specparam_declaration_instance4514();
    specparam_declaration4515 specparam_declaration_instance4515();
    specparam_declaration4516 specparam_declaration_instance4516();
    specparam_declaration4517 specparam_declaration_instance4517();
    specparam_declaration4518 specparam_declaration_instance4518();
    specparam_declaration4519 specparam_declaration_instance4519();
    specparam_declaration4520 specparam_declaration_instance4520();
    specparam_declaration4521 specparam_declaration_instance4521();
    specparam_declaration4522 specparam_declaration_instance4522();
    specparam_declaration4523 specparam_declaration_instance4523();
    specparam_declaration4524 specparam_declaration_instance4524();
    specparam_declaration4525 specparam_declaration_instance4525();
    specparam_declaration4526 specparam_declaration_instance4526();
    specparam_declaration4527 specparam_declaration_instance4527();
    specparam_declaration4528 specparam_declaration_instance4528();
    specparam_declaration4529 specparam_declaration_instance4529();
    specparam_declaration4530 specparam_declaration_instance4530();
    specparam_declaration4531 specparam_declaration_instance4531();
    specparam_declaration4532 specparam_declaration_instance4532();
    specparam_declaration4533 specparam_declaration_instance4533();
    specparam_declaration4534 specparam_declaration_instance4534();
    specparam_declaration4535 specparam_declaration_instance4535();
    specparam_declaration4536 specparam_declaration_instance4536();
    specparam_declaration4537 specparam_declaration_instance4537();
    specparam_declaration4538 specparam_declaration_instance4538();
    specparam_declaration4539 specparam_declaration_instance4539();
    specparam_declaration4540 specparam_declaration_instance4540();
    specparam_declaration4541 specparam_declaration_instance4541();
    specparam_declaration4542 specparam_declaration_instance4542();
    specparam_declaration4543 specparam_declaration_instance4543();
    specparam_declaration4544 specparam_declaration_instance4544();
    specparam_declaration4545 specparam_declaration_instance4545();
    specparam_declaration4546 specparam_declaration_instance4546();
    specparam_declaration4547 specparam_declaration_instance4547();
    specparam_declaration4548 specparam_declaration_instance4548();
    specparam_declaration4549 specparam_declaration_instance4549();
    specparam_declaration4550 specparam_declaration_instance4550();
    specparam_declaration4551 specparam_declaration_instance4551();
    specparam_declaration4552 specparam_declaration_instance4552();
    specparam_declaration4553 specparam_declaration_instance4553();
    specparam_declaration4554 specparam_declaration_instance4554();
    specparam_declaration4555 specparam_declaration_instance4555();
    specparam_declaration4556 specparam_declaration_instance4556();
    specparam_declaration4557 specparam_declaration_instance4557();
    specparam_declaration4558 specparam_declaration_instance4558();
    specparam_declaration4559 specparam_declaration_instance4559();
    specparam_declaration4560 specparam_declaration_instance4560();
    specparam_declaration4561 specparam_declaration_instance4561();
    specparam_declaration4562 specparam_declaration_instance4562();
    specparam_declaration4563 specparam_declaration_instance4563();
    specparam_declaration4564 specparam_declaration_instance4564();
    specparam_declaration4565 specparam_declaration_instance4565();
    specparam_declaration4566 specparam_declaration_instance4566();
    specparam_declaration4567 specparam_declaration_instance4567();
    specparam_declaration4568 specparam_declaration_instance4568();
    specparam_declaration4569 specparam_declaration_instance4569();
    specparam_declaration4570 specparam_declaration_instance4570();
    specparam_declaration4571 specparam_declaration_instance4571();
    specparam_declaration4572 specparam_declaration_instance4572();
    specparam_declaration4573 specparam_declaration_instance4573();
    specparam_declaration4574 specparam_declaration_instance4574();
    specparam_declaration4575 specparam_declaration_instance4575();
    specparam_declaration4576 specparam_declaration_instance4576();
    specparam_declaration4577 specparam_declaration_instance4577();
    specparam_declaration4578 specparam_declaration_instance4578();
    specparam_declaration4579 specparam_declaration_instance4579();
    specparam_declaration4580 specparam_declaration_instance4580();
    specparam_declaration4581 specparam_declaration_instance4581();
    specparam_declaration4582 specparam_declaration_instance4582();
    specparam_declaration4583 specparam_declaration_instance4583();
    specparam_declaration4584 specparam_declaration_instance4584();
    specparam_declaration4585 specparam_declaration_instance4585();
    specparam_declaration4586 specparam_declaration_instance4586();
    specparam_declaration4587 specparam_declaration_instance4587();
    specparam_declaration4588 specparam_declaration_instance4588();
    specparam_declaration4589 specparam_declaration_instance4589();
    specparam_declaration4590 specparam_declaration_instance4590();
    specparam_declaration4591 specparam_declaration_instance4591();
    specparam_declaration4592 specparam_declaration_instance4592();
    specparam_declaration4593 specparam_declaration_instance4593();
    specparam_declaration4594 specparam_declaration_instance4594();
    specparam_declaration4595 specparam_declaration_instance4595();
    specparam_declaration4596 specparam_declaration_instance4596();
    specparam_declaration4597 specparam_declaration_instance4597();
    specparam_declaration4598 specparam_declaration_instance4598();
    specparam_declaration4599 specparam_declaration_instance4599();
    specparam_declaration4600 specparam_declaration_instance4600();
    specparam_declaration4601 specparam_declaration_instance4601();
    specparam_declaration4602 specparam_declaration_instance4602();
    specparam_declaration4603 specparam_declaration_instance4603();
    specparam_declaration4604 specparam_declaration_instance4604();
    specparam_declaration4605 specparam_declaration_instance4605();
    specparam_declaration4606 specparam_declaration_instance4606();
    specparam_declaration4607 specparam_declaration_instance4607();
    specparam_declaration4608 specparam_declaration_instance4608();
    specparam_declaration4609 specparam_declaration_instance4609();
    specparam_declaration4610 specparam_declaration_instance4610();
    specparam_declaration4611 specparam_declaration_instance4611();
    specparam_declaration4612 specparam_declaration_instance4612();
    specparam_declaration4613 specparam_declaration_instance4613();
    specparam_declaration4614 specparam_declaration_instance4614();
    specparam_declaration4615 specparam_declaration_instance4615();
    specparam_declaration4616 specparam_declaration_instance4616();
    specparam_declaration4617 specparam_declaration_instance4617();
    specparam_declaration4618 specparam_declaration_instance4618();
    specparam_declaration4619 specparam_declaration_instance4619();
    specparam_declaration4620 specparam_declaration_instance4620();
    specparam_declaration4621 specparam_declaration_instance4621();
    specparam_declaration4622 specparam_declaration_instance4622();
    specparam_declaration4623 specparam_declaration_instance4623();
    specparam_declaration4624 specparam_declaration_instance4624();
    specparam_declaration4625 specparam_declaration_instance4625();
    specparam_declaration4626 specparam_declaration_instance4626();
    specparam_declaration4627 specparam_declaration_instance4627();
    specparam_declaration4628 specparam_declaration_instance4628();
    specparam_declaration4629 specparam_declaration_instance4629();
    specparam_declaration4630 specparam_declaration_instance4630();
    specparam_declaration4631 specparam_declaration_instance4631();
    specparam_declaration4632 specparam_declaration_instance4632();
    specparam_declaration4633 specparam_declaration_instance4633();
    specparam_declaration4634 specparam_declaration_instance4634();
    specparam_declaration4635 specparam_declaration_instance4635();
    specparam_declaration4636 specparam_declaration_instance4636();
    specparam_declaration4637 specparam_declaration_instance4637();
    specparam_declaration4638 specparam_declaration_instance4638();
    specparam_declaration4639 specparam_declaration_instance4639();
    specparam_declaration4640 specparam_declaration_instance4640();
    specparam_declaration4641 specparam_declaration_instance4641();
    specparam_declaration4642 specparam_declaration_instance4642();
    specparam_declaration4643 specparam_declaration_instance4643();
    specparam_declaration4644 specparam_declaration_instance4644();
    specparam_declaration4645 specparam_declaration_instance4645();
    specparam_declaration4646 specparam_declaration_instance4646();
    specparam_declaration4647 specparam_declaration_instance4647();
    specparam_declaration4648 specparam_declaration_instance4648();
    specparam_declaration4649 specparam_declaration_instance4649();
    specparam_declaration4650 specparam_declaration_instance4650();
    specparam_declaration4651 specparam_declaration_instance4651();
    specparam_declaration4652 specparam_declaration_instance4652();
    specparam_declaration4653 specparam_declaration_instance4653();
    specparam_declaration4654 specparam_declaration_instance4654();
    specparam_declaration4655 specparam_declaration_instance4655();
    specparam_declaration4656 specparam_declaration_instance4656();
    specparam_declaration4657 specparam_declaration_instance4657();
    specparam_declaration4658 specparam_declaration_instance4658();
    specparam_declaration4659 specparam_declaration_instance4659();
    specparam_declaration4660 specparam_declaration_instance4660();
    specparam_declaration4661 specparam_declaration_instance4661();
    specparam_declaration4662 specparam_declaration_instance4662();
    specparam_declaration4663 specparam_declaration_instance4663();
    specparam_declaration4664 specparam_declaration_instance4664();
    specparam_declaration4665 specparam_declaration_instance4665();
    specparam_declaration4666 specparam_declaration_instance4666();
    specparam_declaration4667 specparam_declaration_instance4667();
    specparam_declaration4668 specparam_declaration_instance4668();
    specparam_declaration4669 specparam_declaration_instance4669();
    specparam_declaration4670 specparam_declaration_instance4670();
    specparam_declaration4671 specparam_declaration_instance4671();
    specparam_declaration4672 specparam_declaration_instance4672();
    specparam_declaration4673 specparam_declaration_instance4673();
    specparam_declaration4674 specparam_declaration_instance4674();
    specparam_declaration4675 specparam_declaration_instance4675();
    specparam_declaration4676 specparam_declaration_instance4676();
    specparam_declaration4677 specparam_declaration_instance4677();
    specparam_declaration4678 specparam_declaration_instance4678();
    specparam_declaration4679 specparam_declaration_instance4679();
    specparam_declaration4680 specparam_declaration_instance4680();
    specparam_declaration4681 specparam_declaration_instance4681();
    specparam_declaration4682 specparam_declaration_instance4682();
    specparam_declaration4683 specparam_declaration_instance4683();
    specparam_declaration4684 specparam_declaration_instance4684();
    specparam_declaration4685 specparam_declaration_instance4685();
    specparam_declaration4686 specparam_declaration_instance4686();
    specparam_declaration4687 specparam_declaration_instance4687();
    specparam_declaration4688 specparam_declaration_instance4688();
    specparam_declaration4689 specparam_declaration_instance4689();
    specparam_declaration4690 specparam_declaration_instance4690();
    specparam_declaration4691 specparam_declaration_instance4691();
    specparam_declaration4692 specparam_declaration_instance4692();
    specparam_declaration4693 specparam_declaration_instance4693();
    specparam_declaration4694 specparam_declaration_instance4694();
    specparam_declaration4695 specparam_declaration_instance4695();
    specparam_declaration4696 specparam_declaration_instance4696();
    specparam_declaration4697 specparam_declaration_instance4697();
    specparam_declaration4698 specparam_declaration_instance4698();
    specparam_declaration4699 specparam_declaration_instance4699();
    specparam_declaration4700 specparam_declaration_instance4700();
    specparam_declaration4701 specparam_declaration_instance4701();
    specparam_declaration4702 specparam_declaration_instance4702();
    specparam_declaration4703 specparam_declaration_instance4703();
    specparam_declaration4704 specparam_declaration_instance4704();
    specparam_declaration4705 specparam_declaration_instance4705();
    specparam_declaration4706 specparam_declaration_instance4706();
    specparam_declaration4707 specparam_declaration_instance4707();
    specparam_declaration4708 specparam_declaration_instance4708();
    specparam_declaration4709 specparam_declaration_instance4709();
    specparam_declaration4710 specparam_declaration_instance4710();
    specparam_declaration4711 specparam_declaration_instance4711();
    specparam_declaration4712 specparam_declaration_instance4712();
    specparam_declaration4713 specparam_declaration_instance4713();
    specparam_declaration4714 specparam_declaration_instance4714();
    specparam_declaration4715 specparam_declaration_instance4715();
    specparam_declaration4716 specparam_declaration_instance4716();
    specparam_declaration4717 specparam_declaration_instance4717();
    specparam_declaration4718 specparam_declaration_instance4718();
    specparam_declaration4719 specparam_declaration_instance4719();
    specparam_declaration4720 specparam_declaration_instance4720();
    specparam_declaration4721 specparam_declaration_instance4721();
    specparam_declaration4722 specparam_declaration_instance4722();
    specparam_declaration4723 specparam_declaration_instance4723();
    specparam_declaration4724 specparam_declaration_instance4724();
    specparam_declaration4725 specparam_declaration_instance4725();
    specparam_declaration4726 specparam_declaration_instance4726();
    specparam_declaration4727 specparam_declaration_instance4727();
    specparam_declaration4728 specparam_declaration_instance4728();
    specparam_declaration4729 specparam_declaration_instance4729();
    specparam_declaration4730 specparam_declaration_instance4730();
    specparam_declaration4731 specparam_declaration_instance4731();
    specparam_declaration4732 specparam_declaration_instance4732();
    specparam_declaration4733 specparam_declaration_instance4733();
    specparam_declaration4734 specparam_declaration_instance4734();
    specparam_declaration4735 specparam_declaration_instance4735();
    specparam_declaration4736 specparam_declaration_instance4736();
    specparam_declaration4737 specparam_declaration_instance4737();
    specparam_declaration4738 specparam_declaration_instance4738();
    specparam_declaration4739 specparam_declaration_instance4739();
    specparam_declaration4740 specparam_declaration_instance4740();
    specparam_declaration4741 specparam_declaration_instance4741();
    specparam_declaration4742 specparam_declaration_instance4742();
    specparam_declaration4743 specparam_declaration_instance4743();
    specparam_declaration4744 specparam_declaration_instance4744();
    specparam_declaration4745 specparam_declaration_instance4745();
    specparam_declaration4746 specparam_declaration_instance4746();
    specparam_declaration4747 specparam_declaration_instance4747();
    specparam_declaration4748 specparam_declaration_instance4748();
    specparam_declaration4749 specparam_declaration_instance4749();
    specparam_declaration4750 specparam_declaration_instance4750();
    specparam_declaration4751 specparam_declaration_instance4751();
    specparam_declaration4752 specparam_declaration_instance4752();
    specparam_declaration4753 specparam_declaration_instance4753();
    specparam_declaration4754 specparam_declaration_instance4754();
    specparam_declaration4755 specparam_declaration_instance4755();
    specparam_declaration4756 specparam_declaration_instance4756();
    specparam_declaration4757 specparam_declaration_instance4757();
    specparam_declaration4758 specparam_declaration_instance4758();
    specparam_declaration4759 specparam_declaration_instance4759();
    specparam_declaration4760 specparam_declaration_instance4760();
    specparam_declaration4761 specparam_declaration_instance4761();
    specparam_declaration4762 specparam_declaration_instance4762();
    specparam_declaration4763 specparam_declaration_instance4763();
    specparam_declaration4764 specparam_declaration_instance4764();
    specparam_declaration4765 specparam_declaration_instance4765();
    specparam_declaration4766 specparam_declaration_instance4766();
    specparam_declaration4767 specparam_declaration_instance4767();
    specparam_declaration4768 specparam_declaration_instance4768();
    specparam_declaration4769 specparam_declaration_instance4769();
    specparam_declaration4770 specparam_declaration_instance4770();
    specparam_declaration4771 specparam_declaration_instance4771();
    specparam_declaration4772 specparam_declaration_instance4772();
    specparam_declaration4773 specparam_declaration_instance4773();
    specparam_declaration4774 specparam_declaration_instance4774();
    specparam_declaration4775 specparam_declaration_instance4775();
    specparam_declaration4776 specparam_declaration_instance4776();
    specparam_declaration4777 specparam_declaration_instance4777();
    specparam_declaration4778 specparam_declaration_instance4778();
    specparam_declaration4779 specparam_declaration_instance4779();
    specparam_declaration4780 specparam_declaration_instance4780();
    specparam_declaration4781 specparam_declaration_instance4781();
    specparam_declaration4782 specparam_declaration_instance4782();
    specparam_declaration4783 specparam_declaration_instance4783();
    specparam_declaration4784 specparam_declaration_instance4784();
    specparam_declaration4785 specparam_declaration_instance4785();
    specparam_declaration4786 specparam_declaration_instance4786();
    specparam_declaration4787 specparam_declaration_instance4787();
    specparam_declaration4788 specparam_declaration_instance4788();
    specparam_declaration4789 specparam_declaration_instance4789();
    specparam_declaration4790 specparam_declaration_instance4790();
    specparam_declaration4791 specparam_declaration_instance4791();
    specparam_declaration4792 specparam_declaration_instance4792();
    specparam_declaration4793 specparam_declaration_instance4793();
    specparam_declaration4794 specparam_declaration_instance4794();
    specparam_declaration4795 specparam_declaration_instance4795();
    specparam_declaration4796 specparam_declaration_instance4796();
    specparam_declaration4797 specparam_declaration_instance4797();
    specparam_declaration4798 specparam_declaration_instance4798();
    specparam_declaration4799 specparam_declaration_instance4799();
    specparam_declaration4800 specparam_declaration_instance4800();
    specparam_declaration4801 specparam_declaration_instance4801();
    specparam_declaration4802 specparam_declaration_instance4802();
    specparam_declaration4803 specparam_declaration_instance4803();
    specparam_declaration4804 specparam_declaration_instance4804();
    specparam_declaration4805 specparam_declaration_instance4805();
    specparam_declaration4806 specparam_declaration_instance4806();
    specparam_declaration4807 specparam_declaration_instance4807();
    specparam_declaration4808 specparam_declaration_instance4808();
    specparam_declaration4809 specparam_declaration_instance4809();
    specparam_declaration4810 specparam_declaration_instance4810();
    specparam_declaration4811 specparam_declaration_instance4811();
    specparam_declaration4812 specparam_declaration_instance4812();
    specparam_declaration4813 specparam_declaration_instance4813();
    specparam_declaration4814 specparam_declaration_instance4814();
    specparam_declaration4815 specparam_declaration_instance4815();
    specparam_declaration4816 specparam_declaration_instance4816();
    specparam_declaration4817 specparam_declaration_instance4817();
    specparam_declaration4818 specparam_declaration_instance4818();
    specparam_declaration4819 specparam_declaration_instance4819();
    specparam_declaration4820 specparam_declaration_instance4820();
    specparam_declaration4821 specparam_declaration_instance4821();
    specparam_declaration4822 specparam_declaration_instance4822();
    specparam_declaration4823 specparam_declaration_instance4823();
    specparam_declaration4824 specparam_declaration_instance4824();
    specparam_declaration4825 specparam_declaration_instance4825();
    specparam_declaration4826 specparam_declaration_instance4826();
    specparam_declaration4827 specparam_declaration_instance4827();
    specparam_declaration4828 specparam_declaration_instance4828();
    specparam_declaration4829 specparam_declaration_instance4829();
    specparam_declaration4830 specparam_declaration_instance4830();
    specparam_declaration4831 specparam_declaration_instance4831();
    specparam_declaration4832 specparam_declaration_instance4832();
    specparam_declaration4833 specparam_declaration_instance4833();
    specparam_declaration4834 specparam_declaration_instance4834();
    specparam_declaration4835 specparam_declaration_instance4835();
    specparam_declaration4836 specparam_declaration_instance4836();
    specparam_declaration4837 specparam_declaration_instance4837();
    specparam_declaration4838 specparam_declaration_instance4838();
    specparam_declaration4839 specparam_declaration_instance4839();
    specparam_declaration4840 specparam_declaration_instance4840();
    specparam_declaration4841 specparam_declaration_instance4841();
    specparam_declaration4842 specparam_declaration_instance4842();
    specparam_declaration4843 specparam_declaration_instance4843();
    specparam_declaration4844 specparam_declaration_instance4844();
    specparam_declaration4845 specparam_declaration_instance4845();
    specparam_declaration4846 specparam_declaration_instance4846();
    specparam_declaration4847 specparam_declaration_instance4847();
    specparam_declaration4848 specparam_declaration_instance4848();
    specparam_declaration4849 specparam_declaration_instance4849();
    specparam_declaration4850 specparam_declaration_instance4850();
    specparam_declaration4851 specparam_declaration_instance4851();
    specparam_declaration4852 specparam_declaration_instance4852();
    specparam_declaration4853 specparam_declaration_instance4853();
    specparam_declaration4854 specparam_declaration_instance4854();
    specparam_declaration4855 specparam_declaration_instance4855();
    specparam_declaration4856 specparam_declaration_instance4856();
    specparam_declaration4857 specparam_declaration_instance4857();
    specparam_declaration4858 specparam_declaration_instance4858();
    specparam_declaration4859 specparam_declaration_instance4859();
    specparam_declaration4860 specparam_declaration_instance4860();
    specparam_declaration4861 specparam_declaration_instance4861();
    specparam_declaration4862 specparam_declaration_instance4862();
    specparam_declaration4863 specparam_declaration_instance4863();
    specparam_declaration4864 specparam_declaration_instance4864();
    specparam_declaration4865 specparam_declaration_instance4865();
    specparam_declaration4866 specparam_declaration_instance4866();
    specparam_declaration4867 specparam_declaration_instance4867();
    specparam_declaration4868 specparam_declaration_instance4868();
    specparam_declaration4869 specparam_declaration_instance4869();
    specparam_declaration4870 specparam_declaration_instance4870();
    specparam_declaration4871 specparam_declaration_instance4871();
    specparam_declaration4872 specparam_declaration_instance4872();
    specparam_declaration4873 specparam_declaration_instance4873();
    specparam_declaration4874 specparam_declaration_instance4874();
    specparam_declaration4875 specparam_declaration_instance4875();
    specparam_declaration4876 specparam_declaration_instance4876();
    specparam_declaration4877 specparam_declaration_instance4877();
    specparam_declaration4878 specparam_declaration_instance4878();
    specparam_declaration4879 specparam_declaration_instance4879();
    specparam_declaration4880 specparam_declaration_instance4880();
    specparam_declaration4881 specparam_declaration_instance4881();
    specparam_declaration4882 specparam_declaration_instance4882();
    specparam_declaration4883 specparam_declaration_instance4883();
    specparam_declaration4884 specparam_declaration_instance4884();
    specparam_declaration4885 specparam_declaration_instance4885();
    specparam_declaration4886 specparam_declaration_instance4886();
    specparam_declaration4887 specparam_declaration_instance4887();
    specparam_declaration4888 specparam_declaration_instance4888();
    specparam_declaration4889 specparam_declaration_instance4889();
    specparam_declaration4890 specparam_declaration_instance4890();
    specparam_declaration4891 specparam_declaration_instance4891();
    specparam_declaration4892 specparam_declaration_instance4892();
    specparam_declaration4893 specparam_declaration_instance4893();
    specparam_declaration4894 specparam_declaration_instance4894();
    specparam_declaration4895 specparam_declaration_instance4895();
    specparam_declaration4896 specparam_declaration_instance4896();
    specparam_declaration4897 specparam_declaration_instance4897();
    specparam_declaration4898 specparam_declaration_instance4898();
    specparam_declaration4899 specparam_declaration_instance4899();
    specparam_declaration4900 specparam_declaration_instance4900();
    specparam_declaration4901 specparam_declaration_instance4901();
    specparam_declaration4902 specparam_declaration_instance4902();
    specparam_declaration4903 specparam_declaration_instance4903();
    specparam_declaration4904 specparam_declaration_instance4904();
    specparam_declaration4905 specparam_declaration_instance4905();
    specparam_declaration4906 specparam_declaration_instance4906();
    specparam_declaration4907 specparam_declaration_instance4907();
    specparam_declaration4908 specparam_declaration_instance4908();
    specparam_declaration4909 specparam_declaration_instance4909();
    specparam_declaration4910 specparam_declaration_instance4910();
    specparam_declaration4911 specparam_declaration_instance4911();
    specparam_declaration4912 specparam_declaration_instance4912();
    specparam_declaration4913 specparam_declaration_instance4913();
    specparam_declaration4914 specparam_declaration_instance4914();
    specparam_declaration4915 specparam_declaration_instance4915();
    specparam_declaration4916 specparam_declaration_instance4916();
    specparam_declaration4917 specparam_declaration_instance4917();
    specparam_declaration4918 specparam_declaration_instance4918();
    specparam_declaration4919 specparam_declaration_instance4919();
    specparam_declaration4920 specparam_declaration_instance4920();
    specparam_declaration4921 specparam_declaration_instance4921();
    specparam_declaration4922 specparam_declaration_instance4922();
    specparam_declaration4923 specparam_declaration_instance4923();
    specparam_declaration4924 specparam_declaration_instance4924();
    specparam_declaration4925 specparam_declaration_instance4925();
    specparam_declaration4926 specparam_declaration_instance4926();
    specparam_declaration4927 specparam_declaration_instance4927();
    specparam_declaration4928 specparam_declaration_instance4928();
    specparam_declaration4929 specparam_declaration_instance4929();
    specparam_declaration4930 specparam_declaration_instance4930();
    specparam_declaration4931 specparam_declaration_instance4931();
    specparam_declaration4932 specparam_declaration_instance4932();
    specparam_declaration4933 specparam_declaration_instance4933();
    specparam_declaration4934 specparam_declaration_instance4934();
    specparam_declaration4935 specparam_declaration_instance4935();
    specparam_declaration4936 specparam_declaration_instance4936();
    specparam_declaration4937 specparam_declaration_instance4937();
    specparam_declaration4938 specparam_declaration_instance4938();
    specparam_declaration4939 specparam_declaration_instance4939();
    specparam_declaration4940 specparam_declaration_instance4940();
    specparam_declaration4941 specparam_declaration_instance4941();
    specparam_declaration4942 specparam_declaration_instance4942();
    specparam_declaration4943 specparam_declaration_instance4943();
    specparam_declaration4944 specparam_declaration_instance4944();
    specparam_declaration4945 specparam_declaration_instance4945();
    specparam_declaration4946 specparam_declaration_instance4946();
    specparam_declaration4947 specparam_declaration_instance4947();
    specparam_declaration4948 specparam_declaration_instance4948();
    specparam_declaration4949 specparam_declaration_instance4949();
    specparam_declaration4950 specparam_declaration_instance4950();
    specparam_declaration4951 specparam_declaration_instance4951();
    specparam_declaration4952 specparam_declaration_instance4952();
    specparam_declaration4953 specparam_declaration_instance4953();
    specparam_declaration4954 specparam_declaration_instance4954();
    specparam_declaration4955 specparam_declaration_instance4955();
    specparam_declaration4956 specparam_declaration_instance4956();
    specparam_declaration4957 specparam_declaration_instance4957();
    specparam_declaration4958 specparam_declaration_instance4958();
    specparam_declaration4959 specparam_declaration_instance4959();
    specparam_declaration4960 specparam_declaration_instance4960();
    specparam_declaration4961 specparam_declaration_instance4961();
    specparam_declaration4962 specparam_declaration_instance4962();
    specparam_declaration4963 specparam_declaration_instance4963();
    specparam_declaration4964 specparam_declaration_instance4964();
    specparam_declaration4965 specparam_declaration_instance4965();
    specparam_declaration4966 specparam_declaration_instance4966();
    specparam_declaration4967 specparam_declaration_instance4967();
    specparam_declaration4968 specparam_declaration_instance4968();
    specparam_declaration4969 specparam_declaration_instance4969();
    specparam_declaration4970 specparam_declaration_instance4970();
    specparam_declaration4971 specparam_declaration_instance4971();
    specparam_declaration4972 specparam_declaration_instance4972();
    specparam_declaration4973 specparam_declaration_instance4973();
    specparam_declaration4974 specparam_declaration_instance4974();
    specparam_declaration4975 specparam_declaration_instance4975();
    specparam_declaration4976 specparam_declaration_instance4976();
    specparam_declaration4977 specparam_declaration_instance4977();
    specparam_declaration4978 specparam_declaration_instance4978();
    specparam_declaration4979 specparam_declaration_instance4979();
    specparam_declaration4980 specparam_declaration_instance4980();
    specparam_declaration4981 specparam_declaration_instance4981();
    specparam_declaration4982 specparam_declaration_instance4982();
    specparam_declaration4983 specparam_declaration_instance4983();
    specparam_declaration4984 specparam_declaration_instance4984();
    specparam_declaration4985 specparam_declaration_instance4985();
    specparam_declaration4986 specparam_declaration_instance4986();
    specparam_declaration4987 specparam_declaration_instance4987();
    specparam_declaration4988 specparam_declaration_instance4988();
    specparam_declaration4989 specparam_declaration_instance4989();
    specparam_declaration4990 specparam_declaration_instance4990();
    specparam_declaration4991 specparam_declaration_instance4991();
    specparam_declaration4992 specparam_declaration_instance4992();
    specparam_declaration4993 specparam_declaration_instance4993();
    specparam_declaration4994 specparam_declaration_instance4994();
    specparam_declaration4995 specparam_declaration_instance4995();
    specparam_declaration4996 specparam_declaration_instance4996();
    specparam_declaration4997 specparam_declaration_instance4997();
    specparam_declaration4998 specparam_declaration_instance4998();
    specparam_declaration4999 specparam_declaration_instance4999();
    specparam_declaration5000 specparam_declaration_instance5000();
    specparam_declaration5001 specparam_declaration_instance5001();
    specparam_declaration5002 specparam_declaration_instance5002();
    specparam_declaration5003 specparam_declaration_instance5003();
    specparam_declaration5004 specparam_declaration_instance5004();
    specparam_declaration5005 specparam_declaration_instance5005();
    specparam_declaration5006 specparam_declaration_instance5006();
    specparam_declaration5007 specparam_declaration_instance5007();
    specparam_declaration5008 specparam_declaration_instance5008();
    specparam_declaration5009 specparam_declaration_instance5009();
    specparam_declaration5010 specparam_declaration_instance5010();
    specparam_declaration5011 specparam_declaration_instance5011();
    specparam_declaration5012 specparam_declaration_instance5012();
    specparam_declaration5013 specparam_declaration_instance5013();
    specparam_declaration5014 specparam_declaration_instance5014();
    specparam_declaration5015 specparam_declaration_instance5015();
    specparam_declaration5016 specparam_declaration_instance5016();
    specparam_declaration5017 specparam_declaration_instance5017();
    specparam_declaration5018 specparam_declaration_instance5018();
    specparam_declaration5019 specparam_declaration_instance5019();
    specparam_declaration5020 specparam_declaration_instance5020();
    specparam_declaration5021 specparam_declaration_instance5021();
    specparam_declaration5022 specparam_declaration_instance5022();
    specparam_declaration5023 specparam_declaration_instance5023();
    specparam_declaration5024 specparam_declaration_instance5024();
    specparam_declaration5025 specparam_declaration_instance5025();
    specparam_declaration5026 specparam_declaration_instance5026();
    specparam_declaration5027 specparam_declaration_instance5027();
    specparam_declaration5028 specparam_declaration_instance5028();
    specparam_declaration5029 specparam_declaration_instance5029();
    specparam_declaration5030 specparam_declaration_instance5030();
    specparam_declaration5031 specparam_declaration_instance5031();
    specparam_declaration5032 specparam_declaration_instance5032();
    specparam_declaration5033 specparam_declaration_instance5033();
    specparam_declaration5034 specparam_declaration_instance5034();
    specparam_declaration5035 specparam_declaration_instance5035();
    specparam_declaration5036 specparam_declaration_instance5036();
    specparam_declaration5037 specparam_declaration_instance5037();
    specparam_declaration5038 specparam_declaration_instance5038();
    specparam_declaration5039 specparam_declaration_instance5039();
    specparam_declaration5040 specparam_declaration_instance5040();
    specparam_declaration5041 specparam_declaration_instance5041();
    specparam_declaration5042 specparam_declaration_instance5042();
    specparam_declaration5043 specparam_declaration_instance5043();
    specparam_declaration5044 specparam_declaration_instance5044();
    specparam_declaration5045 specparam_declaration_instance5045();
    specparam_declaration5046 specparam_declaration_instance5046();
    specparam_declaration5047 specparam_declaration_instance5047();
    specparam_declaration5048 specparam_declaration_instance5048();
    specparam_declaration5049 specparam_declaration_instance5049();
    specparam_declaration5050 specparam_declaration_instance5050();
    specparam_declaration5051 specparam_declaration_instance5051();
    specparam_declaration5052 specparam_declaration_instance5052();
    specparam_declaration5053 specparam_declaration_instance5053();
    specparam_declaration5054 specparam_declaration_instance5054();
    specparam_declaration5055 specparam_declaration_instance5055();
    specparam_declaration5056 specparam_declaration_instance5056();
    specparam_declaration5057 specparam_declaration_instance5057();
    specparam_declaration5058 specparam_declaration_instance5058();
    specparam_declaration5059 specparam_declaration_instance5059();
    specparam_declaration5060 specparam_declaration_instance5060();
    specparam_declaration5061 specparam_declaration_instance5061();
    specparam_declaration5062 specparam_declaration_instance5062();
    specparam_declaration5063 specparam_declaration_instance5063();
    specparam_declaration5064 specparam_declaration_instance5064();
    specparam_declaration5065 specparam_declaration_instance5065();
    specparam_declaration5066 specparam_declaration_instance5066();
    specparam_declaration5067 specparam_declaration_instance5067();
    specparam_declaration5068 specparam_declaration_instance5068();
    specparam_declaration5069 specparam_declaration_instance5069();
    specparam_declaration5070 specparam_declaration_instance5070();
    specparam_declaration5071 specparam_declaration_instance5071();
    specparam_declaration5072 specparam_declaration_instance5072();
    specparam_declaration5073 specparam_declaration_instance5073();
    specparam_declaration5074 specparam_declaration_instance5074();
    specparam_declaration5075 specparam_declaration_instance5075();
    specparam_declaration5076 specparam_declaration_instance5076();
    specparam_declaration5077 specparam_declaration_instance5077();
    specparam_declaration5078 specparam_declaration_instance5078();
    specparam_declaration5079 specparam_declaration_instance5079();
    specparam_declaration5080 specparam_declaration_instance5080();
    specparam_declaration5081 specparam_declaration_instance5081();
    specparam_declaration5082 specparam_declaration_instance5082();
    specparam_declaration5083 specparam_declaration_instance5083();
    specparam_declaration5084 specparam_declaration_instance5084();
    specparam_declaration5085 specparam_declaration_instance5085();
    specparam_declaration5086 specparam_declaration_instance5086();
    specparam_declaration5087 specparam_declaration_instance5087();
    specparam_declaration5088 specparam_declaration_instance5088();
    specparam_declaration5089 specparam_declaration_instance5089();
    specparam_declaration5090 specparam_declaration_instance5090();
    specparam_declaration5091 specparam_declaration_instance5091();
    specparam_declaration5092 specparam_declaration_instance5092();
    specparam_declaration5093 specparam_declaration_instance5093();
    specparam_declaration5094 specparam_declaration_instance5094();
    specparam_declaration5095 specparam_declaration_instance5095();
    specparam_declaration5096 specparam_declaration_instance5096();
    specparam_declaration5097 specparam_declaration_instance5097();
    specparam_declaration5098 specparam_declaration_instance5098();
    specparam_declaration5099 specparam_declaration_instance5099();
    specparam_declaration5100 specparam_declaration_instance5100();
    specparam_declaration5101 specparam_declaration_instance5101();
    specparam_declaration5102 specparam_declaration_instance5102();
    specparam_declaration5103 specparam_declaration_instance5103();
    specparam_declaration5104 specparam_declaration_instance5104();
    specparam_declaration5105 specparam_declaration_instance5105();
    specparam_declaration5106 specparam_declaration_instance5106();
    specparam_declaration5107 specparam_declaration_instance5107();
    specparam_declaration5108 specparam_declaration_instance5108();
    specparam_declaration5109 specparam_declaration_instance5109();
    specparam_declaration5110 specparam_declaration_instance5110();
    specparam_declaration5111 specparam_declaration_instance5111();
    specparam_declaration5112 specparam_declaration_instance5112();
    specparam_declaration5113 specparam_declaration_instance5113();
    specparam_declaration5114 specparam_declaration_instance5114();
    specparam_declaration5115 specparam_declaration_instance5115();
    specparam_declaration5116 specparam_declaration_instance5116();
    specparam_declaration5117 specparam_declaration_instance5117();
    specparam_declaration5118 specparam_declaration_instance5118();
    specparam_declaration5119 specparam_declaration_instance5119();
    specparam_declaration5120 specparam_declaration_instance5120();
    specparam_declaration5121 specparam_declaration_instance5121();
    specparam_declaration5122 specparam_declaration_instance5122();
    specparam_declaration5123 specparam_declaration_instance5123();
    specparam_declaration5124 specparam_declaration_instance5124();
    specparam_declaration5125 specparam_declaration_instance5125();
    specparam_declaration5126 specparam_declaration_instance5126();
    specparam_declaration5127 specparam_declaration_instance5127();
    specparam_declaration5128 specparam_declaration_instance5128();
    specparam_declaration5129 specparam_declaration_instance5129();
    specparam_declaration5130 specparam_declaration_instance5130();
    specparam_declaration5131 specparam_declaration_instance5131();
    specparam_declaration5132 specparam_declaration_instance5132();
    specparam_declaration5133 specparam_declaration_instance5133();
    specparam_declaration5134 specparam_declaration_instance5134();
    specparam_declaration5135 specparam_declaration_instance5135();
    specparam_declaration5136 specparam_declaration_instance5136();
    specparam_declaration5137 specparam_declaration_instance5137();
    specparam_declaration5138 specparam_declaration_instance5138();
    specparam_declaration5139 specparam_declaration_instance5139();
    specparam_declaration5140 specparam_declaration_instance5140();
    specparam_declaration5141 specparam_declaration_instance5141();
    specparam_declaration5142 specparam_declaration_instance5142();
    specparam_declaration5143 specparam_declaration_instance5143();
    specparam_declaration5144 specparam_declaration_instance5144();
    specparam_declaration5145 specparam_declaration_instance5145();
    specparam_declaration5146 specparam_declaration_instance5146();
    specparam_declaration5147 specparam_declaration_instance5147();
    specparam_declaration5148 specparam_declaration_instance5148();
    specparam_declaration5149 specparam_declaration_instance5149();
    specparam_declaration5150 specparam_declaration_instance5150();
    specparam_declaration5151 specparam_declaration_instance5151();
    specparam_declaration5152 specparam_declaration_instance5152();
    specparam_declaration5153 specparam_declaration_instance5153();
    specparam_declaration5154 specparam_declaration_instance5154();
    specparam_declaration5155 specparam_declaration_instance5155();
    specparam_declaration5156 specparam_declaration_instance5156();
    specparam_declaration5157 specparam_declaration_instance5157();
    specparam_declaration5158 specparam_declaration_instance5158();
    specparam_declaration5159 specparam_declaration_instance5159();
    specparam_declaration5160 specparam_declaration_instance5160();
    specparam_declaration5161 specparam_declaration_instance5161();
    specparam_declaration5162 specparam_declaration_instance5162();
    specparam_declaration5163 specparam_declaration_instance5163();
    specparam_declaration5164 specparam_declaration_instance5164();
    specparam_declaration5165 specparam_declaration_instance5165();
    specparam_declaration5166 specparam_declaration_instance5166();
    specparam_declaration5167 specparam_declaration_instance5167();
    specparam_declaration5168 specparam_declaration_instance5168();
    specparam_declaration5169 specparam_declaration_instance5169();
    specparam_declaration5170 specparam_declaration_instance5170();
    specparam_declaration5171 specparam_declaration_instance5171();
    specparam_declaration5172 specparam_declaration_instance5172();
    specparam_declaration5173 specparam_declaration_instance5173();
    specparam_declaration5174 specparam_declaration_instance5174();
    specparam_declaration5175 specparam_declaration_instance5175();
    specparam_declaration5176 specparam_declaration_instance5176();
    specparam_declaration5177 specparam_declaration_instance5177();
    specparam_declaration5178 specparam_declaration_instance5178();
    specparam_declaration5179 specparam_declaration_instance5179();
    specparam_declaration5180 specparam_declaration_instance5180();
    specparam_declaration5181 specparam_declaration_instance5181();
    specparam_declaration5182 specparam_declaration_instance5182();
    specparam_declaration5183 specparam_declaration_instance5183();
    specparam_declaration5184 specparam_declaration_instance5184();
    specparam_declaration5185 specparam_declaration_instance5185();
    specparam_declaration5186 specparam_declaration_instance5186();
    specparam_declaration5187 specparam_declaration_instance5187();
    specparam_declaration5188 specparam_declaration_instance5188();
    specparam_declaration5189 specparam_declaration_instance5189();
    specparam_declaration5190 specparam_declaration_instance5190();
    specparam_declaration5191 specparam_declaration_instance5191();
    specparam_declaration5192 specparam_declaration_instance5192();
    specparam_declaration5193 specparam_declaration_instance5193();
    specparam_declaration5194 specparam_declaration_instance5194();
    specparam_declaration5195 specparam_declaration_instance5195();
    specparam_declaration5196 specparam_declaration_instance5196();
    specparam_declaration5197 specparam_declaration_instance5197();
    specparam_declaration5198 specparam_declaration_instance5198();
    specparam_declaration5199 specparam_declaration_instance5199();
    specparam_declaration5200 specparam_declaration_instance5200();
    specparam_declaration5201 specparam_declaration_instance5201();
    specparam_declaration5202 specparam_declaration_instance5202();
    specparam_declaration5203 specparam_declaration_instance5203();
    specparam_declaration5204 specparam_declaration_instance5204();
    specparam_declaration5205 specparam_declaration_instance5205();
    specparam_declaration5206 specparam_declaration_instance5206();
    specparam_declaration5207 specparam_declaration_instance5207();
    specparam_declaration5208 specparam_declaration_instance5208();
    specparam_declaration5209 specparam_declaration_instance5209();
    specparam_declaration5210 specparam_declaration_instance5210();
    specparam_declaration5211 specparam_declaration_instance5211();
    specparam_declaration5212 specparam_declaration_instance5212();
    specparam_declaration5213 specparam_declaration_instance5213();
    specparam_declaration5214 specparam_declaration_instance5214();
    specparam_declaration5215 specparam_declaration_instance5215();
    specparam_declaration5216 specparam_declaration_instance5216();
    specparam_declaration5217 specparam_declaration_instance5217();
    specparam_declaration5218 specparam_declaration_instance5218();
    specparam_declaration5219 specparam_declaration_instance5219();
    specparam_declaration5220 specparam_declaration_instance5220();
    specparam_declaration5221 specparam_declaration_instance5221();
    specparam_declaration5222 specparam_declaration_instance5222();
    specparam_declaration5223 specparam_declaration_instance5223();
    specparam_declaration5224 specparam_declaration_instance5224();
    specparam_declaration5225 specparam_declaration_instance5225();
    specparam_declaration5226 specparam_declaration_instance5226();
    specparam_declaration5227 specparam_declaration_instance5227();
    specparam_declaration5228 specparam_declaration_instance5228();
    specparam_declaration5229 specparam_declaration_instance5229();
    specparam_declaration5230 specparam_declaration_instance5230();
    specparam_declaration5231 specparam_declaration_instance5231();
    specparam_declaration5232 specparam_declaration_instance5232();
    specparam_declaration5233 specparam_declaration_instance5233();
    specparam_declaration5234 specparam_declaration_instance5234();
    specparam_declaration5235 specparam_declaration_instance5235();
    specparam_declaration5236 specparam_declaration_instance5236();
    specparam_declaration5237 specparam_declaration_instance5237();
    specparam_declaration5238 specparam_declaration_instance5238();
    specparam_declaration5239 specparam_declaration_instance5239();
    specparam_declaration5240 specparam_declaration_instance5240();
    specparam_declaration5241 specparam_declaration_instance5241();
    specparam_declaration5242 specparam_declaration_instance5242();
    specparam_declaration5243 specparam_declaration_instance5243();
    specparam_declaration5244 specparam_declaration_instance5244();
    specparam_declaration5245 specparam_declaration_instance5245();
    specparam_declaration5246 specparam_declaration_instance5246();
    specparam_declaration5247 specparam_declaration_instance5247();
    specparam_declaration5248 specparam_declaration_instance5248();
    specparam_declaration5249 specparam_declaration_instance5249();
    specparam_declaration5250 specparam_declaration_instance5250();
    specparam_declaration5251 specparam_declaration_instance5251();
    specparam_declaration5252 specparam_declaration_instance5252();
    specparam_declaration5253 specparam_declaration_instance5253();
    specparam_declaration5254 specparam_declaration_instance5254();
    specparam_declaration5255 specparam_declaration_instance5255();
    specparam_declaration5256 specparam_declaration_instance5256();
    specparam_declaration5257 specparam_declaration_instance5257();
    specparam_declaration5258 specparam_declaration_instance5258();
    specparam_declaration5259 specparam_declaration_instance5259();
    specparam_declaration5260 specparam_declaration_instance5260();
    specparam_declaration5261 specparam_declaration_instance5261();
    specparam_declaration5262 specparam_declaration_instance5262();
    specparam_declaration5263 specparam_declaration_instance5263();
    specparam_declaration5264 specparam_declaration_instance5264();
    specparam_declaration5265 specparam_declaration_instance5265();
    specparam_declaration5266 specparam_declaration_instance5266();
    specparam_declaration5267 specparam_declaration_instance5267();
    specparam_declaration5268 specparam_declaration_instance5268();
    specparam_declaration5269 specparam_declaration_instance5269();
    specparam_declaration5270 specparam_declaration_instance5270();
    specparam_declaration5271 specparam_declaration_instance5271();
    specparam_declaration5272 specparam_declaration_instance5272();
    specparam_declaration5273 specparam_declaration_instance5273();
    specparam_declaration5274 specparam_declaration_instance5274();
    specparam_declaration5275 specparam_declaration_instance5275();
    specparam_declaration5276 specparam_declaration_instance5276();
    specparam_declaration5277 specparam_declaration_instance5277();
    specparam_declaration5278 specparam_declaration_instance5278();
    specparam_declaration5279 specparam_declaration_instance5279();
    specparam_declaration5280 specparam_declaration_instance5280();
    specparam_declaration5281 specparam_declaration_instance5281();
    specparam_declaration5282 specparam_declaration_instance5282();
    specparam_declaration5283 specparam_declaration_instance5283();
    specparam_declaration5284 specparam_declaration_instance5284();
    specparam_declaration5285 specparam_declaration_instance5285();
    specparam_declaration5286 specparam_declaration_instance5286();
    specparam_declaration5287 specparam_declaration_instance5287();
    specparam_declaration5288 specparam_declaration_instance5288();
    specparam_declaration5289 specparam_declaration_instance5289();
    specparam_declaration5290 specparam_declaration_instance5290();
    specparam_declaration5291 specparam_declaration_instance5291();
    specparam_declaration5292 specparam_declaration_instance5292();
    specparam_declaration5293 specparam_declaration_instance5293();
    specparam_declaration5294 specparam_declaration_instance5294();
    specparam_declaration5295 specparam_declaration_instance5295();
    specparam_declaration5296 specparam_declaration_instance5296();
    specparam_declaration5297 specparam_declaration_instance5297();
    specparam_declaration5298 specparam_declaration_instance5298();
    specparam_declaration5299 specparam_declaration_instance5299();
    specparam_declaration5300 specparam_declaration_instance5300();
    specparam_declaration5301 specparam_declaration_instance5301();
    specparam_declaration5302 specparam_declaration_instance5302();
    specparam_declaration5303 specparam_declaration_instance5303();
    specparam_declaration5304 specparam_declaration_instance5304();
    specparam_declaration5305 specparam_declaration_instance5305();
    specparam_declaration5306 specparam_declaration_instance5306();
    specparam_declaration5307 specparam_declaration_instance5307();
    specparam_declaration5308 specparam_declaration_instance5308();
    specparam_declaration5309 specparam_declaration_instance5309();
    specparam_declaration5310 specparam_declaration_instance5310();
    specparam_declaration5311 specparam_declaration_instance5311();
    specparam_declaration5312 specparam_declaration_instance5312();
    specparam_declaration5313 specparam_declaration_instance5313();
    specparam_declaration5314 specparam_declaration_instance5314();
    specparam_declaration5315 specparam_declaration_instance5315();
    specparam_declaration5316 specparam_declaration_instance5316();
    specparam_declaration5317 specparam_declaration_instance5317();
    specparam_declaration5318 specparam_declaration_instance5318();
    specparam_declaration5319 specparam_declaration_instance5319();
    specparam_declaration5320 specparam_declaration_instance5320();
    specparam_declaration5321 specparam_declaration_instance5321();
    specparam_declaration5322 specparam_declaration_instance5322();
    specparam_declaration5323 specparam_declaration_instance5323();
    specparam_declaration5324 specparam_declaration_instance5324();
    specparam_declaration5325 specparam_declaration_instance5325();
    specparam_declaration5326 specparam_declaration_instance5326();
    specparam_declaration5327 specparam_declaration_instance5327();
    specparam_declaration5328 specparam_declaration_instance5328();
    specparam_declaration5329 specparam_declaration_instance5329();
    specparam_declaration5330 specparam_declaration_instance5330();
    specparam_declaration5331 specparam_declaration_instance5331();
    specparam_declaration5332 specparam_declaration_instance5332();
    specparam_declaration5333 specparam_declaration_instance5333();
    specparam_declaration5334 specparam_declaration_instance5334();
    specparam_declaration5335 specparam_declaration_instance5335();
    specparam_declaration5336 specparam_declaration_instance5336();
    specparam_declaration5337 specparam_declaration_instance5337();
    specparam_declaration5338 specparam_declaration_instance5338();
    specparam_declaration5339 specparam_declaration_instance5339();
    specparam_declaration5340 specparam_declaration_instance5340();
    specparam_declaration5341 specparam_declaration_instance5341();
    specparam_declaration5342 specparam_declaration_instance5342();
    specparam_declaration5343 specparam_declaration_instance5343();
    specparam_declaration5344 specparam_declaration_instance5344();
    specparam_declaration5345 specparam_declaration_instance5345();
    specparam_declaration5346 specparam_declaration_instance5346();
    specparam_declaration5347 specparam_declaration_instance5347();
    specparam_declaration5348 specparam_declaration_instance5348();
    specparam_declaration5349 specparam_declaration_instance5349();
    specparam_declaration5350 specparam_declaration_instance5350();
    specparam_declaration5351 specparam_declaration_instance5351();
    specparam_declaration5352 specparam_declaration_instance5352();
    specparam_declaration5353 specparam_declaration_instance5353();
    specparam_declaration5354 specparam_declaration_instance5354();
    specparam_declaration5355 specparam_declaration_instance5355();
    specparam_declaration5356 specparam_declaration_instance5356();
    specparam_declaration5357 specparam_declaration_instance5357();
    specparam_declaration5358 specparam_declaration_instance5358();
    specparam_declaration5359 specparam_declaration_instance5359();
    specparam_declaration5360 specparam_declaration_instance5360();
    specparam_declaration5361 specparam_declaration_instance5361();
    specparam_declaration5362 specparam_declaration_instance5362();
    specparam_declaration5363 specparam_declaration_instance5363();
    specparam_declaration5364 specparam_declaration_instance5364();
    specparam_declaration5365 specparam_declaration_instance5365();
    specparam_declaration5366 specparam_declaration_instance5366();
    specparam_declaration5367 specparam_declaration_instance5367();
    specparam_declaration5368 specparam_declaration_instance5368();
    specparam_declaration5369 specparam_declaration_instance5369();
    specparam_declaration5370 specparam_declaration_instance5370();
    specparam_declaration5371 specparam_declaration_instance5371();
    specparam_declaration5372 specparam_declaration_instance5372();
    specparam_declaration5373 specparam_declaration_instance5373();
    specparam_declaration5374 specparam_declaration_instance5374();
    specparam_declaration5375 specparam_declaration_instance5375();
    specparam_declaration5376 specparam_declaration_instance5376();
    specparam_declaration5377 specparam_declaration_instance5377();
    specparam_declaration5378 specparam_declaration_instance5378();
    specparam_declaration5379 specparam_declaration_instance5379();
    specparam_declaration5380 specparam_declaration_instance5380();
    specparam_declaration5381 specparam_declaration_instance5381();
    specparam_declaration5382 specparam_declaration_instance5382();
    specparam_declaration5383 specparam_declaration_instance5383();
    specparam_declaration5384 specparam_declaration_instance5384();
    specparam_declaration5385 specparam_declaration_instance5385();
    specparam_declaration5386 specparam_declaration_instance5386();
    specparam_declaration5387 specparam_declaration_instance5387();
    specparam_declaration5388 specparam_declaration_instance5388();
    specparam_declaration5389 specparam_declaration_instance5389();
    specparam_declaration5390 specparam_declaration_instance5390();
    specparam_declaration5391 specparam_declaration_instance5391();
    specparam_declaration5392 specparam_declaration_instance5392();
    specparam_declaration5393 specparam_declaration_instance5393();
    specparam_declaration5394 specparam_declaration_instance5394();
    specparam_declaration5395 specparam_declaration_instance5395();
    specparam_declaration5396 specparam_declaration_instance5396();
    specparam_declaration5397 specparam_declaration_instance5397();
    specparam_declaration5398 specparam_declaration_instance5398();
    specparam_declaration5399 specparam_declaration_instance5399();
    specparam_declaration5400 specparam_declaration_instance5400();
    specparam_declaration5401 specparam_declaration_instance5401();
    specparam_declaration5402 specparam_declaration_instance5402();
    specparam_declaration5403 specparam_declaration_instance5403();
    specparam_declaration5404 specparam_declaration_instance5404();
    specparam_declaration5405 specparam_declaration_instance5405();
    specparam_declaration5406 specparam_declaration_instance5406();
    specparam_declaration5407 specparam_declaration_instance5407();
    specparam_declaration5408 specparam_declaration_instance5408();
    specparam_declaration5409 specparam_declaration_instance5409();
    specparam_declaration5410 specparam_declaration_instance5410();
    specparam_declaration5411 specparam_declaration_instance5411();
    specparam_declaration5412 specparam_declaration_instance5412();
    specparam_declaration5413 specparam_declaration_instance5413();
    specparam_declaration5414 specparam_declaration_instance5414();
    specparam_declaration5415 specparam_declaration_instance5415();
    specparam_declaration5416 specparam_declaration_instance5416();
    specparam_declaration5417 specparam_declaration_instance5417();
    specparam_declaration5418 specparam_declaration_instance5418();
    specparam_declaration5419 specparam_declaration_instance5419();
    specparam_declaration5420 specparam_declaration_instance5420();
    specparam_declaration5421 specparam_declaration_instance5421();
    specparam_declaration5422 specparam_declaration_instance5422();
    specparam_declaration5423 specparam_declaration_instance5423();
    specparam_declaration5424 specparam_declaration_instance5424();
    specparam_declaration5425 specparam_declaration_instance5425();
    specparam_declaration5426 specparam_declaration_instance5426();
    specparam_declaration5427 specparam_declaration_instance5427();
    specparam_declaration5428 specparam_declaration_instance5428();
    specparam_declaration5429 specparam_declaration_instance5429();
    specparam_declaration5430 specparam_declaration_instance5430();
    specparam_declaration5431 specparam_declaration_instance5431();
    specparam_declaration5432 specparam_declaration_instance5432();
    specparam_declaration5433 specparam_declaration_instance5433();
    specparam_declaration5434 specparam_declaration_instance5434();
    specparam_declaration5435 specparam_declaration_instance5435();
    specparam_declaration5436 specparam_declaration_instance5436();
    specparam_declaration5437 specparam_declaration_instance5437();
    specparam_declaration5438 specparam_declaration_instance5438();
    specparam_declaration5439 specparam_declaration_instance5439();
    specparam_declaration5440 specparam_declaration_instance5440();
    specparam_declaration5441 specparam_declaration_instance5441();
    specparam_declaration5442 specparam_declaration_instance5442();
    specparam_declaration5443 specparam_declaration_instance5443();
    specparam_declaration5444 specparam_declaration_instance5444();
    specparam_declaration5445 specparam_declaration_instance5445();
    specparam_declaration5446 specparam_declaration_instance5446();
    specparam_declaration5447 specparam_declaration_instance5447();
    specparam_declaration5448 specparam_declaration_instance5448();
    specparam_declaration5449 specparam_declaration_instance5449();
    specparam_declaration5450 specparam_declaration_instance5450();
    specparam_declaration5451 specparam_declaration_instance5451();
    specparam_declaration5452 specparam_declaration_instance5452();
    specparam_declaration5453 specparam_declaration_instance5453();
    specparam_declaration5454 specparam_declaration_instance5454();
    specparam_declaration5455 specparam_declaration_instance5455();
    specparam_declaration5456 specparam_declaration_instance5456();
    specparam_declaration5457 specparam_declaration_instance5457();
    specparam_declaration5458 specparam_declaration_instance5458();
    specparam_declaration5459 specparam_declaration_instance5459();
    specparam_declaration5460 specparam_declaration_instance5460();
    specparam_declaration5461 specparam_declaration_instance5461();
    specparam_declaration5462 specparam_declaration_instance5462();
    specparam_declaration5463 specparam_declaration_instance5463();
    specparam_declaration5464 specparam_declaration_instance5464();
    specparam_declaration5465 specparam_declaration_instance5465();
    specparam_declaration5466 specparam_declaration_instance5466();
    specparam_declaration5467 specparam_declaration_instance5467();
    specparam_declaration5468 specparam_declaration_instance5468();
    specparam_declaration5469 specparam_declaration_instance5469();
    specparam_declaration5470 specparam_declaration_instance5470();
    specparam_declaration5471 specparam_declaration_instance5471();
    specparam_declaration5472 specparam_declaration_instance5472();
    specparam_declaration5473 specparam_declaration_instance5473();
    specparam_declaration5474 specparam_declaration_instance5474();
    specparam_declaration5475 specparam_declaration_instance5475();
    specparam_declaration5476 specparam_declaration_instance5476();
    specparam_declaration5477 specparam_declaration_instance5477();
    specparam_declaration5478 specparam_declaration_instance5478();
    specparam_declaration5479 specparam_declaration_instance5479();
    specparam_declaration5480 specparam_declaration_instance5480();
    specparam_declaration5481 specparam_declaration_instance5481();
    specparam_declaration5482 specparam_declaration_instance5482();
    specparam_declaration5483 specparam_declaration_instance5483();
    specparam_declaration5484 specparam_declaration_instance5484();
    specparam_declaration5485 specparam_declaration_instance5485();
    specparam_declaration5486 specparam_declaration_instance5486();
    specparam_declaration5487 specparam_declaration_instance5487();
    specparam_declaration5488 specparam_declaration_instance5488();
    specparam_declaration5489 specparam_declaration_instance5489();
    specparam_declaration5490 specparam_declaration_instance5490();
    specparam_declaration5491 specparam_declaration_instance5491();
    specparam_declaration5492 specparam_declaration_instance5492();
    specparam_declaration5493 specparam_declaration_instance5493();
    specparam_declaration5494 specparam_declaration_instance5494();
    specparam_declaration5495 specparam_declaration_instance5495();
    specparam_declaration5496 specparam_declaration_instance5496();
    specparam_declaration5497 specparam_declaration_instance5497();
    specparam_declaration5498 specparam_declaration_instance5498();
    specparam_declaration5499 specparam_declaration_instance5499();
    specparam_declaration5500 specparam_declaration_instance5500();
    specparam_declaration5501 specparam_declaration_instance5501();
    specparam_declaration5502 specparam_declaration_instance5502();
    specparam_declaration5503 specparam_declaration_instance5503();
    specparam_declaration5504 specparam_declaration_instance5504();
    specparam_declaration5505 specparam_declaration_instance5505();
    specparam_declaration5506 specparam_declaration_instance5506();
    specparam_declaration5507 specparam_declaration_instance5507();
    specparam_declaration5508 specparam_declaration_instance5508();
    specparam_declaration5509 specparam_declaration_instance5509();
    specparam_declaration5510 specparam_declaration_instance5510();
    specparam_declaration5511 specparam_declaration_instance5511();
    specparam_declaration5512 specparam_declaration_instance5512();
    specparam_declaration5513 specparam_declaration_instance5513();
    specparam_declaration5514 specparam_declaration_instance5514();
    specparam_declaration5515 specparam_declaration_instance5515();
    specparam_declaration5516 specparam_declaration_instance5516();
    specparam_declaration5517 specparam_declaration_instance5517();
    specparam_declaration5518 specparam_declaration_instance5518();
    specparam_declaration5519 specparam_declaration_instance5519();
    specparam_declaration5520 specparam_declaration_instance5520();
    specparam_declaration5521 specparam_declaration_instance5521();
    specparam_declaration5522 specparam_declaration_instance5522();
    specparam_declaration5523 specparam_declaration_instance5523();
    specparam_declaration5524 specparam_declaration_instance5524();
    specparam_declaration5525 specparam_declaration_instance5525();
    specparam_declaration5526 specparam_declaration_instance5526();
    specparam_declaration5527 specparam_declaration_instance5527();
    specparam_declaration5528 specparam_declaration_instance5528();
    specparam_declaration5529 specparam_declaration_instance5529();
    specparam_declaration5530 specparam_declaration_instance5530();
    specparam_declaration5531 specparam_declaration_instance5531();
    specparam_declaration5532 specparam_declaration_instance5532();
    specparam_declaration5533 specparam_declaration_instance5533();
    specparam_declaration5534 specparam_declaration_instance5534();
    specparam_declaration5535 specparam_declaration_instance5535();
    specparam_declaration5536 specparam_declaration_instance5536();
    specparam_declaration5537 specparam_declaration_instance5537();
    specparam_declaration5538 specparam_declaration_instance5538();
    specparam_declaration5539 specparam_declaration_instance5539();
    specparam_declaration5540 specparam_declaration_instance5540();
    specparam_declaration5541 specparam_declaration_instance5541();
    specparam_declaration5542 specparam_declaration_instance5542();
    specparam_declaration5543 specparam_declaration_instance5543();
    specparam_declaration5544 specparam_declaration_instance5544();
    specparam_declaration5545 specparam_declaration_instance5545();
    specparam_declaration5546 specparam_declaration_instance5546();
    specparam_declaration5547 specparam_declaration_instance5547();
    specparam_declaration5548 specparam_declaration_instance5548();
    specparam_declaration5549 specparam_declaration_instance5549();
    specparam_declaration5550 specparam_declaration_instance5550();
    specparam_declaration5551 specparam_declaration_instance5551();
    specparam_declaration5552 specparam_declaration_instance5552();
    specparam_declaration5553 specparam_declaration_instance5553();
    specparam_declaration5554 specparam_declaration_instance5554();
    specparam_declaration5555 specparam_declaration_instance5555();
    specparam_declaration5556 specparam_declaration_instance5556();
    specparam_declaration5557 specparam_declaration_instance5557();
    specparam_declaration5558 specparam_declaration_instance5558();
    specparam_declaration5559 specparam_declaration_instance5559();
    specparam_declaration5560 specparam_declaration_instance5560();
    specparam_declaration5561 specparam_declaration_instance5561();
    specparam_declaration5562 specparam_declaration_instance5562();
    specparam_declaration5563 specparam_declaration_instance5563();
    specparam_declaration5564 specparam_declaration_instance5564();
    specparam_declaration5565 specparam_declaration_instance5565();
    specparam_declaration5566 specparam_declaration_instance5566();
    specparam_declaration5567 specparam_declaration_instance5567();
    specparam_declaration5568 specparam_declaration_instance5568();
    specparam_declaration5569 specparam_declaration_instance5569();
    specparam_declaration5570 specparam_declaration_instance5570();
    specparam_declaration5571 specparam_declaration_instance5571();
    specparam_declaration5572 specparam_declaration_instance5572();
    specparam_declaration5573 specparam_declaration_instance5573();
    specparam_declaration5574 specparam_declaration_instance5574();
    specparam_declaration5575 specparam_declaration_instance5575();
    specparam_declaration5576 specparam_declaration_instance5576();
    specparam_declaration5577 specparam_declaration_instance5577();
    specparam_declaration5578 specparam_declaration_instance5578();
    specparam_declaration5579 specparam_declaration_instance5579();
    specparam_declaration5580 specparam_declaration_instance5580();
    specparam_declaration5581 specparam_declaration_instance5581();
    specparam_declaration5582 specparam_declaration_instance5582();
    specparam_declaration5583 specparam_declaration_instance5583();
    specparam_declaration5584 specparam_declaration_instance5584();
    specparam_declaration5585 specparam_declaration_instance5585();
    specparam_declaration5586 specparam_declaration_instance5586();
    specparam_declaration5587 specparam_declaration_instance5587();
    specparam_declaration5588 specparam_declaration_instance5588();
    specparam_declaration5589 specparam_declaration_instance5589();
    specparam_declaration5590 specparam_declaration_instance5590();
    specparam_declaration5591 specparam_declaration_instance5591();
    specparam_declaration5592 specparam_declaration_instance5592();
    specparam_declaration5593 specparam_declaration_instance5593();
    specparam_declaration5594 specparam_declaration_instance5594();
    specparam_declaration5595 specparam_declaration_instance5595();
    specparam_declaration5596 specparam_declaration_instance5596();
    specparam_declaration5597 specparam_declaration_instance5597();
    specparam_declaration5598 specparam_declaration_instance5598();
    specparam_declaration5599 specparam_declaration_instance5599();
    specparam_declaration5600 specparam_declaration_instance5600();
    specparam_declaration5601 specparam_declaration_instance5601();
    specparam_declaration5602 specparam_declaration_instance5602();
    specparam_declaration5603 specparam_declaration_instance5603();
    specparam_declaration5604 specparam_declaration_instance5604();
    specparam_declaration5605 specparam_declaration_instance5605();
    specparam_declaration5606 specparam_declaration_instance5606();
    specparam_declaration5607 specparam_declaration_instance5607();
    specparam_declaration5608 specparam_declaration_instance5608();
    specparam_declaration5609 specparam_declaration_instance5609();
    specparam_declaration5610 specparam_declaration_instance5610();
    specparam_declaration5611 specparam_declaration_instance5611();
    specparam_declaration5612 specparam_declaration_instance5612();
    specparam_declaration5613 specparam_declaration_instance5613();
    specparam_declaration5614 specparam_declaration_instance5614();
    specparam_declaration5615 specparam_declaration_instance5615();
    specparam_declaration5616 specparam_declaration_instance5616();
    specparam_declaration5617 specparam_declaration_instance5617();
    specparam_declaration5618 specparam_declaration_instance5618();
    specparam_declaration5619 specparam_declaration_instance5619();
    specparam_declaration5620 specparam_declaration_instance5620();
    specparam_declaration5621 specparam_declaration_instance5621();
    specparam_declaration5622 specparam_declaration_instance5622();
    specparam_declaration5623 specparam_declaration_instance5623();
    specparam_declaration5624 specparam_declaration_instance5624();
    specparam_declaration5625 specparam_declaration_instance5625();
    specparam_declaration5626 specparam_declaration_instance5626();
    specparam_declaration5627 specparam_declaration_instance5627();
    specparam_declaration5628 specparam_declaration_instance5628();
    specparam_declaration5629 specparam_declaration_instance5629();
    specparam_declaration5630 specparam_declaration_instance5630();
    specparam_declaration5631 specparam_declaration_instance5631();
    specparam_declaration5632 specparam_declaration_instance5632();
    specparam_declaration5633 specparam_declaration_instance5633();
    specparam_declaration5634 specparam_declaration_instance5634();
    specparam_declaration5635 specparam_declaration_instance5635();
    specparam_declaration5636 specparam_declaration_instance5636();
    specparam_declaration5637 specparam_declaration_instance5637();
    specparam_declaration5638 specparam_declaration_instance5638();
    specparam_declaration5639 specparam_declaration_instance5639();
    specparam_declaration5640 specparam_declaration_instance5640();
    specparam_declaration5641 specparam_declaration_instance5641();
    specparam_declaration5642 specparam_declaration_instance5642();
    specparam_declaration5643 specparam_declaration_instance5643();
    specparam_declaration5644 specparam_declaration_instance5644();
    specparam_declaration5645 specparam_declaration_instance5645();
    specparam_declaration5646 specparam_declaration_instance5646();
    specparam_declaration5647 specparam_declaration_instance5647();
    specparam_declaration5648 specparam_declaration_instance5648();
    specparam_declaration5649 specparam_declaration_instance5649();
    specparam_declaration5650 specparam_declaration_instance5650();
    specparam_declaration5651 specparam_declaration_instance5651();
    specparam_declaration5652 specparam_declaration_instance5652();
    specparam_declaration5653 specparam_declaration_instance5653();
    specparam_declaration5654 specparam_declaration_instance5654();
    specparam_declaration5655 specparam_declaration_instance5655();
    specparam_declaration5656 specparam_declaration_instance5656();
    specparam_declaration5657 specparam_declaration_instance5657();
    specparam_declaration5658 specparam_declaration_instance5658();
    specparam_declaration5659 specparam_declaration_instance5659();
    specparam_declaration5660 specparam_declaration_instance5660();
    specparam_declaration5661 specparam_declaration_instance5661();
    specparam_declaration5662 specparam_declaration_instance5662();
    specparam_declaration5663 specparam_declaration_instance5663();
    specparam_declaration5664 specparam_declaration_instance5664();
    specparam_declaration5665 specparam_declaration_instance5665();
    specparam_declaration5666 specparam_declaration_instance5666();
    specparam_declaration5667 specparam_declaration_instance5667();
    specparam_declaration5668 specparam_declaration_instance5668();
    specparam_declaration5669 specparam_declaration_instance5669();
    specparam_declaration5670 specparam_declaration_instance5670();
    specparam_declaration5671 specparam_declaration_instance5671();
    specparam_declaration5672 specparam_declaration_instance5672();
    specparam_declaration5673 specparam_declaration_instance5673();
    specparam_declaration5674 specparam_declaration_instance5674();
    specparam_declaration5675 specparam_declaration_instance5675();
    specparam_declaration5676 specparam_declaration_instance5676();
    specparam_declaration5677 specparam_declaration_instance5677();
    specparam_declaration5678 specparam_declaration_instance5678();
    specparam_declaration5679 specparam_declaration_instance5679();
    specparam_declaration5680 specparam_declaration_instance5680();
    specparam_declaration5681 specparam_declaration_instance5681();
    specparam_declaration5682 specparam_declaration_instance5682();
    specparam_declaration5683 specparam_declaration_instance5683();
    specparam_declaration5684 specparam_declaration_instance5684();
    specparam_declaration5685 specparam_declaration_instance5685();
    specparam_declaration5686 specparam_declaration_instance5686();
    specparam_declaration5687 specparam_declaration_instance5687();
    specparam_declaration5688 specparam_declaration_instance5688();
    specparam_declaration5689 specparam_declaration_instance5689();
    specparam_declaration5690 specparam_declaration_instance5690();
    specparam_declaration5691 specparam_declaration_instance5691();
    specparam_declaration5692 specparam_declaration_instance5692();
    specparam_declaration5693 specparam_declaration_instance5693();
    specparam_declaration5694 specparam_declaration_instance5694();
    specparam_declaration5695 specparam_declaration_instance5695();
    specparam_declaration5696 specparam_declaration_instance5696();
    specparam_declaration5697 specparam_declaration_instance5697();
    specparam_declaration5698 specparam_declaration_instance5698();
    specparam_declaration5699 specparam_declaration_instance5699();
    specparam_declaration5700 specparam_declaration_instance5700();
    specparam_declaration5701 specparam_declaration_instance5701();
    specparam_declaration5702 specparam_declaration_instance5702();
    specparam_declaration5703 specparam_declaration_instance5703();
    specparam_declaration5704 specparam_declaration_instance5704();
    specparam_declaration5705 specparam_declaration_instance5705();
    specparam_declaration5706 specparam_declaration_instance5706();
    specparam_declaration5707 specparam_declaration_instance5707();
    specparam_declaration5708 specparam_declaration_instance5708();
    specparam_declaration5709 specparam_declaration_instance5709();
    specparam_declaration5710 specparam_declaration_instance5710();
    specparam_declaration5711 specparam_declaration_instance5711();
    specparam_declaration5712 specparam_declaration_instance5712();
    specparam_declaration5713 specparam_declaration_instance5713();
    specparam_declaration5714 specparam_declaration_instance5714();
    specparam_declaration5715 specparam_declaration_instance5715();
    specparam_declaration5716 specparam_declaration_instance5716();
    specparam_declaration5717 specparam_declaration_instance5717();
    specparam_declaration5718 specparam_declaration_instance5718();
    specparam_declaration5719 specparam_declaration_instance5719();
    specparam_declaration5720 specparam_declaration_instance5720();
    specparam_declaration5721 specparam_declaration_instance5721();
    specparam_declaration5722 specparam_declaration_instance5722();
    specparam_declaration5723 specparam_declaration_instance5723();
    specparam_declaration5724 specparam_declaration_instance5724();
    specparam_declaration5725 specparam_declaration_instance5725();
    specparam_declaration5726 specparam_declaration_instance5726();
    specparam_declaration5727 specparam_declaration_instance5727();
    specparam_declaration5728 specparam_declaration_instance5728();
    specparam_declaration5729 specparam_declaration_instance5729();
    specparam_declaration5730 specparam_declaration_instance5730();
    specparam_declaration5731 specparam_declaration_instance5731();
    specparam_declaration5732 specparam_declaration_instance5732();
    specparam_declaration5733 specparam_declaration_instance5733();
    specparam_declaration5734 specparam_declaration_instance5734();
    specparam_declaration5735 specparam_declaration_instance5735();
    specparam_declaration5736 specparam_declaration_instance5736();
    specparam_declaration5737 specparam_declaration_instance5737();
    specparam_declaration5738 specparam_declaration_instance5738();
    specparam_declaration5739 specparam_declaration_instance5739();
    specparam_declaration5740 specparam_declaration_instance5740();
    specparam_declaration5741 specparam_declaration_instance5741();
    specparam_declaration5742 specparam_declaration_instance5742();
    specparam_declaration5743 specparam_declaration_instance5743();
    specparam_declaration5744 specparam_declaration_instance5744();
    specparam_declaration5745 specparam_declaration_instance5745();
    specparam_declaration5746 specparam_declaration_instance5746();
    specparam_declaration5747 specparam_declaration_instance5747();
    specparam_declaration5748 specparam_declaration_instance5748();
    specparam_declaration5749 specparam_declaration_instance5749();
    specparam_declaration5750 specparam_declaration_instance5750();
    specparam_declaration5751 specparam_declaration_instance5751();
    specparam_declaration5752 specparam_declaration_instance5752();
    specparam_declaration5753 specparam_declaration_instance5753();
    specparam_declaration5754 specparam_declaration_instance5754();
    specparam_declaration5755 specparam_declaration_instance5755();
    specparam_declaration5756 specparam_declaration_instance5756();
    specparam_declaration5757 specparam_declaration_instance5757();
    specparam_declaration5758 specparam_declaration_instance5758();
    specparam_declaration5759 specparam_declaration_instance5759();
    specparam_declaration5760 specparam_declaration_instance5760();
    specparam_declaration5761 specparam_declaration_instance5761();
    specparam_declaration5762 specparam_declaration_instance5762();
    specparam_declaration5763 specparam_declaration_instance5763();
    specparam_declaration5764 specparam_declaration_instance5764();
    specparam_declaration5765 specparam_declaration_instance5765();
    specparam_declaration5766 specparam_declaration_instance5766();
    specparam_declaration5767 specparam_declaration_instance5767();
    specparam_declaration5768 specparam_declaration_instance5768();
    specparam_declaration5769 specparam_declaration_instance5769();
    specparam_declaration5770 specparam_declaration_instance5770();
    specparam_declaration5771 specparam_declaration_instance5771();
    specparam_declaration5772 specparam_declaration_instance5772();
    specparam_declaration5773 specparam_declaration_instance5773();
    specparam_declaration5774 specparam_declaration_instance5774();
    specparam_declaration5775 specparam_declaration_instance5775();
    specparam_declaration5776 specparam_declaration_instance5776();
    specparam_declaration5777 specparam_declaration_instance5777();
    specparam_declaration5778 specparam_declaration_instance5778();
    specparam_declaration5779 specparam_declaration_instance5779();
    specparam_declaration5780 specparam_declaration_instance5780();
    specparam_declaration5781 specparam_declaration_instance5781();
    specparam_declaration5782 specparam_declaration_instance5782();
    specparam_declaration5783 specparam_declaration_instance5783();
    specparam_declaration5784 specparam_declaration_instance5784();
    specparam_declaration5785 specparam_declaration_instance5785();
    specparam_declaration5786 specparam_declaration_instance5786();
    specparam_declaration5787 specparam_declaration_instance5787();
    specparam_declaration5788 specparam_declaration_instance5788();
    specparam_declaration5789 specparam_declaration_instance5789();
    specparam_declaration5790 specparam_declaration_instance5790();
    specparam_declaration5791 specparam_declaration_instance5791();
    specparam_declaration5792 specparam_declaration_instance5792();
    specparam_declaration5793 specparam_declaration_instance5793();
    specparam_declaration5794 specparam_declaration_instance5794();
    specparam_declaration5795 specparam_declaration_instance5795();
    specparam_declaration5796 specparam_declaration_instance5796();
    specparam_declaration5797 specparam_declaration_instance5797();
    specparam_declaration5798 specparam_declaration_instance5798();
    specparam_declaration5799 specparam_declaration_instance5799();
    specparam_declaration5800 specparam_declaration_instance5800();
    specparam_declaration5801 specparam_declaration_instance5801();
    specparam_declaration5802 specparam_declaration_instance5802();
    specparam_declaration5803 specparam_declaration_instance5803();
    specparam_declaration5804 specparam_declaration_instance5804();
    specparam_declaration5805 specparam_declaration_instance5805();
    specparam_declaration5806 specparam_declaration_instance5806();
    specparam_declaration5807 specparam_declaration_instance5807();
    specparam_declaration5808 specparam_declaration_instance5808();
    specparam_declaration5809 specparam_declaration_instance5809();
    specparam_declaration5810 specparam_declaration_instance5810();
    specparam_declaration5811 specparam_declaration_instance5811();
    specparam_declaration5812 specparam_declaration_instance5812();
    specparam_declaration5813 specparam_declaration_instance5813();
    specparam_declaration5814 specparam_declaration_instance5814();
    specparam_declaration5815 specparam_declaration_instance5815();
    specparam_declaration5816 specparam_declaration_instance5816();
    specparam_declaration5817 specparam_declaration_instance5817();
    specparam_declaration5818 specparam_declaration_instance5818();
    specparam_declaration5819 specparam_declaration_instance5819();
    specparam_declaration5820 specparam_declaration_instance5820();
    specparam_declaration5821 specparam_declaration_instance5821();
    specparam_declaration5822 specparam_declaration_instance5822();
    specparam_declaration5823 specparam_declaration_instance5823();
    specparam_declaration5824 specparam_declaration_instance5824();
    specparam_declaration5825 specparam_declaration_instance5825();
    specparam_declaration5826 specparam_declaration_instance5826();
    specparam_declaration5827 specparam_declaration_instance5827();
    specparam_declaration5828 specparam_declaration_instance5828();
    specparam_declaration5829 specparam_declaration_instance5829();
    specparam_declaration5830 specparam_declaration_instance5830();
    specparam_declaration5831 specparam_declaration_instance5831();
    specparam_declaration5832 specparam_declaration_instance5832();
    specparam_declaration5833 specparam_declaration_instance5833();
    specparam_declaration5834 specparam_declaration_instance5834();
    specparam_declaration5835 specparam_declaration_instance5835();
    specparam_declaration5836 specparam_declaration_instance5836();
    specparam_declaration5837 specparam_declaration_instance5837();
    specparam_declaration5838 specparam_declaration_instance5838();
    specparam_declaration5839 specparam_declaration_instance5839();
    specparam_declaration5840 specparam_declaration_instance5840();
    specparam_declaration5841 specparam_declaration_instance5841();
    specparam_declaration5842 specparam_declaration_instance5842();
    specparam_declaration5843 specparam_declaration_instance5843();
    specparam_declaration5844 specparam_declaration_instance5844();
    specparam_declaration5845 specparam_declaration_instance5845();
    specparam_declaration5846 specparam_declaration_instance5846();
    specparam_declaration5847 specparam_declaration_instance5847();
    specparam_declaration5848 specparam_declaration_instance5848();
    specparam_declaration5849 specparam_declaration_instance5849();
    specparam_declaration5850 specparam_declaration_instance5850();
    specparam_declaration5851 specparam_declaration_instance5851();
    specparam_declaration5852 specparam_declaration_instance5852();
    specparam_declaration5853 specparam_declaration_instance5853();
    specparam_declaration5854 specparam_declaration_instance5854();
    specparam_declaration5855 specparam_declaration_instance5855();
    specparam_declaration5856 specparam_declaration_instance5856();
    specparam_declaration5857 specparam_declaration_instance5857();
    specparam_declaration5858 specparam_declaration_instance5858();
    specparam_declaration5859 specparam_declaration_instance5859();
    specparam_declaration5860 specparam_declaration_instance5860();
    specparam_declaration5861 specparam_declaration_instance5861();
    specparam_declaration5862 specparam_declaration_instance5862();
    specparam_declaration5863 specparam_declaration_instance5863();
    specparam_declaration5864 specparam_declaration_instance5864();
    specparam_declaration5865 specparam_declaration_instance5865();
    specparam_declaration5866 specparam_declaration_instance5866();
    specparam_declaration5867 specparam_declaration_instance5867();
    specparam_declaration5868 specparam_declaration_instance5868();
    specparam_declaration5869 specparam_declaration_instance5869();
    specparam_declaration5870 specparam_declaration_instance5870();
    specparam_declaration5871 specparam_declaration_instance5871();
    specparam_declaration5872 specparam_declaration_instance5872();
    specparam_declaration5873 specparam_declaration_instance5873();
    specparam_declaration5874 specparam_declaration_instance5874();
    specparam_declaration5875 specparam_declaration_instance5875();
    specparam_declaration5876 specparam_declaration_instance5876();
    specparam_declaration5877 specparam_declaration_instance5877();
    specparam_declaration5878 specparam_declaration_instance5878();
    specparam_declaration5879 specparam_declaration_instance5879();
    specparam_declaration5880 specparam_declaration_instance5880();
    specparam_declaration5881 specparam_declaration_instance5881();
    specparam_declaration5882 specparam_declaration_instance5882();
    specparam_declaration5883 specparam_declaration_instance5883();
    specparam_declaration5884 specparam_declaration_instance5884();
    specparam_declaration5885 specparam_declaration_instance5885();
    specparam_declaration5886 specparam_declaration_instance5886();
    specparam_declaration5887 specparam_declaration_instance5887();
    specparam_declaration5888 specparam_declaration_instance5888();
    specparam_declaration5889 specparam_declaration_instance5889();
    specparam_declaration5890 specparam_declaration_instance5890();
    specparam_declaration5891 specparam_declaration_instance5891();
    specparam_declaration5892 specparam_declaration_instance5892();
    specparam_declaration5893 specparam_declaration_instance5893();
    specparam_declaration5894 specparam_declaration_instance5894();
    specparam_declaration5895 specparam_declaration_instance5895();
    specparam_declaration5896 specparam_declaration_instance5896();
    specparam_declaration5897 specparam_declaration_instance5897();
    specparam_declaration5898 specparam_declaration_instance5898();
    specparam_declaration5899 specparam_declaration_instance5899();
    specparam_declaration5900 specparam_declaration_instance5900();
    specparam_declaration5901 specparam_declaration_instance5901();
    specparam_declaration5902 specparam_declaration_instance5902();
    specparam_declaration5903 specparam_declaration_instance5903();
    specparam_declaration5904 specparam_declaration_instance5904();
    specparam_declaration5905 specparam_declaration_instance5905();
    specparam_declaration5906 specparam_declaration_instance5906();
    specparam_declaration5907 specparam_declaration_instance5907();
    specparam_declaration5908 specparam_declaration_instance5908();
    specparam_declaration5909 specparam_declaration_instance5909();
    specparam_declaration5910 specparam_declaration_instance5910();
    specparam_declaration5911 specparam_declaration_instance5911();
    specparam_declaration5912 specparam_declaration_instance5912();
    specparam_declaration5913 specparam_declaration_instance5913();
    specparam_declaration5914 specparam_declaration_instance5914();
    specparam_declaration5915 specparam_declaration_instance5915();
    specparam_declaration5916 specparam_declaration_instance5916();
    specparam_declaration5917 specparam_declaration_instance5917();
    specparam_declaration5918 specparam_declaration_instance5918();
    specparam_declaration5919 specparam_declaration_instance5919();
    specparam_declaration5920 specparam_declaration_instance5920();
    specparam_declaration5921 specparam_declaration_instance5921();
    specparam_declaration5922 specparam_declaration_instance5922();
    specparam_declaration5923 specparam_declaration_instance5923();
    specparam_declaration5924 specparam_declaration_instance5924();
    specparam_declaration5925 specparam_declaration_instance5925();
    specparam_declaration5926 specparam_declaration_instance5926();
    specparam_declaration5927 specparam_declaration_instance5927();
    specparam_declaration5928 specparam_declaration_instance5928();
    specparam_declaration5929 specparam_declaration_instance5929();
    specparam_declaration5930 specparam_declaration_instance5930();
    specparam_declaration5931 specparam_declaration_instance5931();
    specparam_declaration5932 specparam_declaration_instance5932();
    specparam_declaration5933 specparam_declaration_instance5933();
    specparam_declaration5934 specparam_declaration_instance5934();
    specparam_declaration5935 specparam_declaration_instance5935();
    specparam_declaration5936 specparam_declaration_instance5936();
    specparam_declaration5937 specparam_declaration_instance5937();
    specparam_declaration5938 specparam_declaration_instance5938();
    specparam_declaration5939 specparam_declaration_instance5939();
    specparam_declaration5940 specparam_declaration_instance5940();
    specparam_declaration5941 specparam_declaration_instance5941();
    specparam_declaration5942 specparam_declaration_instance5942();
    specparam_declaration5943 specparam_declaration_instance5943();
    specparam_declaration5944 specparam_declaration_instance5944();
    specparam_declaration5945 specparam_declaration_instance5945();
    specparam_declaration5946 specparam_declaration_instance5946();
    specparam_declaration5947 specparam_declaration_instance5947();
    specparam_declaration5948 specparam_declaration_instance5948();
    specparam_declaration5949 specparam_declaration_instance5949();
    specparam_declaration5950 specparam_declaration_instance5950();
    specparam_declaration5951 specparam_declaration_instance5951();
    specparam_declaration5952 specparam_declaration_instance5952();
    specparam_declaration5953 specparam_declaration_instance5953();
    specparam_declaration5954 specparam_declaration_instance5954();
    specparam_declaration5955 specparam_declaration_instance5955();
    specparam_declaration5956 specparam_declaration_instance5956();
    specparam_declaration5957 specparam_declaration_instance5957();
    specparam_declaration5958 specparam_declaration_instance5958();
    specparam_declaration5959 specparam_declaration_instance5959();
    specparam_declaration5960 specparam_declaration_instance5960();
    specparam_declaration5961 specparam_declaration_instance5961();
    specparam_declaration5962 specparam_declaration_instance5962();
    specparam_declaration5963 specparam_declaration_instance5963();
    specparam_declaration5964 specparam_declaration_instance5964();
    specparam_declaration5965 specparam_declaration_instance5965();
    specparam_declaration5966 specparam_declaration_instance5966();
    specparam_declaration5967 specparam_declaration_instance5967();
    specparam_declaration5968 specparam_declaration_instance5968();
    specparam_declaration5969 specparam_declaration_instance5969();
    specparam_declaration5970 specparam_declaration_instance5970();
    specparam_declaration5971 specparam_declaration_instance5971();
    specparam_declaration5972 specparam_declaration_instance5972();
    specparam_declaration5973 specparam_declaration_instance5973();
    specparam_declaration5974 specparam_declaration_instance5974();
    specparam_declaration5975 specparam_declaration_instance5975();
    specparam_declaration5976 specparam_declaration_instance5976();
    specparam_declaration5977 specparam_declaration_instance5977();
    specparam_declaration5978 specparam_declaration_instance5978();
    specparam_declaration5979 specparam_declaration_instance5979();
    specparam_declaration5980 specparam_declaration_instance5980();
    specparam_declaration5981 specparam_declaration_instance5981();
    specparam_declaration5982 specparam_declaration_instance5982();
    specparam_declaration5983 specparam_declaration_instance5983();
    specparam_declaration5984 specparam_declaration_instance5984();
    specparam_declaration5985 specparam_declaration_instance5985();
    specparam_declaration5986 specparam_declaration_instance5986();
    specparam_declaration5987 specparam_declaration_instance5987();
    specparam_declaration5988 specparam_declaration_instance5988();
    specparam_declaration5989 specparam_declaration_instance5989();
    specparam_declaration5990 specparam_declaration_instance5990();
    specparam_declaration5991 specparam_declaration_instance5991();
    specparam_declaration5992 specparam_declaration_instance5992();
    specparam_declaration5993 specparam_declaration_instance5993();
    specparam_declaration5994 specparam_declaration_instance5994();
    specparam_declaration5995 specparam_declaration_instance5995();
    specparam_declaration5996 specparam_declaration_instance5996();
    specparam_declaration5997 specparam_declaration_instance5997();
    specparam_declaration5998 specparam_declaration_instance5998();
    specparam_declaration5999 specparam_declaration_instance5999();
    specparam_declaration6000 specparam_declaration_instance6000();
    specparam_declaration6001 specparam_declaration_instance6001();
    specparam_declaration6002 specparam_declaration_instance6002();
    specparam_declaration6003 specparam_declaration_instance6003();
    specparam_declaration6004 specparam_declaration_instance6004();
    specparam_declaration6005 specparam_declaration_instance6005();
    specparam_declaration6006 specparam_declaration_instance6006();
    specparam_declaration6007 specparam_declaration_instance6007();
    specparam_declaration6008 specparam_declaration_instance6008();
    specparam_declaration6009 specparam_declaration_instance6009();
    specparam_declaration6010 specparam_declaration_instance6010();
    specparam_declaration6011 specparam_declaration_instance6011();
    specparam_declaration6012 specparam_declaration_instance6012();
    specparam_declaration6013 specparam_declaration_instance6013();
    specparam_declaration6014 specparam_declaration_instance6014();
    specparam_declaration6015 specparam_declaration_instance6015();
    specparam_declaration6016 specparam_declaration_instance6016();
    specparam_declaration6017 specparam_declaration_instance6017();
    specparam_declaration6018 specparam_declaration_instance6018();
    specparam_declaration6019 specparam_declaration_instance6019();
    specparam_declaration6020 specparam_declaration_instance6020();
    specparam_declaration6021 specparam_declaration_instance6021();
    specparam_declaration6022 specparam_declaration_instance6022();
    specparam_declaration6023 specparam_declaration_instance6023();
    specparam_declaration6024 specparam_declaration_instance6024();
    specparam_declaration6025 specparam_declaration_instance6025();
    specparam_declaration6026 specparam_declaration_instance6026();
    specparam_declaration6027 specparam_declaration_instance6027();
    specparam_declaration6028 specparam_declaration_instance6028();
    specparam_declaration6029 specparam_declaration_instance6029();
    specparam_declaration6030 specparam_declaration_instance6030();
    specparam_declaration6031 specparam_declaration_instance6031();
    specparam_declaration6032 specparam_declaration_instance6032();
    specparam_declaration6033 specparam_declaration_instance6033();
    specparam_declaration6034 specparam_declaration_instance6034();
    specparam_declaration6035 specparam_declaration_instance6035();
    specparam_declaration6036 specparam_declaration_instance6036();
    specparam_declaration6037 specparam_declaration_instance6037();
    specparam_declaration6038 specparam_declaration_instance6038();
    specparam_declaration6039 specparam_declaration_instance6039();
    specparam_declaration6040 specparam_declaration_instance6040();
    specparam_declaration6041 specparam_declaration_instance6041();
    specparam_declaration6042 specparam_declaration_instance6042();
    specparam_declaration6043 specparam_declaration_instance6043();
    specparam_declaration6044 specparam_declaration_instance6044();
    specparam_declaration6045 specparam_declaration_instance6045();
    specparam_declaration6046 specparam_declaration_instance6046();
    specparam_declaration6047 specparam_declaration_instance6047();
    specparam_declaration6048 specparam_declaration_instance6048();
    specparam_declaration6049 specparam_declaration_instance6049();
    specparam_declaration6050 specparam_declaration_instance6050();
    specparam_declaration6051 specparam_declaration_instance6051();
    specparam_declaration6052 specparam_declaration_instance6052();
    specparam_declaration6053 specparam_declaration_instance6053();
    specparam_declaration6054 specparam_declaration_instance6054();
    specparam_declaration6055 specparam_declaration_instance6055();
    specparam_declaration6056 specparam_declaration_instance6056();
    specparam_declaration6057 specparam_declaration_instance6057();
    specparam_declaration6058 specparam_declaration_instance6058();
    specparam_declaration6059 specparam_declaration_instance6059();
    specparam_declaration6060 specparam_declaration_instance6060();
    specparam_declaration6061 specparam_declaration_instance6061();
    specparam_declaration6062 specparam_declaration_instance6062();
    specparam_declaration6063 specparam_declaration_instance6063();
    specparam_declaration6064 specparam_declaration_instance6064();
    specparam_declaration6065 specparam_declaration_instance6065();
    specparam_declaration6066 specparam_declaration_instance6066();
    specparam_declaration6067 specparam_declaration_instance6067();
    specparam_declaration6068 specparam_declaration_instance6068();
    specparam_declaration6069 specparam_declaration_instance6069();
    specparam_declaration6070 specparam_declaration_instance6070();
    specparam_declaration6071 specparam_declaration_instance6071();
    specparam_declaration6072 specparam_declaration_instance6072();
    specparam_declaration6073 specparam_declaration_instance6073();
    specparam_declaration6074 specparam_declaration_instance6074();
    specparam_declaration6075 specparam_declaration_instance6075();
    specparam_declaration6076 specparam_declaration_instance6076();
    specparam_declaration6077 specparam_declaration_instance6077();
    specparam_declaration6078 specparam_declaration_instance6078();
    specparam_declaration6079 specparam_declaration_instance6079();
    specparam_declaration6080 specparam_declaration_instance6080();
    specparam_declaration6081 specparam_declaration_instance6081();
    specparam_declaration6082 specparam_declaration_instance6082();
    specparam_declaration6083 specparam_declaration_instance6083();
    specparam_declaration6084 specparam_declaration_instance6084();
    specparam_declaration6085 specparam_declaration_instance6085();
    specparam_declaration6086 specparam_declaration_instance6086();
    specparam_declaration6087 specparam_declaration_instance6087();
    specparam_declaration6088 specparam_declaration_instance6088();
    specparam_declaration6089 specparam_declaration_instance6089();
    specparam_declaration6090 specparam_declaration_instance6090();
    specparam_declaration6091 specparam_declaration_instance6091();
    specparam_declaration6092 specparam_declaration_instance6092();
    specparam_declaration6093 specparam_declaration_instance6093();
    specparam_declaration6094 specparam_declaration_instance6094();
    specparam_declaration6095 specparam_declaration_instance6095();
    specparam_declaration6096 specparam_declaration_instance6096();
    specparam_declaration6097 specparam_declaration_instance6097();
    specparam_declaration6098 specparam_declaration_instance6098();
    specparam_declaration6099 specparam_declaration_instance6099();
    specparam_declaration6100 specparam_declaration_instance6100();
    specparam_declaration6101 specparam_declaration_instance6101();
    specparam_declaration6102 specparam_declaration_instance6102();
    specparam_declaration6103 specparam_declaration_instance6103();
    specparam_declaration6104 specparam_declaration_instance6104();
    specparam_declaration6105 specparam_declaration_instance6105();
    specparam_declaration6106 specparam_declaration_instance6106();
    specparam_declaration6107 specparam_declaration_instance6107();
    specparam_declaration6108 specparam_declaration_instance6108();
    specparam_declaration6109 specparam_declaration_instance6109();
    specparam_declaration6110 specparam_declaration_instance6110();
    specparam_declaration6111 specparam_declaration_instance6111();
    specparam_declaration6112 specparam_declaration_instance6112();
    specparam_declaration6113 specparam_declaration_instance6113();
    specparam_declaration6114 specparam_declaration_instance6114();
    specparam_declaration6115 specparam_declaration_instance6115();
    specparam_declaration6116 specparam_declaration_instance6116();
    specparam_declaration6117 specparam_declaration_instance6117();
    specparam_declaration6118 specparam_declaration_instance6118();
    specparam_declaration6119 specparam_declaration_instance6119();
    specparam_declaration6120 specparam_declaration_instance6120();
    specparam_declaration6121 specparam_declaration_instance6121();
    specparam_declaration6122 specparam_declaration_instance6122();
    specparam_declaration6123 specparam_declaration_instance6123();
    specparam_declaration6124 specparam_declaration_instance6124();
    specparam_declaration6125 specparam_declaration_instance6125();
    specparam_declaration6126 specparam_declaration_instance6126();
    specparam_declaration6127 specparam_declaration_instance6127();
    specparam_declaration6128 specparam_declaration_instance6128();
    specparam_declaration6129 specparam_declaration_instance6129();
    specparam_declaration6130 specparam_declaration_instance6130();
    specparam_declaration6131 specparam_declaration_instance6131();
    specparam_declaration6132 specparam_declaration_instance6132();
    specparam_declaration6133 specparam_declaration_instance6133();
    specparam_declaration6134 specparam_declaration_instance6134();
    specparam_declaration6135 specparam_declaration_instance6135();
    specparam_declaration6136 specparam_declaration_instance6136();
    specparam_declaration6137 specparam_declaration_instance6137();
    specparam_declaration6138 specparam_declaration_instance6138();
    specparam_declaration6139 specparam_declaration_instance6139();
    specparam_declaration6140 specparam_declaration_instance6140();
    specparam_declaration6141 specparam_declaration_instance6141();
    specparam_declaration6142 specparam_declaration_instance6142();
    specparam_declaration6143 specparam_declaration_instance6143();
    specparam_declaration6144 specparam_declaration_instance6144();
    specparam_declaration6145 specparam_declaration_instance6145();
    specparam_declaration6146 specparam_declaration_instance6146();
    specparam_declaration6147 specparam_declaration_instance6147();
    specparam_declaration6148 specparam_declaration_instance6148();
    specparam_declaration6149 specparam_declaration_instance6149();
    specparam_declaration6150 specparam_declaration_instance6150();
    specparam_declaration6151 specparam_declaration_instance6151();
    specparam_declaration6152 specparam_declaration_instance6152();
    specparam_declaration6153 specparam_declaration_instance6153();
    specparam_declaration6154 specparam_declaration_instance6154();
    specparam_declaration6155 specparam_declaration_instance6155();
    specparam_declaration6156 specparam_declaration_instance6156();
    specparam_declaration6157 specparam_declaration_instance6157();
    specparam_declaration6158 specparam_declaration_instance6158();
    specparam_declaration6159 specparam_declaration_instance6159();
    specparam_declaration6160 specparam_declaration_instance6160();
    specparam_declaration6161 specparam_declaration_instance6161();
    specparam_declaration6162 specparam_declaration_instance6162();
    specparam_declaration6163 specparam_declaration_instance6163();
    specparam_declaration6164 specparam_declaration_instance6164();
    specparam_declaration6165 specparam_declaration_instance6165();
    specparam_declaration6166 specparam_declaration_instance6166();
    specparam_declaration6167 specparam_declaration_instance6167();
    specparam_declaration6168 specparam_declaration_instance6168();
    specparam_declaration6169 specparam_declaration_instance6169();
    specparam_declaration6170 specparam_declaration_instance6170();
    specparam_declaration6171 specparam_declaration_instance6171();
    specparam_declaration6172 specparam_declaration_instance6172();
    specparam_declaration6173 specparam_declaration_instance6173();
    specparam_declaration6174 specparam_declaration_instance6174();
    specparam_declaration6175 specparam_declaration_instance6175();
    specparam_declaration6176 specparam_declaration_instance6176();
    specparam_declaration6177 specparam_declaration_instance6177();
    specparam_declaration6178 specparam_declaration_instance6178();
    specparam_declaration6179 specparam_declaration_instance6179();
    specparam_declaration6180 specparam_declaration_instance6180();
    specparam_declaration6181 specparam_declaration_instance6181();
    specparam_declaration6182 specparam_declaration_instance6182();
    specparam_declaration6183 specparam_declaration_instance6183();
    specparam_declaration6184 specparam_declaration_instance6184();
    specparam_declaration6185 specparam_declaration_instance6185();
    specparam_declaration6186 specparam_declaration_instance6186();
    specparam_declaration6187 specparam_declaration_instance6187();
    specparam_declaration6188 specparam_declaration_instance6188();
    specparam_declaration6189 specparam_declaration_instance6189();
    specparam_declaration6190 specparam_declaration_instance6190();
    specparam_declaration6191 specparam_declaration_instance6191();
    specparam_declaration6192 specparam_declaration_instance6192();
    specparam_declaration6193 specparam_declaration_instance6193();
    specparam_declaration6194 specparam_declaration_instance6194();
    specparam_declaration6195 specparam_declaration_instance6195();
    specparam_declaration6196 specparam_declaration_instance6196();
    specparam_declaration6197 specparam_declaration_instance6197();
    specparam_declaration6198 specparam_declaration_instance6198();
    specparam_declaration6199 specparam_declaration_instance6199();
    specparam_declaration6200 specparam_declaration_instance6200();
    specparam_declaration6201 specparam_declaration_instance6201();
    specparam_declaration6202 specparam_declaration_instance6202();
    specparam_declaration6203 specparam_declaration_instance6203();
    specparam_declaration6204 specparam_declaration_instance6204();
    specparam_declaration6205 specparam_declaration_instance6205();
    specparam_declaration6206 specparam_declaration_instance6206();
    specparam_declaration6207 specparam_declaration_instance6207();
    specparam_declaration6208 specparam_declaration_instance6208();
    specparam_declaration6209 specparam_declaration_instance6209();
    specparam_declaration6210 specparam_declaration_instance6210();
    specparam_declaration6211 specparam_declaration_instance6211();
    specparam_declaration6212 specparam_declaration_instance6212();
    specparam_declaration6213 specparam_declaration_instance6213();
    specparam_declaration6214 specparam_declaration_instance6214();
    specparam_declaration6215 specparam_declaration_instance6215();
    specparam_declaration6216 specparam_declaration_instance6216();
    specparam_declaration6217 specparam_declaration_instance6217();
    specparam_declaration6218 specparam_declaration_instance6218();
    specparam_declaration6219 specparam_declaration_instance6219();
    specparam_declaration6220 specparam_declaration_instance6220();
    specparam_declaration6221 specparam_declaration_instance6221();
    specparam_declaration6222 specparam_declaration_instance6222();
    specparam_declaration6223 specparam_declaration_instance6223();
    specparam_declaration6224 specparam_declaration_instance6224();
    specparam_declaration6225 specparam_declaration_instance6225();
    specparam_declaration6226 specparam_declaration_instance6226();
    specparam_declaration6227 specparam_declaration_instance6227();
    specparam_declaration6228 specparam_declaration_instance6228();
    specparam_declaration6229 specparam_declaration_instance6229();
    specparam_declaration6230 specparam_declaration_instance6230();
    specparam_declaration6231 specparam_declaration_instance6231();
    specparam_declaration6232 specparam_declaration_instance6232();
    specparam_declaration6233 specparam_declaration_instance6233();
    specparam_declaration6234 specparam_declaration_instance6234();
    specparam_declaration6235 specparam_declaration_instance6235();
    specparam_declaration6236 specparam_declaration_instance6236();
    specparam_declaration6237 specparam_declaration_instance6237();
    specparam_declaration6238 specparam_declaration_instance6238();
    specparam_declaration6239 specparam_declaration_instance6239();
    specparam_declaration6240 specparam_declaration_instance6240();
    specparam_declaration6241 specparam_declaration_instance6241();
    specparam_declaration6242 specparam_declaration_instance6242();
    specparam_declaration6243 specparam_declaration_instance6243();
    specparam_declaration6244 specparam_declaration_instance6244();
    specparam_declaration6245 specparam_declaration_instance6245();
    specparam_declaration6246 specparam_declaration_instance6246();
    specparam_declaration6247 specparam_declaration_instance6247();
    specparam_declaration6248 specparam_declaration_instance6248();
    specparam_declaration6249 specparam_declaration_instance6249();
    specparam_declaration6250 specparam_declaration_instance6250();
    specparam_declaration6251 specparam_declaration_instance6251();
    specparam_declaration6252 specparam_declaration_instance6252();
    specparam_declaration6253 specparam_declaration_instance6253();
    specparam_declaration6254 specparam_declaration_instance6254();
    specparam_declaration6255 specparam_declaration_instance6255();
    specparam_declaration6256 specparam_declaration_instance6256();
    specparam_declaration6257 specparam_declaration_instance6257();
    specparam_declaration6258 specparam_declaration_instance6258();
    specparam_declaration6259 specparam_declaration_instance6259();
    specparam_declaration6260 specparam_declaration_instance6260();
    specparam_declaration6261 specparam_declaration_instance6261();
    specparam_declaration6262 specparam_declaration_instance6262();
    specparam_declaration6263 specparam_declaration_instance6263();
    specparam_declaration6264 specparam_declaration_instance6264();
    specparam_declaration6265 specparam_declaration_instance6265();
    specparam_declaration6266 specparam_declaration_instance6266();
    specparam_declaration6267 specparam_declaration_instance6267();
    specparam_declaration6268 specparam_declaration_instance6268();
    specparam_declaration6269 specparam_declaration_instance6269();
    specparam_declaration6270 specparam_declaration_instance6270();
    specparam_declaration6271 specparam_declaration_instance6271();
    specparam_declaration6272 specparam_declaration_instance6272();
    specparam_declaration6273 specparam_declaration_instance6273();
    specparam_declaration6274 specparam_declaration_instance6274();
    specparam_declaration6275 specparam_declaration_instance6275();
    specparam_declaration6276 specparam_declaration_instance6276();
    specparam_declaration6277 specparam_declaration_instance6277();
    specparam_declaration6278 specparam_declaration_instance6278();
    specparam_declaration6279 specparam_declaration_instance6279();
    specparam_declaration6280 specparam_declaration_instance6280();
    specparam_declaration6281 specparam_declaration_instance6281();
    specparam_declaration6282 specparam_declaration_instance6282();
    specparam_declaration6283 specparam_declaration_instance6283();
    specparam_declaration6284 specparam_declaration_instance6284();
    specparam_declaration6285 specparam_declaration_instance6285();
    specparam_declaration6286 specparam_declaration_instance6286();
    specparam_declaration6287 specparam_declaration_instance6287();
    specparam_declaration6288 specparam_declaration_instance6288();
    specparam_declaration6289 specparam_declaration_instance6289();
    specparam_declaration6290 specparam_declaration_instance6290();
    specparam_declaration6291 specparam_declaration_instance6291();
    specparam_declaration6292 specparam_declaration_instance6292();
    specparam_declaration6293 specparam_declaration_instance6293();
    specparam_declaration6294 specparam_declaration_instance6294();
    specparam_declaration6295 specparam_declaration_instance6295();
    specparam_declaration6296 specparam_declaration_instance6296();
    specparam_declaration6297 specparam_declaration_instance6297();
    specparam_declaration6298 specparam_declaration_instance6298();
    specparam_declaration6299 specparam_declaration_instance6299();
    specparam_declaration6300 specparam_declaration_instance6300();
    specparam_declaration6301 specparam_declaration_instance6301();
    specparam_declaration6302 specparam_declaration_instance6302();
    specparam_declaration6303 specparam_declaration_instance6303();
    specparam_declaration6304 specparam_declaration_instance6304();
    specparam_declaration6305 specparam_declaration_instance6305();
    specparam_declaration6306 specparam_declaration_instance6306();
    specparam_declaration6307 specparam_declaration_instance6307();
    specparam_declaration6308 specparam_declaration_instance6308();
    specparam_declaration6309 specparam_declaration_instance6309();
    specparam_declaration6310 specparam_declaration_instance6310();
    specparam_declaration6311 specparam_declaration_instance6311();
    specparam_declaration6312 specparam_declaration_instance6312();
    specparam_declaration6313 specparam_declaration_instance6313();
    specparam_declaration6314 specparam_declaration_instance6314();
    specparam_declaration6315 specparam_declaration_instance6315();
    specparam_declaration6316 specparam_declaration_instance6316();
    specparam_declaration6317 specparam_declaration_instance6317();
    specparam_declaration6318 specparam_declaration_instance6318();
    specparam_declaration6319 specparam_declaration_instance6319();
    specparam_declaration6320 specparam_declaration_instance6320();
    specparam_declaration6321 specparam_declaration_instance6321();
    specparam_declaration6322 specparam_declaration_instance6322();
    specparam_declaration6323 specparam_declaration_instance6323();
    specparam_declaration6324 specparam_declaration_instance6324();
    specparam_declaration6325 specparam_declaration_instance6325();
    specparam_declaration6326 specparam_declaration_instance6326();
    specparam_declaration6327 specparam_declaration_instance6327();
    specparam_declaration6328 specparam_declaration_instance6328();
    specparam_declaration6329 specparam_declaration_instance6329();
    specparam_declaration6330 specparam_declaration_instance6330();
    specparam_declaration6331 specparam_declaration_instance6331();
    specparam_declaration6332 specparam_declaration_instance6332();
    specparam_declaration6333 specparam_declaration_instance6333();
    specparam_declaration6334 specparam_declaration_instance6334();
    specparam_declaration6335 specparam_declaration_instance6335();
    specparam_declaration6336 specparam_declaration_instance6336();
    specparam_declaration6337 specparam_declaration_instance6337();
    specparam_declaration6338 specparam_declaration_instance6338();
    specparam_declaration6339 specparam_declaration_instance6339();
    specparam_declaration6340 specparam_declaration_instance6340();
    specparam_declaration6341 specparam_declaration_instance6341();
    specparam_declaration6342 specparam_declaration_instance6342();
    specparam_declaration6343 specparam_declaration_instance6343();
    specparam_declaration6344 specparam_declaration_instance6344();
    specparam_declaration6345 specparam_declaration_instance6345();
    specparam_declaration6346 specparam_declaration_instance6346();
    specparam_declaration6347 specparam_declaration_instance6347();
    specparam_declaration6348 specparam_declaration_instance6348();
    specparam_declaration6349 specparam_declaration_instance6349();
    specparam_declaration6350 specparam_declaration_instance6350();
    specparam_declaration6351 specparam_declaration_instance6351();
    specparam_declaration6352 specparam_declaration_instance6352();
    specparam_declaration6353 specparam_declaration_instance6353();
    specparam_declaration6354 specparam_declaration_instance6354();
    specparam_declaration6355 specparam_declaration_instance6355();
    specparam_declaration6356 specparam_declaration_instance6356();
    specparam_declaration6357 specparam_declaration_instance6357();
    specparam_declaration6358 specparam_declaration_instance6358();
    specparam_declaration6359 specparam_declaration_instance6359();
    specparam_declaration6360 specparam_declaration_instance6360();
    specparam_declaration6361 specparam_declaration_instance6361();
    specparam_declaration6362 specparam_declaration_instance6362();
    specparam_declaration6363 specparam_declaration_instance6363();
    specparam_declaration6364 specparam_declaration_instance6364();
    specparam_declaration6365 specparam_declaration_instance6365();
    specparam_declaration6366 specparam_declaration_instance6366();
    specparam_declaration6367 specparam_declaration_instance6367();
    specparam_declaration6368 specparam_declaration_instance6368();
    specparam_declaration6369 specparam_declaration_instance6369();
    specparam_declaration6370 specparam_declaration_instance6370();
    specparam_declaration6371 specparam_declaration_instance6371();
    specparam_declaration6372 specparam_declaration_instance6372();
    specparam_declaration6373 specparam_declaration_instance6373();
    specparam_declaration6374 specparam_declaration_instance6374();
    specparam_declaration6375 specparam_declaration_instance6375();
    specparam_declaration6376 specparam_declaration_instance6376();
    specparam_declaration6377 specparam_declaration_instance6377();
    specparam_declaration6378 specparam_declaration_instance6378();
    specparam_declaration6379 specparam_declaration_instance6379();
    specparam_declaration6380 specparam_declaration_instance6380();
    specparam_declaration6381 specparam_declaration_instance6381();
    specparam_declaration6382 specparam_declaration_instance6382();
    specparam_declaration6383 specparam_declaration_instance6383();
    specparam_declaration6384 specparam_declaration_instance6384();
    specparam_declaration6385 specparam_declaration_instance6385();
    specparam_declaration6386 specparam_declaration_instance6386();
    specparam_declaration6387 specparam_declaration_instance6387();
    specparam_declaration6388 specparam_declaration_instance6388();
    specparam_declaration6389 specparam_declaration_instance6389();
    specparam_declaration6390 specparam_declaration_instance6390();
    specparam_declaration6391 specparam_declaration_instance6391();
    specparam_declaration6392 specparam_declaration_instance6392();
    specparam_declaration6393 specparam_declaration_instance6393();
    specparam_declaration6394 specparam_declaration_instance6394();
    specparam_declaration6395 specparam_declaration_instance6395();
    specparam_declaration6396 specparam_declaration_instance6396();
    specparam_declaration6397 specparam_declaration_instance6397();
    specparam_declaration6398 specparam_declaration_instance6398();
    specparam_declaration6399 specparam_declaration_instance6399();
    specparam_declaration6400 specparam_declaration_instance6400();
    specparam_declaration6401 specparam_declaration_instance6401();
    specparam_declaration6402 specparam_declaration_instance6402();
    specparam_declaration6403 specparam_declaration_instance6403();
    specparam_declaration6404 specparam_declaration_instance6404();
    specparam_declaration6405 specparam_declaration_instance6405();
    specparam_declaration6406 specparam_declaration_instance6406();
    specparam_declaration6407 specparam_declaration_instance6407();
    specparam_declaration6408 specparam_declaration_instance6408();
    specparam_declaration6409 specparam_declaration_instance6409();
    specparam_declaration6410 specparam_declaration_instance6410();
    specparam_declaration6411 specparam_declaration_instance6411();
    specparam_declaration6412 specparam_declaration_instance6412();
    specparam_declaration6413 specparam_declaration_instance6413();
    specparam_declaration6414 specparam_declaration_instance6414();
    specparam_declaration6415 specparam_declaration_instance6415();
    specparam_declaration6416 specparam_declaration_instance6416();
    specparam_declaration6417 specparam_declaration_instance6417();
    specparam_declaration6418 specparam_declaration_instance6418();
    specparam_declaration6419 specparam_declaration_instance6419();
    specparam_declaration6420 specparam_declaration_instance6420();
    specparam_declaration6421 specparam_declaration_instance6421();
    specparam_declaration6422 specparam_declaration_instance6422();
    specparam_declaration6423 specparam_declaration_instance6423();
    specparam_declaration6424 specparam_declaration_instance6424();
    specparam_declaration6425 specparam_declaration_instance6425();
    specparam_declaration6426 specparam_declaration_instance6426();
    specparam_declaration6427 specparam_declaration_instance6427();
    specparam_declaration6428 specparam_declaration_instance6428();
    specparam_declaration6429 specparam_declaration_instance6429();
    specparam_declaration6430 specparam_declaration_instance6430();
    specparam_declaration6431 specparam_declaration_instance6431();
    specparam_declaration6432 specparam_declaration_instance6432();
    specparam_declaration6433 specparam_declaration_instance6433();
    specparam_declaration6434 specparam_declaration_instance6434();
    specparam_declaration6435 specparam_declaration_instance6435();
    specparam_declaration6436 specparam_declaration_instance6436();
    specparam_declaration6437 specparam_declaration_instance6437();
    specparam_declaration6438 specparam_declaration_instance6438();
    specparam_declaration6439 specparam_declaration_instance6439();
    specparam_declaration6440 specparam_declaration_instance6440();
    specparam_declaration6441 specparam_declaration_instance6441();
    specparam_declaration6442 specparam_declaration_instance6442();
    specparam_declaration6443 specparam_declaration_instance6443();
    specparam_declaration6444 specparam_declaration_instance6444();
    specparam_declaration6445 specparam_declaration_instance6445();
    specparam_declaration6446 specparam_declaration_instance6446();
    specparam_declaration6447 specparam_declaration_instance6447();
    specparam_declaration6448 specparam_declaration_instance6448();
    specparam_declaration6449 specparam_declaration_instance6449();
    specparam_declaration6450 specparam_declaration_instance6450();
    specparam_declaration6451 specparam_declaration_instance6451();
    specparam_declaration6452 specparam_declaration_instance6452();
    specparam_declaration6453 specparam_declaration_instance6453();
    specparam_declaration6454 specparam_declaration_instance6454();
    specparam_declaration6455 specparam_declaration_instance6455();
    specparam_declaration6456 specparam_declaration_instance6456();
    specparam_declaration6457 specparam_declaration_instance6457();
    specparam_declaration6458 specparam_declaration_instance6458();
    specparam_declaration6459 specparam_declaration_instance6459();
    specparam_declaration6460 specparam_declaration_instance6460();
    specparam_declaration6461 specparam_declaration_instance6461();
    specparam_declaration6462 specparam_declaration_instance6462();
    specparam_declaration6463 specparam_declaration_instance6463();
    specparam_declaration6464 specparam_declaration_instance6464();
    specparam_declaration6465 specparam_declaration_instance6465();
    specparam_declaration6466 specparam_declaration_instance6466();
    specparam_declaration6467 specparam_declaration_instance6467();
    specparam_declaration6468 specparam_declaration_instance6468();
    specparam_declaration6469 specparam_declaration_instance6469();
    specparam_declaration6470 specparam_declaration_instance6470();
    specparam_declaration6471 specparam_declaration_instance6471();
    specparam_declaration6472 specparam_declaration_instance6472();
    specparam_declaration6473 specparam_declaration_instance6473();
    specparam_declaration6474 specparam_declaration_instance6474();
    specparam_declaration6475 specparam_declaration_instance6475();
    specparam_declaration6476 specparam_declaration_instance6476();
    specparam_declaration6477 specparam_declaration_instance6477();
    specparam_declaration6478 specparam_declaration_instance6478();
    specparam_declaration6479 specparam_declaration_instance6479();
    specparam_declaration6480 specparam_declaration_instance6480();
    specparam_declaration6481 specparam_declaration_instance6481();
    specparam_declaration6482 specparam_declaration_instance6482();
    specparam_declaration6483 specparam_declaration_instance6483();
    specparam_declaration6484 specparam_declaration_instance6484();
    specparam_declaration6485 specparam_declaration_instance6485();
    specparam_declaration6486 specparam_declaration_instance6486();
    specparam_declaration6487 specparam_declaration_instance6487();
    specparam_declaration6488 specparam_declaration_instance6488();
    specparam_declaration6489 specparam_declaration_instance6489();
    specparam_declaration6490 specparam_declaration_instance6490();
    specparam_declaration6491 specparam_declaration_instance6491();
    specparam_declaration6492 specparam_declaration_instance6492();
    specparam_declaration6493 specparam_declaration_instance6493();
    specparam_declaration6494 specparam_declaration_instance6494();
    specparam_declaration6495 specparam_declaration_instance6495();
    specparam_declaration6496 specparam_declaration_instance6496();
    specparam_declaration6497 specparam_declaration_instance6497();
    specparam_declaration6498 specparam_declaration_instance6498();
    specparam_declaration6499 specparam_declaration_instance6499();
    specparam_declaration6500 specparam_declaration_instance6500();
    specparam_declaration6501 specparam_declaration_instance6501();
    specparam_declaration6502 specparam_declaration_instance6502();
    specparam_declaration6503 specparam_declaration_instance6503();
    specparam_declaration6504 specparam_declaration_instance6504();
    specparam_declaration6505 specparam_declaration_instance6505();
    specparam_declaration6506 specparam_declaration_instance6506();
    specparam_declaration6507 specparam_declaration_instance6507();
    specparam_declaration6508 specparam_declaration_instance6508();
    specparam_declaration6509 specparam_declaration_instance6509();
    specparam_declaration6510 specparam_declaration_instance6510();
    specparam_declaration6511 specparam_declaration_instance6511();
    specparam_declaration6512 specparam_declaration_instance6512();
    specparam_declaration6513 specparam_declaration_instance6513();
    specparam_declaration6514 specparam_declaration_instance6514();
    specparam_declaration6515 specparam_declaration_instance6515();
    specparam_declaration6516 specparam_declaration_instance6516();
    specparam_declaration6517 specparam_declaration_instance6517();
    specparam_declaration6518 specparam_declaration_instance6518();
    specparam_declaration6519 specparam_declaration_instance6519();
    specparam_declaration6520 specparam_declaration_instance6520();
    specparam_declaration6521 specparam_declaration_instance6521();
    specparam_declaration6522 specparam_declaration_instance6522();
    specparam_declaration6523 specparam_declaration_instance6523();
    specparam_declaration6524 specparam_declaration_instance6524();
    specparam_declaration6525 specparam_declaration_instance6525();
    specparam_declaration6526 specparam_declaration_instance6526();
    specparam_declaration6527 specparam_declaration_instance6527();
    specparam_declaration6528 specparam_declaration_instance6528();
    specparam_declaration6529 specparam_declaration_instance6529();
    specparam_declaration6530 specparam_declaration_instance6530();
    specparam_declaration6531 specparam_declaration_instance6531();
    specparam_declaration6532 specparam_declaration_instance6532();
    specparam_declaration6533 specparam_declaration_instance6533();
    specparam_declaration6534 specparam_declaration_instance6534();
    specparam_declaration6535 specparam_declaration_instance6535();
    specparam_declaration6536 specparam_declaration_instance6536();
    specparam_declaration6537 specparam_declaration_instance6537();
    specparam_declaration6538 specparam_declaration_instance6538();
    specparam_declaration6539 specparam_declaration_instance6539();
    specparam_declaration6540 specparam_declaration_instance6540();
    specparam_declaration6541 specparam_declaration_instance6541();
    specparam_declaration6542 specparam_declaration_instance6542();
    specparam_declaration6543 specparam_declaration_instance6543();
    specparam_declaration6544 specparam_declaration_instance6544();
    specparam_declaration6545 specparam_declaration_instance6545();
    specparam_declaration6546 specparam_declaration_instance6546();
    specparam_declaration6547 specparam_declaration_instance6547();
    specparam_declaration6548 specparam_declaration_instance6548();
    specparam_declaration6549 specparam_declaration_instance6549();
    specparam_declaration6550 specparam_declaration_instance6550();
    specparam_declaration6551 specparam_declaration_instance6551();
    specparam_declaration6552 specparam_declaration_instance6552();
    specparam_declaration6553 specparam_declaration_instance6553();
    specparam_declaration6554 specparam_declaration_instance6554();
    specparam_declaration6555 specparam_declaration_instance6555();
    specparam_declaration6556 specparam_declaration_instance6556();
    specparam_declaration6557 specparam_declaration_instance6557();
    specparam_declaration6558 specparam_declaration_instance6558();
    specparam_declaration6559 specparam_declaration_instance6559();
    specparam_declaration6560 specparam_declaration_instance6560();
    specparam_declaration6561 specparam_declaration_instance6561();
    specparam_declaration6562 specparam_declaration_instance6562();
    specparam_declaration6563 specparam_declaration_instance6563();
    specparam_declaration6564 specparam_declaration_instance6564();
    specparam_declaration6565 specparam_declaration_instance6565();
    specparam_declaration6566 specparam_declaration_instance6566();
    specparam_declaration6567 specparam_declaration_instance6567();
    specparam_declaration6568 specparam_declaration_instance6568();
    specparam_declaration6569 specparam_declaration_instance6569();
    specparam_declaration6570 specparam_declaration_instance6570();
    specparam_declaration6571 specparam_declaration_instance6571();
    specparam_declaration6572 specparam_declaration_instance6572();
    specparam_declaration6573 specparam_declaration_instance6573();
    specparam_declaration6574 specparam_declaration_instance6574();
    specparam_declaration6575 specparam_declaration_instance6575();
    specparam_declaration6576 specparam_declaration_instance6576();
    specparam_declaration6577 specparam_declaration_instance6577();
    specparam_declaration6578 specparam_declaration_instance6578();
    specparam_declaration6579 specparam_declaration_instance6579();
    specparam_declaration6580 specparam_declaration_instance6580();
    specparam_declaration6581 specparam_declaration_instance6581();
    specparam_declaration6582 specparam_declaration_instance6582();
    specparam_declaration6583 specparam_declaration_instance6583();
    specparam_declaration6584 specparam_declaration_instance6584();
    specparam_declaration6585 specparam_declaration_instance6585();
    specparam_declaration6586 specparam_declaration_instance6586();
    specparam_declaration6587 specparam_declaration_instance6587();
    specparam_declaration6588 specparam_declaration_instance6588();
    specparam_declaration6589 specparam_declaration_instance6589();
    specparam_declaration6590 specparam_declaration_instance6590();
    specparam_declaration6591 specparam_declaration_instance6591();
    specparam_declaration6592 specparam_declaration_instance6592();
    specparam_declaration6593 specparam_declaration_instance6593();
    specparam_declaration6594 specparam_declaration_instance6594();
    specparam_declaration6595 specparam_declaration_instance6595();
    specparam_declaration6596 specparam_declaration_instance6596();
    specparam_declaration6597 specparam_declaration_instance6597();
    specparam_declaration6598 specparam_declaration_instance6598();
    specparam_declaration6599 specparam_declaration_instance6599();
    specparam_declaration6600 specparam_declaration_instance6600();
    specparam_declaration6601 specparam_declaration_instance6601();
    specparam_declaration6602 specparam_declaration_instance6602();
    specparam_declaration6603 specparam_declaration_instance6603();
    specparam_declaration6604 specparam_declaration_instance6604();
    specparam_declaration6605 specparam_declaration_instance6605();
    specparam_declaration6606 specparam_declaration_instance6606();
    specparam_declaration6607 specparam_declaration_instance6607();
    specparam_declaration6608 specparam_declaration_instance6608();
    specparam_declaration6609 specparam_declaration_instance6609();
    specparam_declaration6610 specparam_declaration_instance6610();
    specparam_declaration6611 specparam_declaration_instance6611();
    specparam_declaration6612 specparam_declaration_instance6612();
    specparam_declaration6613 specparam_declaration_instance6613();
    specparam_declaration6614 specparam_declaration_instance6614();
    specparam_declaration6615 specparam_declaration_instance6615();
    specparam_declaration6616 specparam_declaration_instance6616();
    specparam_declaration6617 specparam_declaration_instance6617();
    specparam_declaration6618 specparam_declaration_instance6618();
    specparam_declaration6619 specparam_declaration_instance6619();
    specparam_declaration6620 specparam_declaration_instance6620();
    specparam_declaration6621 specparam_declaration_instance6621();
    specparam_declaration6622 specparam_declaration_instance6622();
    specparam_declaration6623 specparam_declaration_instance6623();
    specparam_declaration6624 specparam_declaration_instance6624();
    specparam_declaration6625 specparam_declaration_instance6625();
    specparam_declaration6626 specparam_declaration_instance6626();
    specparam_declaration6627 specparam_declaration_instance6627();
    specparam_declaration6628 specparam_declaration_instance6628();
    specparam_declaration6629 specparam_declaration_instance6629();
    specparam_declaration6630 specparam_declaration_instance6630();
    specparam_declaration6631 specparam_declaration_instance6631();
    specparam_declaration6632 specparam_declaration_instance6632();
    specparam_declaration6633 specparam_declaration_instance6633();
    specparam_declaration6634 specparam_declaration_instance6634();
    specparam_declaration6635 specparam_declaration_instance6635();
    specparam_declaration6636 specparam_declaration_instance6636();
    specparam_declaration6637 specparam_declaration_instance6637();
    specparam_declaration6638 specparam_declaration_instance6638();
    specparam_declaration6639 specparam_declaration_instance6639();
    specparam_declaration6640 specparam_declaration_instance6640();
    specparam_declaration6641 specparam_declaration_instance6641();
    specparam_declaration6642 specparam_declaration_instance6642();
    specparam_declaration6643 specparam_declaration_instance6643();
    specparam_declaration6644 specparam_declaration_instance6644();
    specparam_declaration6645 specparam_declaration_instance6645();
    specparam_declaration6646 specparam_declaration_instance6646();
    specparam_declaration6647 specparam_declaration_instance6647();
    specparam_declaration6648 specparam_declaration_instance6648();
    specparam_declaration6649 specparam_declaration_instance6649();
    specparam_declaration6650 specparam_declaration_instance6650();
    specparam_declaration6651 specparam_declaration_instance6651();
    specparam_declaration6652 specparam_declaration_instance6652();
    specparam_declaration6653 specparam_declaration_instance6653();
    specparam_declaration6654 specparam_declaration_instance6654();
    specparam_declaration6655 specparam_declaration_instance6655();
    specparam_declaration6656 specparam_declaration_instance6656();
    specparam_declaration6657 specparam_declaration_instance6657();
    specparam_declaration6658 specparam_declaration_instance6658();
    specparam_declaration6659 specparam_declaration_instance6659();
    specparam_declaration6660 specparam_declaration_instance6660();
    specparam_declaration6661 specparam_declaration_instance6661();
    specparam_declaration6662 specparam_declaration_instance6662();
    specparam_declaration6663 specparam_declaration_instance6663();
    specparam_declaration6664 specparam_declaration_instance6664();
    specparam_declaration6665 specparam_declaration_instance6665();
    specparam_declaration6666 specparam_declaration_instance6666();
    specparam_declaration6667 specparam_declaration_instance6667();
    specparam_declaration6668 specparam_declaration_instance6668();
    specparam_declaration6669 specparam_declaration_instance6669();
    specparam_declaration6670 specparam_declaration_instance6670();
    specparam_declaration6671 specparam_declaration_instance6671();
    specparam_declaration6672 specparam_declaration_instance6672();
    specparam_declaration6673 specparam_declaration_instance6673();
    specparam_declaration6674 specparam_declaration_instance6674();
    specparam_declaration6675 specparam_declaration_instance6675();
    specparam_declaration6676 specparam_declaration_instance6676();
    specparam_declaration6677 specparam_declaration_instance6677();
    specparam_declaration6678 specparam_declaration_instance6678();
    specparam_declaration6679 specparam_declaration_instance6679();
    specparam_declaration6680 specparam_declaration_instance6680();
    specparam_declaration6681 specparam_declaration_instance6681();
    specparam_declaration6682 specparam_declaration_instance6682();
    specparam_declaration6683 specparam_declaration_instance6683();
    specparam_declaration6684 specparam_declaration_instance6684();
    specparam_declaration6685 specparam_declaration_instance6685();
    specparam_declaration6686 specparam_declaration_instance6686();
    specparam_declaration6687 specparam_declaration_instance6687();
    specparam_declaration6688 specparam_declaration_instance6688();
    specparam_declaration6689 specparam_declaration_instance6689();
    specparam_declaration6690 specparam_declaration_instance6690();
    specparam_declaration6691 specparam_declaration_instance6691();
    specparam_declaration6692 specparam_declaration_instance6692();
    specparam_declaration6693 specparam_declaration_instance6693();
    specparam_declaration6694 specparam_declaration_instance6694();
    specparam_declaration6695 specparam_declaration_instance6695();
    specparam_declaration6696 specparam_declaration_instance6696();
    specparam_declaration6697 specparam_declaration_instance6697();
    specparam_declaration6698 specparam_declaration_instance6698();
    specparam_declaration6699 specparam_declaration_instance6699();
    specparam_declaration6700 specparam_declaration_instance6700();
    specparam_declaration6701 specparam_declaration_instance6701();
    specparam_declaration6702 specparam_declaration_instance6702();
    specparam_declaration6703 specparam_declaration_instance6703();
    specparam_declaration6704 specparam_declaration_instance6704();
    specparam_declaration6705 specparam_declaration_instance6705();
    specparam_declaration6706 specparam_declaration_instance6706();
    specparam_declaration6707 specparam_declaration_instance6707();
    specparam_declaration6708 specparam_declaration_instance6708();
    specparam_declaration6709 specparam_declaration_instance6709();
    specparam_declaration6710 specparam_declaration_instance6710();
    specparam_declaration6711 specparam_declaration_instance6711();
    specparam_declaration6712 specparam_declaration_instance6712();
    specparam_declaration6713 specparam_declaration_instance6713();
    specparam_declaration6714 specparam_declaration_instance6714();
    specparam_declaration6715 specparam_declaration_instance6715();
    specparam_declaration6716 specparam_declaration_instance6716();
    specparam_declaration6717 specparam_declaration_instance6717();
    specparam_declaration6718 specparam_declaration_instance6718();
    specparam_declaration6719 specparam_declaration_instance6719();
    specparam_declaration6720 specparam_declaration_instance6720();
    specparam_declaration6721 specparam_declaration_instance6721();
    specparam_declaration6722 specparam_declaration_instance6722();
    specparam_declaration6723 specparam_declaration_instance6723();
    specparam_declaration6724 specparam_declaration_instance6724();
    specparam_declaration6725 specparam_declaration_instance6725();
    specparam_declaration6726 specparam_declaration_instance6726();
    specparam_declaration6727 specparam_declaration_instance6727();
    specparam_declaration6728 specparam_declaration_instance6728();
    specparam_declaration6729 specparam_declaration_instance6729();
    specparam_declaration6730 specparam_declaration_instance6730();
    specparam_declaration6731 specparam_declaration_instance6731();
    specparam_declaration6732 specparam_declaration_instance6732();
    specparam_declaration6733 specparam_declaration_instance6733();
    specparam_declaration6734 specparam_declaration_instance6734();
    specparam_declaration6735 specparam_declaration_instance6735();
    specparam_declaration6736 specparam_declaration_instance6736();
    specparam_declaration6737 specparam_declaration_instance6737();
    specparam_declaration6738 specparam_declaration_instance6738();
    specparam_declaration6739 specparam_declaration_instance6739();
    specparam_declaration6740 specparam_declaration_instance6740();
    specparam_declaration6741 specparam_declaration_instance6741();
    specparam_declaration6742 specparam_declaration_instance6742();
    specparam_declaration6743 specparam_declaration_instance6743();
    specparam_declaration6744 specparam_declaration_instance6744();
    specparam_declaration6745 specparam_declaration_instance6745();
    specparam_declaration6746 specparam_declaration_instance6746();
    specparam_declaration6747 specparam_declaration_instance6747();
    specparam_declaration6748 specparam_declaration_instance6748();
    specparam_declaration6749 specparam_declaration_instance6749();
    specparam_declaration6750 specparam_declaration_instance6750();
    specparam_declaration6751 specparam_declaration_instance6751();
    specparam_declaration6752 specparam_declaration_instance6752();
    specparam_declaration6753 specparam_declaration_instance6753();
    specparam_declaration6754 specparam_declaration_instance6754();
    specparam_declaration6755 specparam_declaration_instance6755();
    specparam_declaration6756 specparam_declaration_instance6756();
    specparam_declaration6757 specparam_declaration_instance6757();
    specparam_declaration6758 specparam_declaration_instance6758();
    specparam_declaration6759 specparam_declaration_instance6759();
    specparam_declaration6760 specparam_declaration_instance6760();
    specparam_declaration6761 specparam_declaration_instance6761();
    specparam_declaration6762 specparam_declaration_instance6762();
    specparam_declaration6763 specparam_declaration_instance6763();
    specparam_declaration6764 specparam_declaration_instance6764();
    specparam_declaration6765 specparam_declaration_instance6765();
    specparam_declaration6766 specparam_declaration_instance6766();
    specparam_declaration6767 specparam_declaration_instance6767();
    specparam_declaration6768 specparam_declaration_instance6768();
    specparam_declaration6769 specparam_declaration_instance6769();
    specparam_declaration6770 specparam_declaration_instance6770();
    specparam_declaration6771 specparam_declaration_instance6771();
    specparam_declaration6772 specparam_declaration_instance6772();
    specparam_declaration6773 specparam_declaration_instance6773();
    specparam_declaration6774 specparam_declaration_instance6774();
    specparam_declaration6775 specparam_declaration_instance6775();
    specparam_declaration6776 specparam_declaration_instance6776();
    specparam_declaration6777 specparam_declaration_instance6777();
    specparam_declaration6778 specparam_declaration_instance6778();
    specparam_declaration6779 specparam_declaration_instance6779();
    specparam_declaration6780 specparam_declaration_instance6780();
    specparam_declaration6781 specparam_declaration_instance6781();
    specparam_declaration6782 specparam_declaration_instance6782();
    specparam_declaration6783 specparam_declaration_instance6783();
    specparam_declaration6784 specparam_declaration_instance6784();
    specparam_declaration6785 specparam_declaration_instance6785();
    specparam_declaration6786 specparam_declaration_instance6786();
    specparam_declaration6787 specparam_declaration_instance6787();
    specparam_declaration6788 specparam_declaration_instance6788();
    specparam_declaration6789 specparam_declaration_instance6789();
    specparam_declaration6790 specparam_declaration_instance6790();
    specparam_declaration6791 specparam_declaration_instance6791();
    specparam_declaration6792 specparam_declaration_instance6792();
    specparam_declaration6793 specparam_declaration_instance6793();
    specparam_declaration6794 specparam_declaration_instance6794();
    specparam_declaration6795 specparam_declaration_instance6795();
    specparam_declaration6796 specparam_declaration_instance6796();
    specparam_declaration6797 specparam_declaration_instance6797();
    specparam_declaration6798 specparam_declaration_instance6798();
    specparam_declaration6799 specparam_declaration_instance6799();
    specparam_declaration6800 specparam_declaration_instance6800();
    specparam_declaration6801 specparam_declaration_instance6801();
    specparam_declaration6802 specparam_declaration_instance6802();
    specparam_declaration6803 specparam_declaration_instance6803();
    specparam_declaration6804 specparam_declaration_instance6804();
    specparam_declaration6805 specparam_declaration_instance6805();
    specparam_declaration6806 specparam_declaration_instance6806();
    specparam_declaration6807 specparam_declaration_instance6807();
    specparam_declaration6808 specparam_declaration_instance6808();
    specparam_declaration6809 specparam_declaration_instance6809();
    specparam_declaration6810 specparam_declaration_instance6810();
    specparam_declaration6811 specparam_declaration_instance6811();
    specparam_declaration6812 specparam_declaration_instance6812();
    specparam_declaration6813 specparam_declaration_instance6813();
    specparam_declaration6814 specparam_declaration_instance6814();
    specparam_declaration6815 specparam_declaration_instance6815();
    specparam_declaration6816 specparam_declaration_instance6816();
    specparam_declaration6817 specparam_declaration_instance6817();
    specparam_declaration6818 specparam_declaration_instance6818();
    specparam_declaration6819 specparam_declaration_instance6819();
    specparam_declaration6820 specparam_declaration_instance6820();
    specparam_declaration6821 specparam_declaration_instance6821();
    specparam_declaration6822 specparam_declaration_instance6822();
    specparam_declaration6823 specparam_declaration_instance6823();
    specparam_declaration6824 specparam_declaration_instance6824();
    specparam_declaration6825 specparam_declaration_instance6825();
    specparam_declaration6826 specparam_declaration_instance6826();
    specparam_declaration6827 specparam_declaration_instance6827();
    specparam_declaration6828 specparam_declaration_instance6828();
    specparam_declaration6829 specparam_declaration_instance6829();
    specparam_declaration6830 specparam_declaration_instance6830();
    specparam_declaration6831 specparam_declaration_instance6831();
    specparam_declaration6832 specparam_declaration_instance6832();
    specparam_declaration6833 specparam_declaration_instance6833();
    specparam_declaration6834 specparam_declaration_instance6834();
    specparam_declaration6835 specparam_declaration_instance6835();
    specparam_declaration6836 specparam_declaration_instance6836();
    specparam_declaration6837 specparam_declaration_instance6837();
    specparam_declaration6838 specparam_declaration_instance6838();
    specparam_declaration6839 specparam_declaration_instance6839();
    specparam_declaration6840 specparam_declaration_instance6840();
    specparam_declaration6841 specparam_declaration_instance6841();
    specparam_declaration6842 specparam_declaration_instance6842();
    specparam_declaration6843 specparam_declaration_instance6843();
    specparam_declaration6844 specparam_declaration_instance6844();
    specparam_declaration6845 specparam_declaration_instance6845();
    specparam_declaration6846 specparam_declaration_instance6846();
    specparam_declaration6847 specparam_declaration_instance6847();
    specparam_declaration6848 specparam_declaration_instance6848();
    specparam_declaration6849 specparam_declaration_instance6849();
    specparam_declaration6850 specparam_declaration_instance6850();
    specparam_declaration6851 specparam_declaration_instance6851();
    specparam_declaration6852 specparam_declaration_instance6852();
    specparam_declaration6853 specparam_declaration_instance6853();
    specparam_declaration6854 specparam_declaration_instance6854();
    specparam_declaration6855 specparam_declaration_instance6855();
    specparam_declaration6856 specparam_declaration_instance6856();
    specparam_declaration6857 specparam_declaration_instance6857();
    specparam_declaration6858 specparam_declaration_instance6858();
    specparam_declaration6859 specparam_declaration_instance6859();
    specparam_declaration6860 specparam_declaration_instance6860();
    specparam_declaration6861 specparam_declaration_instance6861();
    specparam_declaration6862 specparam_declaration_instance6862();
    specparam_declaration6863 specparam_declaration_instance6863();
    specparam_declaration6864 specparam_declaration_instance6864();
    specparam_declaration6865 specparam_declaration_instance6865();
    specparam_declaration6866 specparam_declaration_instance6866();
    specparam_declaration6867 specparam_declaration_instance6867();
    specparam_declaration6868 specparam_declaration_instance6868();
    specparam_declaration6869 specparam_declaration_instance6869();
    specparam_declaration6870 specparam_declaration_instance6870();
    specparam_declaration6871 specparam_declaration_instance6871();
    specparam_declaration6872 specparam_declaration_instance6872();
    specparam_declaration6873 specparam_declaration_instance6873();
    specparam_declaration6874 specparam_declaration_instance6874();
    specparam_declaration6875 specparam_declaration_instance6875();
    specparam_declaration6876 specparam_declaration_instance6876();
    specparam_declaration6877 specparam_declaration_instance6877();
    specparam_declaration6878 specparam_declaration_instance6878();
    specparam_declaration6879 specparam_declaration_instance6879();
    specparam_declaration6880 specparam_declaration_instance6880();
    specparam_declaration6881 specparam_declaration_instance6881();
    specparam_declaration6882 specparam_declaration_instance6882();
    specparam_declaration6883 specparam_declaration_instance6883();
    specparam_declaration6884 specparam_declaration_instance6884();
    specparam_declaration6885 specparam_declaration_instance6885();
    specparam_declaration6886 specparam_declaration_instance6886();
    specparam_declaration6887 specparam_declaration_instance6887();
    specparam_declaration6888 specparam_declaration_instance6888();
    specparam_declaration6889 specparam_declaration_instance6889();
    specparam_declaration6890 specparam_declaration_instance6890();
    specparam_declaration6891 specparam_declaration_instance6891();
    specparam_declaration6892 specparam_declaration_instance6892();
    specparam_declaration6893 specparam_declaration_instance6893();
    specparam_declaration6894 specparam_declaration_instance6894();
    specparam_declaration6895 specparam_declaration_instance6895();
    specparam_declaration6896 specparam_declaration_instance6896();
    specparam_declaration6897 specparam_declaration_instance6897();
    specparam_declaration6898 specparam_declaration_instance6898();
    specparam_declaration6899 specparam_declaration_instance6899();
    specparam_declaration6900 specparam_declaration_instance6900();
    specparam_declaration6901 specparam_declaration_instance6901();
    specparam_declaration6902 specparam_declaration_instance6902();
    specparam_declaration6903 specparam_declaration_instance6903();
    specparam_declaration6904 specparam_declaration_instance6904();
    specparam_declaration6905 specparam_declaration_instance6905();
    specparam_declaration6906 specparam_declaration_instance6906();
    specparam_declaration6907 specparam_declaration_instance6907();
    specparam_declaration6908 specparam_declaration_instance6908();
    specparam_declaration6909 specparam_declaration_instance6909();
    specparam_declaration6910 specparam_declaration_instance6910();
    specparam_declaration6911 specparam_declaration_instance6911();
    specparam_declaration6912 specparam_declaration_instance6912();
    specparam_declaration6913 specparam_declaration_instance6913();
    specparam_declaration6914 specparam_declaration_instance6914();
    specparam_declaration6915 specparam_declaration_instance6915();
    specparam_declaration6916 specparam_declaration_instance6916();
    specparam_declaration6917 specparam_declaration_instance6917();
    specparam_declaration6918 specparam_declaration_instance6918();
    specparam_declaration6919 specparam_declaration_instance6919();
    specparam_declaration6920 specparam_declaration_instance6920();
    specparam_declaration6921 specparam_declaration_instance6921();
    specparam_declaration6922 specparam_declaration_instance6922();
    specparam_declaration6923 specparam_declaration_instance6923();
    specparam_declaration6924 specparam_declaration_instance6924();
    specparam_declaration6925 specparam_declaration_instance6925();
    specparam_declaration6926 specparam_declaration_instance6926();
    specparam_declaration6927 specparam_declaration_instance6927();
    specparam_declaration6928 specparam_declaration_instance6928();
    specparam_declaration6929 specparam_declaration_instance6929();
    specparam_declaration6930 specparam_declaration_instance6930();
    specparam_declaration6931 specparam_declaration_instance6931();
    specparam_declaration6932 specparam_declaration_instance6932();
    specparam_declaration6933 specparam_declaration_instance6933();
    specparam_declaration6934 specparam_declaration_instance6934();
    specparam_declaration6935 specparam_declaration_instance6935();
    specparam_declaration6936 specparam_declaration_instance6936();
    specparam_declaration6937 specparam_declaration_instance6937();
    specparam_declaration6938 specparam_declaration_instance6938();
    specparam_declaration6939 specparam_declaration_instance6939();
    specparam_declaration6940 specparam_declaration_instance6940();
    specparam_declaration6941 specparam_declaration_instance6941();
    specparam_declaration6942 specparam_declaration_instance6942();
    specparam_declaration6943 specparam_declaration_instance6943();
    specparam_declaration6944 specparam_declaration_instance6944();
    specparam_declaration6945 specparam_declaration_instance6945();
    specparam_declaration6946 specparam_declaration_instance6946();
    specparam_declaration6947 specparam_declaration_instance6947();
    specparam_declaration6948 specparam_declaration_instance6948();
    specparam_declaration6949 specparam_declaration_instance6949();
    specparam_declaration6950 specparam_declaration_instance6950();
    specparam_declaration6951 specparam_declaration_instance6951();
    specparam_declaration6952 specparam_declaration_instance6952();
    specparam_declaration6953 specparam_declaration_instance6953();
    specparam_declaration6954 specparam_declaration_instance6954();
    specparam_declaration6955 specparam_declaration_instance6955();
    specparam_declaration6956 specparam_declaration_instance6956();
    specparam_declaration6957 specparam_declaration_instance6957();
    specparam_declaration6958 specparam_declaration_instance6958();
    specparam_declaration6959 specparam_declaration_instance6959();
    specparam_declaration6960 specparam_declaration_instance6960();
    specparam_declaration6961 specparam_declaration_instance6961();
    specparam_declaration6962 specparam_declaration_instance6962();
    specparam_declaration6963 specparam_declaration_instance6963();
    specparam_declaration6964 specparam_declaration_instance6964();
    specparam_declaration6965 specparam_declaration_instance6965();
    specparam_declaration6966 specparam_declaration_instance6966();
    specparam_declaration6967 specparam_declaration_instance6967();
    specparam_declaration6968 specparam_declaration_instance6968();
    specparam_declaration6969 specparam_declaration_instance6969();
    specparam_declaration6970 specparam_declaration_instance6970();
    specparam_declaration6971 specparam_declaration_instance6971();
    specparam_declaration6972 specparam_declaration_instance6972();
    specparam_declaration6973 specparam_declaration_instance6973();
    specparam_declaration6974 specparam_declaration_instance6974();
    specparam_declaration6975 specparam_declaration_instance6975();
    specparam_declaration6976 specparam_declaration_instance6976();
    specparam_declaration6977 specparam_declaration_instance6977();
    specparam_declaration6978 specparam_declaration_instance6978();
    specparam_declaration6979 specparam_declaration_instance6979();
    specparam_declaration6980 specparam_declaration_instance6980();
    specparam_declaration6981 specparam_declaration_instance6981();
    specparam_declaration6982 specparam_declaration_instance6982();
    specparam_declaration6983 specparam_declaration_instance6983();
    specparam_declaration6984 specparam_declaration_instance6984();
    specparam_declaration6985 specparam_declaration_instance6985();
    specparam_declaration6986 specparam_declaration_instance6986();
    specparam_declaration6987 specparam_declaration_instance6987();
    specparam_declaration6988 specparam_declaration_instance6988();
    specparam_declaration6989 specparam_declaration_instance6989();
    specparam_declaration6990 specparam_declaration_instance6990();
    specparam_declaration6991 specparam_declaration_instance6991();
    specparam_declaration6992 specparam_declaration_instance6992();
    specparam_declaration6993 specparam_declaration_instance6993();
    specparam_declaration6994 specparam_declaration_instance6994();
    specparam_declaration6995 specparam_declaration_instance6995();
    specparam_declaration6996 specparam_declaration_instance6996();
    specparam_declaration6997 specparam_declaration_instance6997();
    specparam_declaration6998 specparam_declaration_instance6998();
    specparam_declaration6999 specparam_declaration_instance6999();
    specparam_declaration7000 specparam_declaration_instance7000();
    specparam_declaration7001 specparam_declaration_instance7001();
    specparam_declaration7002 specparam_declaration_instance7002();
    specparam_declaration7003 specparam_declaration_instance7003();
    specparam_declaration7004 specparam_declaration_instance7004();
    specparam_declaration7005 specparam_declaration_instance7005();
    specparam_declaration7006 specparam_declaration_instance7006();
    specparam_declaration7007 specparam_declaration_instance7007();
    specparam_declaration7008 specparam_declaration_instance7008();
    specparam_declaration7009 specparam_declaration_instance7009();
    specparam_declaration7010 specparam_declaration_instance7010();
    specparam_declaration7011 specparam_declaration_instance7011();
    specparam_declaration7012 specparam_declaration_instance7012();
    specparam_declaration7013 specparam_declaration_instance7013();
    specparam_declaration7014 specparam_declaration_instance7014();
    specparam_declaration7015 specparam_declaration_instance7015();
    specparam_declaration7016 specparam_declaration_instance7016();
    specparam_declaration7017 specparam_declaration_instance7017();
    specparam_declaration7018 specparam_declaration_instance7018();
    specparam_declaration7019 specparam_declaration_instance7019();
    specparam_declaration7020 specparam_declaration_instance7020();
    specparam_declaration7021 specparam_declaration_instance7021();
    specparam_declaration7022 specparam_declaration_instance7022();
    specparam_declaration7023 specparam_declaration_instance7023();
    specparam_declaration7024 specparam_declaration_instance7024();
    specparam_declaration7025 specparam_declaration_instance7025();
    specparam_declaration7026 specparam_declaration_instance7026();
    specparam_declaration7027 specparam_declaration_instance7027();
    specparam_declaration7028 specparam_declaration_instance7028();
    specparam_declaration7029 specparam_declaration_instance7029();
    specparam_declaration7030 specparam_declaration_instance7030();
    specparam_declaration7031 specparam_declaration_instance7031();
    specparam_declaration7032 specparam_declaration_instance7032();
    specparam_declaration7033 specparam_declaration_instance7033();
    specparam_declaration7034 specparam_declaration_instance7034();
    specparam_declaration7035 specparam_declaration_instance7035();
    specparam_declaration7036 specparam_declaration_instance7036();
    specparam_declaration7037 specparam_declaration_instance7037();
    specparam_declaration7038 specparam_declaration_instance7038();
    specparam_declaration7039 specparam_declaration_instance7039();
    specparam_declaration7040 specparam_declaration_instance7040();
    specparam_declaration7041 specparam_declaration_instance7041();
    specparam_declaration7042 specparam_declaration_instance7042();
    specparam_declaration7043 specparam_declaration_instance7043();
    specparam_declaration7044 specparam_declaration_instance7044();
    specparam_declaration7045 specparam_declaration_instance7045();
    specparam_declaration7046 specparam_declaration_instance7046();
    specparam_declaration7047 specparam_declaration_instance7047();
    specparam_declaration7048 specparam_declaration_instance7048();
    specparam_declaration7049 specparam_declaration_instance7049();
    specparam_declaration7050 specparam_declaration_instance7050();
    specparam_declaration7051 specparam_declaration_instance7051();
    specparam_declaration7052 specparam_declaration_instance7052();
    specparam_declaration7053 specparam_declaration_instance7053();
    specparam_declaration7054 specparam_declaration_instance7054();
    specparam_declaration7055 specparam_declaration_instance7055();
    specparam_declaration7056 specparam_declaration_instance7056();
    specparam_declaration7057 specparam_declaration_instance7057();
    specparam_declaration7058 specparam_declaration_instance7058();
    specparam_declaration7059 specparam_declaration_instance7059();
    specparam_declaration7060 specparam_declaration_instance7060();
    specparam_declaration7061 specparam_declaration_instance7061();
    specparam_declaration7062 specparam_declaration_instance7062();
    specparam_declaration7063 specparam_declaration_instance7063();
    specparam_declaration7064 specparam_declaration_instance7064();
    specparam_declaration7065 specparam_declaration_instance7065();
    specparam_declaration7066 specparam_declaration_instance7066();
    specparam_declaration7067 specparam_declaration_instance7067();
    specparam_declaration7068 specparam_declaration_instance7068();
    specparam_declaration7069 specparam_declaration_instance7069();
    specparam_declaration7070 specparam_declaration_instance7070();
    specparam_declaration7071 specparam_declaration_instance7071();
    specparam_declaration7072 specparam_declaration_instance7072();
    specparam_declaration7073 specparam_declaration_instance7073();
    specparam_declaration7074 specparam_declaration_instance7074();
    specparam_declaration7075 specparam_declaration_instance7075();
    specparam_declaration7076 specparam_declaration_instance7076();
    specparam_declaration7077 specparam_declaration_instance7077();
    specparam_declaration7078 specparam_declaration_instance7078();
    specparam_declaration7079 specparam_declaration_instance7079();
    specparam_declaration7080 specparam_declaration_instance7080();
    specparam_declaration7081 specparam_declaration_instance7081();
    specparam_declaration7082 specparam_declaration_instance7082();
    specparam_declaration7083 specparam_declaration_instance7083();
    specparam_declaration7084 specparam_declaration_instance7084();
    specparam_declaration7085 specparam_declaration_instance7085();
    specparam_declaration7086 specparam_declaration_instance7086();
    specparam_declaration7087 specparam_declaration_instance7087();
    specparam_declaration7088 specparam_declaration_instance7088();
    specparam_declaration7089 specparam_declaration_instance7089();
    specparam_declaration7090 specparam_declaration_instance7090();
    specparam_declaration7091 specparam_declaration_instance7091();
    specparam_declaration7092 specparam_declaration_instance7092();
    specparam_declaration7093 specparam_declaration_instance7093();
    specparam_declaration7094 specparam_declaration_instance7094();
    specparam_declaration7095 specparam_declaration_instance7095();
    specparam_declaration7096 specparam_declaration_instance7096();
    specparam_declaration7097 specparam_declaration_instance7097();
    specparam_declaration7098 specparam_declaration_instance7098();
    specparam_declaration7099 specparam_declaration_instance7099();
    specparam_declaration7100 specparam_declaration_instance7100();
    specparam_declaration7101 specparam_declaration_instance7101();
    specparam_declaration7102 specparam_declaration_instance7102();
    specparam_declaration7103 specparam_declaration_instance7103();
    specparam_declaration7104 specparam_declaration_instance7104();
    specparam_declaration7105 specparam_declaration_instance7105();
    specparam_declaration7106 specparam_declaration_instance7106();
    specparam_declaration7107 specparam_declaration_instance7107();
    specparam_declaration7108 specparam_declaration_instance7108();
    specparam_declaration7109 specparam_declaration_instance7109();
    specparam_declaration7110 specparam_declaration_instance7110();
    specparam_declaration7111 specparam_declaration_instance7111();
    specparam_declaration7112 specparam_declaration_instance7112();
    specparam_declaration7113 specparam_declaration_instance7113();
    specparam_declaration7114 specparam_declaration_instance7114();
    specparam_declaration7115 specparam_declaration_instance7115();
    specparam_declaration7116 specparam_declaration_instance7116();
    specparam_declaration7117 specparam_declaration_instance7117();
    specparam_declaration7118 specparam_declaration_instance7118();
    specparam_declaration7119 specparam_declaration_instance7119();
    specparam_declaration7120 specparam_declaration_instance7120();
    specparam_declaration7121 specparam_declaration_instance7121();
    specparam_declaration7122 specparam_declaration_instance7122();
    specparam_declaration7123 specparam_declaration_instance7123();
    specparam_declaration7124 specparam_declaration_instance7124();
    specparam_declaration7125 specparam_declaration_instance7125();
    specparam_declaration7126 specparam_declaration_instance7126();
    specparam_declaration7127 specparam_declaration_instance7127();
    specparam_declaration7128 specparam_declaration_instance7128();
    specparam_declaration7129 specparam_declaration_instance7129();
    specparam_declaration7130 specparam_declaration_instance7130();
    specparam_declaration7131 specparam_declaration_instance7131();
    specparam_declaration7132 specparam_declaration_instance7132();
    specparam_declaration7133 specparam_declaration_instance7133();
    specparam_declaration7134 specparam_declaration_instance7134();
    specparam_declaration7135 specparam_declaration_instance7135();
    specparam_declaration7136 specparam_declaration_instance7136();
    specparam_declaration7137 specparam_declaration_instance7137();
    specparam_declaration7138 specparam_declaration_instance7138();
    specparam_declaration7139 specparam_declaration_instance7139();
    specparam_declaration7140 specparam_declaration_instance7140();
    specparam_declaration7141 specparam_declaration_instance7141();
    specparam_declaration7142 specparam_declaration_instance7142();
    specparam_declaration7143 specparam_declaration_instance7143();
    specparam_declaration7144 specparam_declaration_instance7144();
    specparam_declaration7145 specparam_declaration_instance7145();
    specparam_declaration7146 specparam_declaration_instance7146();
    specparam_declaration7147 specparam_declaration_instance7147();
    specparam_declaration7148 specparam_declaration_instance7148();
    specparam_declaration7149 specparam_declaration_instance7149();
    specparam_declaration7150 specparam_declaration_instance7150();
    specparam_declaration7151 specparam_declaration_instance7151();
    specparam_declaration7152 specparam_declaration_instance7152();
    specparam_declaration7153 specparam_declaration_instance7153();
    specparam_declaration7154 specparam_declaration_instance7154();
    specparam_declaration7155 specparam_declaration_instance7155();
    specparam_declaration7156 specparam_declaration_instance7156();
    specparam_declaration7157 specparam_declaration_instance7157();
    specparam_declaration7158 specparam_declaration_instance7158();
    specparam_declaration7159 specparam_declaration_instance7159();
    specparam_declaration7160 specparam_declaration_instance7160();
    specparam_declaration7161 specparam_declaration_instance7161();
    specparam_declaration7162 specparam_declaration_instance7162();
    specparam_declaration7163 specparam_declaration_instance7163();
    specparam_declaration7164 specparam_declaration_instance7164();
    specparam_declaration7165 specparam_declaration_instance7165();
    specparam_declaration7166 specparam_declaration_instance7166();
    specparam_declaration7167 specparam_declaration_instance7167();
    specparam_declaration7168 specparam_declaration_instance7168();
    specparam_declaration7169 specparam_declaration_instance7169();
    specparam_declaration7170 specparam_declaration_instance7170();
    specparam_declaration7171 specparam_declaration_instance7171();
    specparam_declaration7172 specparam_declaration_instance7172();
    specparam_declaration7173 specparam_declaration_instance7173();
    specparam_declaration7174 specparam_declaration_instance7174();
    specparam_declaration7175 specparam_declaration_instance7175();
    specparam_declaration7176 specparam_declaration_instance7176();
    specparam_declaration7177 specparam_declaration_instance7177();
    specparam_declaration7178 specparam_declaration_instance7178();
    specparam_declaration7179 specparam_declaration_instance7179();
    specparam_declaration7180 specparam_declaration_instance7180();
    specparam_declaration7181 specparam_declaration_instance7181();
    specparam_declaration7182 specparam_declaration_instance7182();
    specparam_declaration7183 specparam_declaration_instance7183();
    specparam_declaration7184 specparam_declaration_instance7184();
    specparam_declaration7185 specparam_declaration_instance7185();
    specparam_declaration7186 specparam_declaration_instance7186();
    specparam_declaration7187 specparam_declaration_instance7187();
    specparam_declaration7188 specparam_declaration_instance7188();
    specparam_declaration7189 specparam_declaration_instance7189();
    specparam_declaration7190 specparam_declaration_instance7190();
    specparam_declaration7191 specparam_declaration_instance7191();
    specparam_declaration7192 specparam_declaration_instance7192();
    specparam_declaration7193 specparam_declaration_instance7193();
    specparam_declaration7194 specparam_declaration_instance7194();
    specparam_declaration7195 specparam_declaration_instance7195();
    specparam_declaration7196 specparam_declaration_instance7196();
    specparam_declaration7197 specparam_declaration_instance7197();
    specparam_declaration7198 specparam_declaration_instance7198();
    specparam_declaration7199 specparam_declaration_instance7199();
    specparam_declaration7200 specparam_declaration_instance7200();
    specparam_declaration7201 specparam_declaration_instance7201();
    specparam_declaration7202 specparam_declaration_instance7202();
    specparam_declaration7203 specparam_declaration_instance7203();
    specparam_declaration7204 specparam_declaration_instance7204();
    specparam_declaration7205 specparam_declaration_instance7205();
    specparam_declaration7206 specparam_declaration_instance7206();
    specparam_declaration7207 specparam_declaration_instance7207();
    specparam_declaration7208 specparam_declaration_instance7208();
    specparam_declaration7209 specparam_declaration_instance7209();
    specparam_declaration7210 specparam_declaration_instance7210();
    specparam_declaration7211 specparam_declaration_instance7211();
    specparam_declaration7212 specparam_declaration_instance7212();
    specparam_declaration7213 specparam_declaration_instance7213();
    specparam_declaration7214 specparam_declaration_instance7214();
    specparam_declaration7215 specparam_declaration_instance7215();
    specparam_declaration7216 specparam_declaration_instance7216();
    specparam_declaration7217 specparam_declaration_instance7217();
    specparam_declaration7218 specparam_declaration_instance7218();
    specparam_declaration7219 specparam_declaration_instance7219();
    specparam_declaration7220 specparam_declaration_instance7220();
    specparam_declaration7221 specparam_declaration_instance7221();
    specparam_declaration7222 specparam_declaration_instance7222();
    specparam_declaration7223 specparam_declaration_instance7223();
    specparam_declaration7224 specparam_declaration_instance7224();
    specparam_declaration7225 specparam_declaration_instance7225();
    specparam_declaration7226 specparam_declaration_instance7226();
    specparam_declaration7227 specparam_declaration_instance7227();
    specparam_declaration7228 specparam_declaration_instance7228();
    specparam_declaration7229 specparam_declaration_instance7229();
    specparam_declaration7230 specparam_declaration_instance7230();
    specparam_declaration7231 specparam_declaration_instance7231();
    specparam_declaration7232 specparam_declaration_instance7232();
    specparam_declaration7233 specparam_declaration_instance7233();
    specparam_declaration7234 specparam_declaration_instance7234();
    specparam_declaration7235 specparam_declaration_instance7235();
    specparam_declaration7236 specparam_declaration_instance7236();
    specparam_declaration7237 specparam_declaration_instance7237();
    specparam_declaration7238 specparam_declaration_instance7238();
    specparam_declaration7239 specparam_declaration_instance7239();
    specparam_declaration7240 specparam_declaration_instance7240();
    specparam_declaration7241 specparam_declaration_instance7241();
    specparam_declaration7242 specparam_declaration_instance7242();
    specparam_declaration7243 specparam_declaration_instance7243();
    specparam_declaration7244 specparam_declaration_instance7244();
    specparam_declaration7245 specparam_declaration_instance7245();
    specparam_declaration7246 specparam_declaration_instance7246();
    specparam_declaration7247 specparam_declaration_instance7247();
    specparam_declaration7248 specparam_declaration_instance7248();
    specparam_declaration7249 specparam_declaration_instance7249();
    specparam_declaration7250 specparam_declaration_instance7250();
    specparam_declaration7251 specparam_declaration_instance7251();
    specparam_declaration7252 specparam_declaration_instance7252();
    specparam_declaration7253 specparam_declaration_instance7253();
    specparam_declaration7254 specparam_declaration_instance7254();
    specparam_declaration7255 specparam_declaration_instance7255();
    specparam_declaration7256 specparam_declaration_instance7256();
    specparam_declaration7257 specparam_declaration_instance7257();
    specparam_declaration7258 specparam_declaration_instance7258();
    specparam_declaration7259 specparam_declaration_instance7259();
    specparam_declaration7260 specparam_declaration_instance7260();
    specparam_declaration7261 specparam_declaration_instance7261();
    specparam_declaration7262 specparam_declaration_instance7262();
    specparam_declaration7263 specparam_declaration_instance7263();
    specparam_declaration7264 specparam_declaration_instance7264();
    specparam_declaration7265 specparam_declaration_instance7265();
    specparam_declaration7266 specparam_declaration_instance7266();
    specparam_declaration7267 specparam_declaration_instance7267();
    specparam_declaration7268 specparam_declaration_instance7268();
    specparam_declaration7269 specparam_declaration_instance7269();
    specparam_declaration7270 specparam_declaration_instance7270();
    specparam_declaration7271 specparam_declaration_instance7271();
    specparam_declaration7272 specparam_declaration_instance7272();
    specparam_declaration7273 specparam_declaration_instance7273();
    specparam_declaration7274 specparam_declaration_instance7274();
    specparam_declaration7275 specparam_declaration_instance7275();
    specparam_declaration7276 specparam_declaration_instance7276();
    specparam_declaration7277 specparam_declaration_instance7277();
    specparam_declaration7278 specparam_declaration_instance7278();
    specparam_declaration7279 specparam_declaration_instance7279();
    specparam_declaration7280 specparam_declaration_instance7280();
    specparam_declaration7281 specparam_declaration_instance7281();
    specparam_declaration7282 specparam_declaration_instance7282();
    specparam_declaration7283 specparam_declaration_instance7283();
    specparam_declaration7284 specparam_declaration_instance7284();
    specparam_declaration7285 specparam_declaration_instance7285();
    specparam_declaration7286 specparam_declaration_instance7286();
    specparam_declaration7287 specparam_declaration_instance7287();
    specparam_declaration7288 specparam_declaration_instance7288();
    specparam_declaration7289 specparam_declaration_instance7289();
    specparam_declaration7290 specparam_declaration_instance7290();
    specparam_declaration7291 specparam_declaration_instance7291();
    specparam_declaration7292 specparam_declaration_instance7292();
    specparam_declaration7293 specparam_declaration_instance7293();
    specparam_declaration7294 specparam_declaration_instance7294();
    specparam_declaration7295 specparam_declaration_instance7295();
    specparam_declaration7296 specparam_declaration_instance7296();
    specparam_declaration7297 specparam_declaration_instance7297();
    specparam_declaration7298 specparam_declaration_instance7298();
    specparam_declaration7299 specparam_declaration_instance7299();
    specparam_declaration7300 specparam_declaration_instance7300();
    specparam_declaration7301 specparam_declaration_instance7301();
    specparam_declaration7302 specparam_declaration_instance7302();
    specparam_declaration7303 specparam_declaration_instance7303();
    specparam_declaration7304 specparam_declaration_instance7304();
    specparam_declaration7305 specparam_declaration_instance7305();
    specparam_declaration7306 specparam_declaration_instance7306();
    specparam_declaration7307 specparam_declaration_instance7307();
    specparam_declaration7308 specparam_declaration_instance7308();
    specparam_declaration7309 specparam_declaration_instance7309();
    specparam_declaration7310 specparam_declaration_instance7310();
    specparam_declaration7311 specparam_declaration_instance7311();
    specparam_declaration7312 specparam_declaration_instance7312();
    specparam_declaration7313 specparam_declaration_instance7313();
    specparam_declaration7314 specparam_declaration_instance7314();
    specparam_declaration7315 specparam_declaration_instance7315();
    specparam_declaration7316 specparam_declaration_instance7316();
    specparam_declaration7317 specparam_declaration_instance7317();
    specparam_declaration7318 specparam_declaration_instance7318();
    specparam_declaration7319 specparam_declaration_instance7319();
    specparam_declaration7320 specparam_declaration_instance7320();
    specparam_declaration7321 specparam_declaration_instance7321();
    specparam_declaration7322 specparam_declaration_instance7322();
    specparam_declaration7323 specparam_declaration_instance7323();
    specparam_declaration7324 specparam_declaration_instance7324();
    specparam_declaration7325 specparam_declaration_instance7325();
    specparam_declaration7326 specparam_declaration_instance7326();
    specparam_declaration7327 specparam_declaration_instance7327();
    specparam_declaration7328 specparam_declaration_instance7328();
    specparam_declaration7329 specparam_declaration_instance7329();
    specparam_declaration7330 specparam_declaration_instance7330();
    specparam_declaration7331 specparam_declaration_instance7331();
    specparam_declaration7332 specparam_declaration_instance7332();
    specparam_declaration7333 specparam_declaration_instance7333();
    specparam_declaration7334 specparam_declaration_instance7334();
    specparam_declaration7335 specparam_declaration_instance7335();
    specparam_declaration7336 specparam_declaration_instance7336();
    specparam_declaration7337 specparam_declaration_instance7337();
    specparam_declaration7338 specparam_declaration_instance7338();
    specparam_declaration7339 specparam_declaration_instance7339();
    specparam_declaration7340 specparam_declaration_instance7340();
    specparam_declaration7341 specparam_declaration_instance7341();
    specparam_declaration7342 specparam_declaration_instance7342();
    specparam_declaration7343 specparam_declaration_instance7343();
    specparam_declaration7344 specparam_declaration_instance7344();
    specparam_declaration7345 specparam_declaration_instance7345();
    specparam_declaration7346 specparam_declaration_instance7346();
    specparam_declaration7347 specparam_declaration_instance7347();
    specparam_declaration7348 specparam_declaration_instance7348();
    specparam_declaration7349 specparam_declaration_instance7349();
    specparam_declaration7350 specparam_declaration_instance7350();
    specparam_declaration7351 specparam_declaration_instance7351();
    specparam_declaration7352 specparam_declaration_instance7352();
    specparam_declaration7353 specparam_declaration_instance7353();
    specparam_declaration7354 specparam_declaration_instance7354();
    specparam_declaration7355 specparam_declaration_instance7355();
    specparam_declaration7356 specparam_declaration_instance7356();
    specparam_declaration7357 specparam_declaration_instance7357();
    specparam_declaration7358 specparam_declaration_instance7358();
    specparam_declaration7359 specparam_declaration_instance7359();
    specparam_declaration7360 specparam_declaration_instance7360();
    specparam_declaration7361 specparam_declaration_instance7361();
    specparam_declaration7362 specparam_declaration_instance7362();
    specparam_declaration7363 specparam_declaration_instance7363();
    specparam_declaration7364 specparam_declaration_instance7364();
    specparam_declaration7365 specparam_declaration_instance7365();
    specparam_declaration7366 specparam_declaration_instance7366();
    specparam_declaration7367 specparam_declaration_instance7367();
    specparam_declaration7368 specparam_declaration_instance7368();
    specparam_declaration7369 specparam_declaration_instance7369();
    specparam_declaration7370 specparam_declaration_instance7370();
    specparam_declaration7371 specparam_declaration_instance7371();
    specparam_declaration7372 specparam_declaration_instance7372();
    specparam_declaration7373 specparam_declaration_instance7373();
    specparam_declaration7374 specparam_declaration_instance7374();
    specparam_declaration7375 specparam_declaration_instance7375();
    specparam_declaration7376 specparam_declaration_instance7376();
    specparam_declaration7377 specparam_declaration_instance7377();
    specparam_declaration7378 specparam_declaration_instance7378();
    specparam_declaration7379 specparam_declaration_instance7379();
    specparam_declaration7380 specparam_declaration_instance7380();
    specparam_declaration7381 specparam_declaration_instance7381();
    specparam_declaration7382 specparam_declaration_instance7382();
    specparam_declaration7383 specparam_declaration_instance7383();
    specparam_declaration7384 specparam_declaration_instance7384();
    specparam_declaration7385 specparam_declaration_instance7385();
    specparam_declaration7386 specparam_declaration_instance7386();
    specparam_declaration7387 specparam_declaration_instance7387();
    specparam_declaration7388 specparam_declaration_instance7388();
    specparam_declaration7389 specparam_declaration_instance7389();
    specparam_declaration7390 specparam_declaration_instance7390();
    specparam_declaration7391 specparam_declaration_instance7391();
    specparam_declaration7392 specparam_declaration_instance7392();
    specparam_declaration7393 specparam_declaration_instance7393();
    specparam_declaration7394 specparam_declaration_instance7394();
    specparam_declaration7395 specparam_declaration_instance7395();
    specparam_declaration7396 specparam_declaration_instance7396();
    specparam_declaration7397 specparam_declaration_instance7397();
    specparam_declaration7398 specparam_declaration_instance7398();
    specparam_declaration7399 specparam_declaration_instance7399();
    specparam_declaration7400 specparam_declaration_instance7400();
    specparam_declaration7401 specparam_declaration_instance7401();
    specparam_declaration7402 specparam_declaration_instance7402();
    specparam_declaration7403 specparam_declaration_instance7403();
    specparam_declaration7404 specparam_declaration_instance7404();
    specparam_declaration7405 specparam_declaration_instance7405();
    specparam_declaration7406 specparam_declaration_instance7406();
    specparam_declaration7407 specparam_declaration_instance7407();
    specparam_declaration7408 specparam_declaration_instance7408();
    specparam_declaration7409 specparam_declaration_instance7409();
    specparam_declaration7410 specparam_declaration_instance7410();
    specparam_declaration7411 specparam_declaration_instance7411();
    specparam_declaration7412 specparam_declaration_instance7412();
    specparam_declaration7413 specparam_declaration_instance7413();
    specparam_declaration7414 specparam_declaration_instance7414();
    specparam_declaration7415 specparam_declaration_instance7415();
    specparam_declaration7416 specparam_declaration_instance7416();
    specparam_declaration7417 specparam_declaration_instance7417();
    specparam_declaration7418 specparam_declaration_instance7418();
    specparam_declaration7419 specparam_declaration_instance7419();
    specparam_declaration7420 specparam_declaration_instance7420();
    specparam_declaration7421 specparam_declaration_instance7421();
    specparam_declaration7422 specparam_declaration_instance7422();
    specparam_declaration7423 specparam_declaration_instance7423();
    specparam_declaration7424 specparam_declaration_instance7424();
    specparam_declaration7425 specparam_declaration_instance7425();
    specparam_declaration7426 specparam_declaration_instance7426();
    specparam_declaration7427 specparam_declaration_instance7427();
    specparam_declaration7428 specparam_declaration_instance7428();
    specparam_declaration7429 specparam_declaration_instance7429();
    specparam_declaration7430 specparam_declaration_instance7430();
    specparam_declaration7431 specparam_declaration_instance7431();
    specparam_declaration7432 specparam_declaration_instance7432();
    specparam_declaration7433 specparam_declaration_instance7433();
    specparam_declaration7434 specparam_declaration_instance7434();
    specparam_declaration7435 specparam_declaration_instance7435();
    specparam_declaration7436 specparam_declaration_instance7436();
    specparam_declaration7437 specparam_declaration_instance7437();
    specparam_declaration7438 specparam_declaration_instance7438();
    specparam_declaration7439 specparam_declaration_instance7439();
    specparam_declaration7440 specparam_declaration_instance7440();
    specparam_declaration7441 specparam_declaration_instance7441();
    specparam_declaration7442 specparam_declaration_instance7442();
    specparam_declaration7443 specparam_declaration_instance7443();
    specparam_declaration7444 specparam_declaration_instance7444();
    specparam_declaration7445 specparam_declaration_instance7445();
    specparam_declaration7446 specparam_declaration_instance7446();
    specparam_declaration7447 specparam_declaration_instance7447();
    specparam_declaration7448 specparam_declaration_instance7448();
    specparam_declaration7449 specparam_declaration_instance7449();
    specparam_declaration7450 specparam_declaration_instance7450();
    specparam_declaration7451 specparam_declaration_instance7451();
    specparam_declaration7452 specparam_declaration_instance7452();
    specparam_declaration7453 specparam_declaration_instance7453();
    specparam_declaration7454 specparam_declaration_instance7454();
    specparam_declaration7455 specparam_declaration_instance7455();
    specparam_declaration7456 specparam_declaration_instance7456();
    specparam_declaration7457 specparam_declaration_instance7457();
    specparam_declaration7458 specparam_declaration_instance7458();
    specparam_declaration7459 specparam_declaration_instance7459();
    specparam_declaration7460 specparam_declaration_instance7460();
    specparam_declaration7461 specparam_declaration_instance7461();
    specparam_declaration7462 specparam_declaration_instance7462();
    specparam_declaration7463 specparam_declaration_instance7463();
    specparam_declaration7464 specparam_declaration_instance7464();
    specparam_declaration7465 specparam_declaration_instance7465();
    specparam_declaration7466 specparam_declaration_instance7466();
    specparam_declaration7467 specparam_declaration_instance7467();
    specparam_declaration7468 specparam_declaration_instance7468();
    specparam_declaration7469 specparam_declaration_instance7469();
    specparam_declaration7470 specparam_declaration_instance7470();
    specparam_declaration7471 specparam_declaration_instance7471();
    specparam_declaration7472 specparam_declaration_instance7472();
    specparam_declaration7473 specparam_declaration_instance7473();
    specparam_declaration7474 specparam_declaration_instance7474();
    specparam_declaration7475 specparam_declaration_instance7475();
    specparam_declaration7476 specparam_declaration_instance7476();
    specparam_declaration7477 specparam_declaration_instance7477();
    specparam_declaration7478 specparam_declaration_instance7478();
    specparam_declaration7479 specparam_declaration_instance7479();
    specparam_declaration7480 specparam_declaration_instance7480();
    specparam_declaration7481 specparam_declaration_instance7481();
    specparam_declaration7482 specparam_declaration_instance7482();
    specparam_declaration7483 specparam_declaration_instance7483();
    specparam_declaration7484 specparam_declaration_instance7484();
    specparam_declaration7485 specparam_declaration_instance7485();
    specparam_declaration7486 specparam_declaration_instance7486();
    specparam_declaration7487 specparam_declaration_instance7487();
    specparam_declaration7488 specparam_declaration_instance7488();
    specparam_declaration7489 specparam_declaration_instance7489();
    specparam_declaration7490 specparam_declaration_instance7490();
    specparam_declaration7491 specparam_declaration_instance7491();
    specparam_declaration7492 specparam_declaration_instance7492();
    specparam_declaration7493 specparam_declaration_instance7493();
    specparam_declaration7494 specparam_declaration_instance7494();
    specparam_declaration7495 specparam_declaration_instance7495();
    specparam_declaration7496 specparam_declaration_instance7496();
    specparam_declaration7497 specparam_declaration_instance7497();
    specparam_declaration7498 specparam_declaration_instance7498();
    specparam_declaration7499 specparam_declaration_instance7499();
    specparam_declaration7500 specparam_declaration_instance7500();
    specparam_declaration7501 specparam_declaration_instance7501();
    specparam_declaration7502 specparam_declaration_instance7502();
    specparam_declaration7503 specparam_declaration_instance7503();
    specparam_declaration7504 specparam_declaration_instance7504();
    specparam_declaration7505 specparam_declaration_instance7505();
    specparam_declaration7506 specparam_declaration_instance7506();
    specparam_declaration7507 specparam_declaration_instance7507();
    specparam_declaration7508 specparam_declaration_instance7508();
    specparam_declaration7509 specparam_declaration_instance7509();
    specparam_declaration7510 specparam_declaration_instance7510();
    specparam_declaration7511 specparam_declaration_instance7511();
    specparam_declaration7512 specparam_declaration_instance7512();
    specparam_declaration7513 specparam_declaration_instance7513();
    specparam_declaration7514 specparam_declaration_instance7514();
    specparam_declaration7515 specparam_declaration_instance7515();
    specparam_declaration7516 specparam_declaration_instance7516();
    specparam_declaration7517 specparam_declaration_instance7517();
    specparam_declaration7518 specparam_declaration_instance7518();
    specparam_declaration7519 specparam_declaration_instance7519();
    specparam_declaration7520 specparam_declaration_instance7520();
    specparam_declaration7521 specparam_declaration_instance7521();
    specparam_declaration7522 specparam_declaration_instance7522();
    specparam_declaration7523 specparam_declaration_instance7523();
    specparam_declaration7524 specparam_declaration_instance7524();
    specparam_declaration7525 specparam_declaration_instance7525();
    specparam_declaration7526 specparam_declaration_instance7526();
    specparam_declaration7527 specparam_declaration_instance7527();
    specparam_declaration7528 specparam_declaration_instance7528();
    specparam_declaration7529 specparam_declaration_instance7529();
    specparam_declaration7530 specparam_declaration_instance7530();
    specparam_declaration7531 specparam_declaration_instance7531();
    specparam_declaration7532 specparam_declaration_instance7532();
    specparam_declaration7533 specparam_declaration_instance7533();
    specparam_declaration7534 specparam_declaration_instance7534();
    specparam_declaration7535 specparam_declaration_instance7535();
    specparam_declaration7536 specparam_declaration_instance7536();
    specparam_declaration7537 specparam_declaration_instance7537();
    specparam_declaration7538 specparam_declaration_instance7538();
    specparam_declaration7539 specparam_declaration_instance7539();
    specparam_declaration7540 specparam_declaration_instance7540();
    specparam_declaration7541 specparam_declaration_instance7541();
    specparam_declaration7542 specparam_declaration_instance7542();
    specparam_declaration7543 specparam_declaration_instance7543();
    specparam_declaration7544 specparam_declaration_instance7544();
    specparam_declaration7545 specparam_declaration_instance7545();
    specparam_declaration7546 specparam_declaration_instance7546();
    specparam_declaration7547 specparam_declaration_instance7547();
    specparam_declaration7548 specparam_declaration_instance7548();
    specparam_declaration7549 specparam_declaration_instance7549();
    specparam_declaration7550 specparam_declaration_instance7550();
    specparam_declaration7551 specparam_declaration_instance7551();
    specparam_declaration7552 specparam_declaration_instance7552();
    specparam_declaration7553 specparam_declaration_instance7553();
    specparam_declaration7554 specparam_declaration_instance7554();
    specparam_declaration7555 specparam_declaration_instance7555();
    specparam_declaration7556 specparam_declaration_instance7556();
    specparam_declaration7557 specparam_declaration_instance7557();
    specparam_declaration7558 specparam_declaration_instance7558();
    specparam_declaration7559 specparam_declaration_instance7559();
    specparam_declaration7560 specparam_declaration_instance7560();
    specparam_declaration7561 specparam_declaration_instance7561();
    specparam_declaration7562 specparam_declaration_instance7562();
    specparam_declaration7563 specparam_declaration_instance7563();
    specparam_declaration7564 specparam_declaration_instance7564();
    specparam_declaration7565 specparam_declaration_instance7565();
    specparam_declaration7566 specparam_declaration_instance7566();
    specparam_declaration7567 specparam_declaration_instance7567();
    specparam_declaration7568 specparam_declaration_instance7568();
    specparam_declaration7569 specparam_declaration_instance7569();
    specparam_declaration7570 specparam_declaration_instance7570();
    specparam_declaration7571 specparam_declaration_instance7571();
    specparam_declaration7572 specparam_declaration_instance7572();
    specparam_declaration7573 specparam_declaration_instance7573();
    specparam_declaration7574 specparam_declaration_instance7574();
    specparam_declaration7575 specparam_declaration_instance7575();
    specparam_declaration7576 specparam_declaration_instance7576();
    specparam_declaration7577 specparam_declaration_instance7577();
    specparam_declaration7578 specparam_declaration_instance7578();
    specparam_declaration7579 specparam_declaration_instance7579();
    specparam_declaration7580 specparam_declaration_instance7580();
    specparam_declaration7581 specparam_declaration_instance7581();
    specparam_declaration7582 specparam_declaration_instance7582();
    specparam_declaration7583 specparam_declaration_instance7583();
    specparam_declaration7584 specparam_declaration_instance7584();
    specparam_declaration7585 specparam_declaration_instance7585();
    specparam_declaration7586 specparam_declaration_instance7586();
    specparam_declaration7587 specparam_declaration_instance7587();
    specparam_declaration7588 specparam_declaration_instance7588();
    specparam_declaration7589 specparam_declaration_instance7589();
    specparam_declaration7590 specparam_declaration_instance7590();
    specparam_declaration7591 specparam_declaration_instance7591();
    specparam_declaration7592 specparam_declaration_instance7592();
    specparam_declaration7593 specparam_declaration_instance7593();
    specparam_declaration7594 specparam_declaration_instance7594();
    specparam_declaration7595 specparam_declaration_instance7595();
    specparam_declaration7596 specparam_declaration_instance7596();
    specparam_declaration7597 specparam_declaration_instance7597();
    specparam_declaration7598 specparam_declaration_instance7598();
    specparam_declaration7599 specparam_declaration_instance7599();
    specparam_declaration7600 specparam_declaration_instance7600();
    specparam_declaration7601 specparam_declaration_instance7601();
    specparam_declaration7602 specparam_declaration_instance7602();
    specparam_declaration7603 specparam_declaration_instance7603();
    specparam_declaration7604 specparam_declaration_instance7604();
    specparam_declaration7605 specparam_declaration_instance7605();
    specparam_declaration7606 specparam_declaration_instance7606();
    specparam_declaration7607 specparam_declaration_instance7607();
    specparam_declaration7608 specparam_declaration_instance7608();
    specparam_declaration7609 specparam_declaration_instance7609();
    specparam_declaration7610 specparam_declaration_instance7610();
    specparam_declaration7611 specparam_declaration_instance7611();
    specparam_declaration7612 specparam_declaration_instance7612();
    specparam_declaration7613 specparam_declaration_instance7613();
    specparam_declaration7614 specparam_declaration_instance7614();
    specparam_declaration7615 specparam_declaration_instance7615();
    specparam_declaration7616 specparam_declaration_instance7616();
    specparam_declaration7617 specparam_declaration_instance7617();
    specparam_declaration7618 specparam_declaration_instance7618();
    specparam_declaration7619 specparam_declaration_instance7619();
    specparam_declaration7620 specparam_declaration_instance7620();
    specparam_declaration7621 specparam_declaration_instance7621();
    specparam_declaration7622 specparam_declaration_instance7622();
    specparam_declaration7623 specparam_declaration_instance7623();
    specparam_declaration7624 specparam_declaration_instance7624();
    specparam_declaration7625 specparam_declaration_instance7625();
    specparam_declaration7626 specparam_declaration_instance7626();
    specparam_declaration7627 specparam_declaration_instance7627();
    specparam_declaration7628 specparam_declaration_instance7628();
    specparam_declaration7629 specparam_declaration_instance7629();
    specparam_declaration7630 specparam_declaration_instance7630();
    specparam_declaration7631 specparam_declaration_instance7631();
    specparam_declaration7632 specparam_declaration_instance7632();
    specparam_declaration7633 specparam_declaration_instance7633();
    specparam_declaration7634 specparam_declaration_instance7634();
    specparam_declaration7635 specparam_declaration_instance7635();
    specparam_declaration7636 specparam_declaration_instance7636();
    specparam_declaration7637 specparam_declaration_instance7637();
    specparam_declaration7638 specparam_declaration_instance7638();
    specparam_declaration7639 specparam_declaration_instance7639();
    specparam_declaration7640 specparam_declaration_instance7640();
    specparam_declaration7641 specparam_declaration_instance7641();
    specparam_declaration7642 specparam_declaration_instance7642();
    specparam_declaration7643 specparam_declaration_instance7643();
    specparam_declaration7644 specparam_declaration_instance7644();
    specparam_declaration7645 specparam_declaration_instance7645();
    specparam_declaration7646 specparam_declaration_instance7646();
    specparam_declaration7647 specparam_declaration_instance7647();
    specparam_declaration7648 specparam_declaration_instance7648();
    specparam_declaration7649 specparam_declaration_instance7649();
    specparam_declaration7650 specparam_declaration_instance7650();
    specparam_declaration7651 specparam_declaration_instance7651();
    specparam_declaration7652 specparam_declaration_instance7652();
    specparam_declaration7653 specparam_declaration_instance7653();
    specparam_declaration7654 specparam_declaration_instance7654();
    specparam_declaration7655 specparam_declaration_instance7655();
    specparam_declaration7656 specparam_declaration_instance7656();
    specparam_declaration7657 specparam_declaration_instance7657();
    specparam_declaration7658 specparam_declaration_instance7658();
    specparam_declaration7659 specparam_declaration_instance7659();
    specparam_declaration7660 specparam_declaration_instance7660();
    specparam_declaration7661 specparam_declaration_instance7661();
    specparam_declaration7662 specparam_declaration_instance7662();
    specparam_declaration7663 specparam_declaration_instance7663();
    specparam_declaration7664 specparam_declaration_instance7664();
    specparam_declaration7665 specparam_declaration_instance7665();
    specparam_declaration7666 specparam_declaration_instance7666();
    specparam_declaration7667 specparam_declaration_instance7667();
    specparam_declaration7668 specparam_declaration_instance7668();
    specparam_declaration7669 specparam_declaration_instance7669();
    specparam_declaration7670 specparam_declaration_instance7670();
    specparam_declaration7671 specparam_declaration_instance7671();
    specparam_declaration7672 specparam_declaration_instance7672();
    specparam_declaration7673 specparam_declaration_instance7673();
    specparam_declaration7674 specparam_declaration_instance7674();
    specparam_declaration7675 specparam_declaration_instance7675();
    specparam_declaration7676 specparam_declaration_instance7676();
    specparam_declaration7677 specparam_declaration_instance7677();
    specparam_declaration7678 specparam_declaration_instance7678();
    specparam_declaration7679 specparam_declaration_instance7679();
    specparam_declaration7680 specparam_declaration_instance7680();
    specparam_declaration7681 specparam_declaration_instance7681();
    specparam_declaration7682 specparam_declaration_instance7682();
    specparam_declaration7683 specparam_declaration_instance7683();
    specparam_declaration7684 specparam_declaration_instance7684();
    specparam_declaration7685 specparam_declaration_instance7685();
    specparam_declaration7686 specparam_declaration_instance7686();
    specparam_declaration7687 specparam_declaration_instance7687();
    specparam_declaration7688 specparam_declaration_instance7688();
    specparam_declaration7689 specparam_declaration_instance7689();
    specparam_declaration7690 specparam_declaration_instance7690();
    specparam_declaration7691 specparam_declaration_instance7691();
    specparam_declaration7692 specparam_declaration_instance7692();
    specparam_declaration7693 specparam_declaration_instance7693();
    specparam_declaration7694 specparam_declaration_instance7694();
    specparam_declaration7695 specparam_declaration_instance7695();
    specparam_declaration7696 specparam_declaration_instance7696();
    specparam_declaration7697 specparam_declaration_instance7697();
    specparam_declaration7698 specparam_declaration_instance7698();
    specparam_declaration7699 specparam_declaration_instance7699();
    specparam_declaration7700 specparam_declaration_instance7700();
    specparam_declaration7701 specparam_declaration_instance7701();
    specparam_declaration7702 specparam_declaration_instance7702();
    specparam_declaration7703 specparam_declaration_instance7703();
    specparam_declaration7704 specparam_declaration_instance7704();
    specparam_declaration7705 specparam_declaration_instance7705();
    specparam_declaration7706 specparam_declaration_instance7706();
    specparam_declaration7707 specparam_declaration_instance7707();
    specparam_declaration7708 specparam_declaration_instance7708();
    specparam_declaration7709 specparam_declaration_instance7709();
    specparam_declaration7710 specparam_declaration_instance7710();
    specparam_declaration7711 specparam_declaration_instance7711();
    specparam_declaration7712 specparam_declaration_instance7712();
    specparam_declaration7713 specparam_declaration_instance7713();
    specparam_declaration7714 specparam_declaration_instance7714();
    specparam_declaration7715 specparam_declaration_instance7715();
    specparam_declaration7716 specparam_declaration_instance7716();
    specparam_declaration7717 specparam_declaration_instance7717();
    specparam_declaration7718 specparam_declaration_instance7718();
    specparam_declaration7719 specparam_declaration_instance7719();
    specparam_declaration7720 specparam_declaration_instance7720();
    specparam_declaration7721 specparam_declaration_instance7721();
    specparam_declaration7722 specparam_declaration_instance7722();
    specparam_declaration7723 specparam_declaration_instance7723();
    specparam_declaration7724 specparam_declaration_instance7724();
    specparam_declaration7725 specparam_declaration_instance7725();
    specparam_declaration7726 specparam_declaration_instance7726();
    specparam_declaration7727 specparam_declaration_instance7727();
    specparam_declaration7728 specparam_declaration_instance7728();
    specparam_declaration7729 specparam_declaration_instance7729();
    specparam_declaration7730 specparam_declaration_instance7730();
    specparam_declaration7731 specparam_declaration_instance7731();
    specparam_declaration7732 specparam_declaration_instance7732();
    specparam_declaration7733 specparam_declaration_instance7733();
    specparam_declaration7734 specparam_declaration_instance7734();
    specparam_declaration7735 specparam_declaration_instance7735();
    specparam_declaration7736 specparam_declaration_instance7736();
    specparam_declaration7737 specparam_declaration_instance7737();
    specparam_declaration7738 specparam_declaration_instance7738();
    specparam_declaration7739 specparam_declaration_instance7739();
    specparam_declaration7740 specparam_declaration_instance7740();
    specparam_declaration7741 specparam_declaration_instance7741();
    specparam_declaration7742 specparam_declaration_instance7742();
    specparam_declaration7743 specparam_declaration_instance7743();
    specparam_declaration7744 specparam_declaration_instance7744();
    specparam_declaration7745 specparam_declaration_instance7745();
    specparam_declaration7746 specparam_declaration_instance7746();
    specparam_declaration7747 specparam_declaration_instance7747();
    specparam_declaration7748 specparam_declaration_instance7748();
    specparam_declaration7749 specparam_declaration_instance7749();
    specparam_declaration7750 specparam_declaration_instance7750();
    specparam_declaration7751 specparam_declaration_instance7751();
    specparam_declaration7752 specparam_declaration_instance7752();
    specparam_declaration7753 specparam_declaration_instance7753();
    specparam_declaration7754 specparam_declaration_instance7754();
    specparam_declaration7755 specparam_declaration_instance7755();
    specparam_declaration7756 specparam_declaration_instance7756();
    specparam_declaration7757 specparam_declaration_instance7757();
    specparam_declaration7758 specparam_declaration_instance7758();
    specparam_declaration7759 specparam_declaration_instance7759();
    specparam_declaration7760 specparam_declaration_instance7760();
    specparam_declaration7761 specparam_declaration_instance7761();
    specparam_declaration7762 specparam_declaration_instance7762();
    specparam_declaration7763 specparam_declaration_instance7763();
    specparam_declaration7764 specparam_declaration_instance7764();
    specparam_declaration7765 specparam_declaration_instance7765();
    specparam_declaration7766 specparam_declaration_instance7766();
    specparam_declaration7767 specparam_declaration_instance7767();
    specparam_declaration7768 specparam_declaration_instance7768();
    specparam_declaration7769 specparam_declaration_instance7769();
    specparam_declaration7770 specparam_declaration_instance7770();
    specparam_declaration7771 specparam_declaration_instance7771();
    specparam_declaration7772 specparam_declaration_instance7772();
    specparam_declaration7773 specparam_declaration_instance7773();
    specparam_declaration7774 specparam_declaration_instance7774();
    specparam_declaration7775 specparam_declaration_instance7775();
    specparam_declaration7776 specparam_declaration_instance7776();
    specparam_declaration7777 specparam_declaration_instance7777();
    specparam_declaration7778 specparam_declaration_instance7778();
    specparam_declaration7779 specparam_declaration_instance7779();
    specparam_declaration7780 specparam_declaration_instance7780();
    specparam_declaration7781 specparam_declaration_instance7781();
    specparam_declaration7782 specparam_declaration_instance7782();
    specparam_declaration7783 specparam_declaration_instance7783();
    specparam_declaration7784 specparam_declaration_instance7784();
    specparam_declaration7785 specparam_declaration_instance7785();
    specparam_declaration7786 specparam_declaration_instance7786();
    specparam_declaration7787 specparam_declaration_instance7787();
    specparam_declaration7788 specparam_declaration_instance7788();
    specparam_declaration7789 specparam_declaration_instance7789();
    specparam_declaration7790 specparam_declaration_instance7790();
    specparam_declaration7791 specparam_declaration_instance7791();
    specparam_declaration7792 specparam_declaration_instance7792();
    specparam_declaration7793 specparam_declaration_instance7793();
    specparam_declaration7794 specparam_declaration_instance7794();
    specparam_declaration7795 specparam_declaration_instance7795();
    specparam_declaration7796 specparam_declaration_instance7796();
    specparam_declaration7797 specparam_declaration_instance7797();
    specparam_declaration7798 specparam_declaration_instance7798();
    specparam_declaration7799 specparam_declaration_instance7799();
    specparam_declaration7800 specparam_declaration_instance7800();
    specparam_declaration7801 specparam_declaration_instance7801();
    specparam_declaration7802 specparam_declaration_instance7802();
    specparam_declaration7803 specparam_declaration_instance7803();
    specparam_declaration7804 specparam_declaration_instance7804();
    specparam_declaration7805 specparam_declaration_instance7805();
    specparam_declaration7806 specparam_declaration_instance7806();
    specparam_declaration7807 specparam_declaration_instance7807();
    specparam_declaration7808 specparam_declaration_instance7808();
    specparam_declaration7809 specparam_declaration_instance7809();
    specparam_declaration7810 specparam_declaration_instance7810();
    specparam_declaration7811 specparam_declaration_instance7811();
    specparam_declaration7812 specparam_declaration_instance7812();
    specparam_declaration7813 specparam_declaration_instance7813();
    specparam_declaration7814 specparam_declaration_instance7814();
    specparam_declaration7815 specparam_declaration_instance7815();
    specparam_declaration7816 specparam_declaration_instance7816();
    specparam_declaration7817 specparam_declaration_instance7817();
    specparam_declaration7818 specparam_declaration_instance7818();
    specparam_declaration7819 specparam_declaration_instance7819();
    specparam_declaration7820 specparam_declaration_instance7820();
    specparam_declaration7821 specparam_declaration_instance7821();
    specparam_declaration7822 specparam_declaration_instance7822();
    specparam_declaration7823 specparam_declaration_instance7823();
    specparam_declaration7824 specparam_declaration_instance7824();
    specparam_declaration7825 specparam_declaration_instance7825();
    specparam_declaration7826 specparam_declaration_instance7826();
    specparam_declaration7827 specparam_declaration_instance7827();
    specparam_declaration7828 specparam_declaration_instance7828();
    specparam_declaration7829 specparam_declaration_instance7829();
    specparam_declaration7830 specparam_declaration_instance7830();
    specparam_declaration7831 specparam_declaration_instance7831();
    specparam_declaration7832 specparam_declaration_instance7832();
    specparam_declaration7833 specparam_declaration_instance7833();
    specparam_declaration7834 specparam_declaration_instance7834();
    specparam_declaration7835 specparam_declaration_instance7835();
    specparam_declaration7836 specparam_declaration_instance7836();
    specparam_declaration7837 specparam_declaration_instance7837();
    specparam_declaration7838 specparam_declaration_instance7838();
    specparam_declaration7839 specparam_declaration_instance7839();
    specparam_declaration7840 specparam_declaration_instance7840();
    specparam_declaration7841 specparam_declaration_instance7841();
    specparam_declaration7842 specparam_declaration_instance7842();
    specparam_declaration7843 specparam_declaration_instance7843();
    specparam_declaration7844 specparam_declaration_instance7844();
    specparam_declaration7845 specparam_declaration_instance7845();
    specparam_declaration7846 specparam_declaration_instance7846();
    specparam_declaration7847 specparam_declaration_instance7847();
    specparam_declaration7848 specparam_declaration_instance7848();
    specparam_declaration7849 specparam_declaration_instance7849();
    specparam_declaration7850 specparam_declaration_instance7850();
    specparam_declaration7851 specparam_declaration_instance7851();
    specparam_declaration7852 specparam_declaration_instance7852();
    specparam_declaration7853 specparam_declaration_instance7853();
    specparam_declaration7854 specparam_declaration_instance7854();
    specparam_declaration7855 specparam_declaration_instance7855();
    specparam_declaration7856 specparam_declaration_instance7856();
    specparam_declaration7857 specparam_declaration_instance7857();
    specparam_declaration7858 specparam_declaration_instance7858();
    specparam_declaration7859 specparam_declaration_instance7859();
    specparam_declaration7860 specparam_declaration_instance7860();
    specparam_declaration7861 specparam_declaration_instance7861();
    specparam_declaration7862 specparam_declaration_instance7862();
    specparam_declaration7863 specparam_declaration_instance7863();
    specparam_declaration7864 specparam_declaration_instance7864();
    specparam_declaration7865 specparam_declaration_instance7865();
    specparam_declaration7866 specparam_declaration_instance7866();
    specparam_declaration7867 specparam_declaration_instance7867();
    specparam_declaration7868 specparam_declaration_instance7868();
    specparam_declaration7869 specparam_declaration_instance7869();
    specparam_declaration7870 specparam_declaration_instance7870();
    specparam_declaration7871 specparam_declaration_instance7871();
    specparam_declaration7872 specparam_declaration_instance7872();
    specparam_declaration7873 specparam_declaration_instance7873();
    specparam_declaration7874 specparam_declaration_instance7874();
    specparam_declaration7875 specparam_declaration_instance7875();
    specparam_declaration7876 specparam_declaration_instance7876();
    specparam_declaration7877 specparam_declaration_instance7877();
    specparam_declaration7878 specparam_declaration_instance7878();
    specparam_declaration7879 specparam_declaration_instance7879();
    specparam_declaration7880 specparam_declaration_instance7880();
    specparam_declaration7881 specparam_declaration_instance7881();
    specparam_declaration7882 specparam_declaration_instance7882();
    specparam_declaration7883 specparam_declaration_instance7883();
    specparam_declaration7884 specparam_declaration_instance7884();
    specparam_declaration7885 specparam_declaration_instance7885();
    specparam_declaration7886 specparam_declaration_instance7886();
    specparam_declaration7887 specparam_declaration_instance7887();
    specparam_declaration7888 specparam_declaration_instance7888();
    specparam_declaration7889 specparam_declaration_instance7889();
    specparam_declaration7890 specparam_declaration_instance7890();
    specparam_declaration7891 specparam_declaration_instance7891();
    specparam_declaration7892 specparam_declaration_instance7892();
    specparam_declaration7893 specparam_declaration_instance7893();
    specparam_declaration7894 specparam_declaration_instance7894();
    specparam_declaration7895 specparam_declaration_instance7895();
    specparam_declaration7896 specparam_declaration_instance7896();
    specparam_declaration7897 specparam_declaration_instance7897();
    specparam_declaration7898 specparam_declaration_instance7898();
    specparam_declaration7899 specparam_declaration_instance7899();
    specparam_declaration7900 specparam_declaration_instance7900();
    specparam_declaration7901 specparam_declaration_instance7901();
    specparam_declaration7902 specparam_declaration_instance7902();
    specparam_declaration7903 specparam_declaration_instance7903();
    specparam_declaration7904 specparam_declaration_instance7904();
    specparam_declaration7905 specparam_declaration_instance7905();
    specparam_declaration7906 specparam_declaration_instance7906();
    specparam_declaration7907 specparam_declaration_instance7907();
    specparam_declaration7908 specparam_declaration_instance7908();
    specparam_declaration7909 specparam_declaration_instance7909();
    specparam_declaration7910 specparam_declaration_instance7910();
    specparam_declaration7911 specparam_declaration_instance7911();
    specparam_declaration7912 specparam_declaration_instance7912();
    specparam_declaration7913 specparam_declaration_instance7913();
    specparam_declaration7914 specparam_declaration_instance7914();
    specparam_declaration7915 specparam_declaration_instance7915();
    specparam_declaration7916 specparam_declaration_instance7916();
    specparam_declaration7917 specparam_declaration_instance7917();
    specparam_declaration7918 specparam_declaration_instance7918();
    specparam_declaration7919 specparam_declaration_instance7919();
    specparam_declaration7920 specparam_declaration_instance7920();
    specparam_declaration7921 specparam_declaration_instance7921();
    specparam_declaration7922 specparam_declaration_instance7922();
    specparam_declaration7923 specparam_declaration_instance7923();
    specparam_declaration7924 specparam_declaration_instance7924();
    specparam_declaration7925 specparam_declaration_instance7925();
    specparam_declaration7926 specparam_declaration_instance7926();
    specparam_declaration7927 specparam_declaration_instance7927();
    specparam_declaration7928 specparam_declaration_instance7928();
    specparam_declaration7929 specparam_declaration_instance7929();
    specparam_declaration7930 specparam_declaration_instance7930();
    specparam_declaration7931 specparam_declaration_instance7931();
    specparam_declaration7932 specparam_declaration_instance7932();
    specparam_declaration7933 specparam_declaration_instance7933();
    specparam_declaration7934 specparam_declaration_instance7934();
    specparam_declaration7935 specparam_declaration_instance7935();
    specparam_declaration7936 specparam_declaration_instance7936();
    specparam_declaration7937 specparam_declaration_instance7937();
    specparam_declaration7938 specparam_declaration_instance7938();
    specparam_declaration7939 specparam_declaration_instance7939();
    specparam_declaration7940 specparam_declaration_instance7940();
    specparam_declaration7941 specparam_declaration_instance7941();
    specparam_declaration7942 specparam_declaration_instance7942();
    specparam_declaration7943 specparam_declaration_instance7943();
    specparam_declaration7944 specparam_declaration_instance7944();
    specparam_declaration7945 specparam_declaration_instance7945();
    specparam_declaration7946 specparam_declaration_instance7946();
    specparam_declaration7947 specparam_declaration_instance7947();
    specparam_declaration7948 specparam_declaration_instance7948();
    specparam_declaration7949 specparam_declaration_instance7949();
    specparam_declaration7950 specparam_declaration_instance7950();
    specparam_declaration7951 specparam_declaration_instance7951();
    specparam_declaration7952 specparam_declaration_instance7952();
    specparam_declaration7953 specparam_declaration_instance7953();
    specparam_declaration7954 specparam_declaration_instance7954();
    specparam_declaration7955 specparam_declaration_instance7955();
    specparam_declaration7956 specparam_declaration_instance7956();
    specparam_declaration7957 specparam_declaration_instance7957();
    specparam_declaration7958 specparam_declaration_instance7958();
    specparam_declaration7959 specparam_declaration_instance7959();
    specparam_declaration7960 specparam_declaration_instance7960();
    specparam_declaration7961 specparam_declaration_instance7961();
    specparam_declaration7962 specparam_declaration_instance7962();
    specparam_declaration7963 specparam_declaration_instance7963();
    specparam_declaration7964 specparam_declaration_instance7964();
    specparam_declaration7965 specparam_declaration_instance7965();
    specparam_declaration7966 specparam_declaration_instance7966();
    specparam_declaration7967 specparam_declaration_instance7967();
    specparam_declaration7968 specparam_declaration_instance7968();
    specparam_declaration7969 specparam_declaration_instance7969();
    specparam_declaration7970 specparam_declaration_instance7970();
    specparam_declaration7971 specparam_declaration_instance7971();
    specparam_declaration7972 specparam_declaration_instance7972();
    specparam_declaration7973 specparam_declaration_instance7973();
    specparam_declaration7974 specparam_declaration_instance7974();
    specparam_declaration7975 specparam_declaration_instance7975();
    specparam_declaration7976 specparam_declaration_instance7976();
    specparam_declaration7977 specparam_declaration_instance7977();
    specparam_declaration7978 specparam_declaration_instance7978();
    specparam_declaration7979 specparam_declaration_instance7979();
    specparam_declaration7980 specparam_declaration_instance7980();
    specparam_declaration7981 specparam_declaration_instance7981();
    specparam_declaration7982 specparam_declaration_instance7982();
    specparam_declaration7983 specparam_declaration_instance7983();
    specparam_declaration7984 specparam_declaration_instance7984();
    specparam_declaration7985 specparam_declaration_instance7985();
    specparam_declaration7986 specparam_declaration_instance7986();
    specparam_declaration7987 specparam_declaration_instance7987();
    specparam_declaration7988 specparam_declaration_instance7988();
    specparam_declaration7989 specparam_declaration_instance7989();
    specparam_declaration7990 specparam_declaration_instance7990();
    specparam_declaration7991 specparam_declaration_instance7991();
    specparam_declaration7992 specparam_declaration_instance7992();
    specparam_declaration7993 specparam_declaration_instance7993();
    specparam_declaration7994 specparam_declaration_instance7994();
    specparam_declaration7995 specparam_declaration_instance7995();
    specparam_declaration7996 specparam_declaration_instance7996();
    specparam_declaration7997 specparam_declaration_instance7997();
    specparam_declaration7998 specparam_declaration_instance7998();
    specparam_declaration7999 specparam_declaration_instance7999();
    specparam_declaration8000 specparam_declaration_instance8000();
    specparam_declaration8001 specparam_declaration_instance8001();
    specparam_declaration8002 specparam_declaration_instance8002();
    specparam_declaration8003 specparam_declaration_instance8003();
    specparam_declaration8004 specparam_declaration_instance8004();
    specparam_declaration8005 specparam_declaration_instance8005();
    specparam_declaration8006 specparam_declaration_instance8006();
    specparam_declaration8007 specparam_declaration_instance8007();
    specparam_declaration8008 specparam_declaration_instance8008();
    specparam_declaration8009 specparam_declaration_instance8009();
    specparam_declaration8010 specparam_declaration_instance8010();
    specparam_declaration8011 specparam_declaration_instance8011();
    specparam_declaration8012 specparam_declaration_instance8012();
    specparam_declaration8013 specparam_declaration_instance8013();
    specparam_declaration8014 specparam_declaration_instance8014();
    specparam_declaration8015 specparam_declaration_instance8015();
    specparam_declaration8016 specparam_declaration_instance8016();
    specparam_declaration8017 specparam_declaration_instance8017();
    specparam_declaration8018 specparam_declaration_instance8018();
    specparam_declaration8019 specparam_declaration_instance8019();
    specparam_declaration8020 specparam_declaration_instance8020();
    specparam_declaration8021 specparam_declaration_instance8021();
    specparam_declaration8022 specparam_declaration_instance8022();
    specparam_declaration8023 specparam_declaration_instance8023();
    specparam_declaration8024 specparam_declaration_instance8024();
    specparam_declaration8025 specparam_declaration_instance8025();
    specparam_declaration8026 specparam_declaration_instance8026();
    specparam_declaration8027 specparam_declaration_instance8027();
    specparam_declaration8028 specparam_declaration_instance8028();
    specparam_declaration8029 specparam_declaration_instance8029();
    specparam_declaration8030 specparam_declaration_instance8030();
    specparam_declaration8031 specparam_declaration_instance8031();
    specparam_declaration8032 specparam_declaration_instance8032();
    specparam_declaration8033 specparam_declaration_instance8033();
    specparam_declaration8034 specparam_declaration_instance8034();
    specparam_declaration8035 specparam_declaration_instance8035();
    specparam_declaration8036 specparam_declaration_instance8036();
    specparam_declaration8037 specparam_declaration_instance8037();
    specparam_declaration8038 specparam_declaration_instance8038();
    specparam_declaration8039 specparam_declaration_instance8039();
    specparam_declaration8040 specparam_declaration_instance8040();
    specparam_declaration8041 specparam_declaration_instance8041();
    specparam_declaration8042 specparam_declaration_instance8042();
    specparam_declaration8043 specparam_declaration_instance8043();
    specparam_declaration8044 specparam_declaration_instance8044();
    specparam_declaration8045 specparam_declaration_instance8045();
    specparam_declaration8046 specparam_declaration_instance8046();
    specparam_declaration8047 specparam_declaration_instance8047();
    specparam_declaration8048 specparam_declaration_instance8048();
    specparam_declaration8049 specparam_declaration_instance8049();
    specparam_declaration8050 specparam_declaration_instance8050();
    specparam_declaration8051 specparam_declaration_instance8051();
    specparam_declaration8052 specparam_declaration_instance8052();
    specparam_declaration8053 specparam_declaration_instance8053();
    specparam_declaration8054 specparam_declaration_instance8054();
    specparam_declaration8055 specparam_declaration_instance8055();
    specparam_declaration8056 specparam_declaration_instance8056();
    specparam_declaration8057 specparam_declaration_instance8057();
    specparam_declaration8058 specparam_declaration_instance8058();
    specparam_declaration8059 specparam_declaration_instance8059();
    specparam_declaration8060 specparam_declaration_instance8060();
    specparam_declaration8061 specparam_declaration_instance8061();
    specparam_declaration8062 specparam_declaration_instance8062();
    specparam_declaration8063 specparam_declaration_instance8063();
    specparam_declaration8064 specparam_declaration_instance8064();
    specparam_declaration8065 specparam_declaration_instance8065();
    specparam_declaration8066 specparam_declaration_instance8066();
    specparam_declaration8067 specparam_declaration_instance8067();
    specparam_declaration8068 specparam_declaration_instance8068();
    specparam_declaration8069 specparam_declaration_instance8069();
    specparam_declaration8070 specparam_declaration_instance8070();
    specparam_declaration8071 specparam_declaration_instance8071();
    specparam_declaration8072 specparam_declaration_instance8072();
    specparam_declaration8073 specparam_declaration_instance8073();
    specparam_declaration8074 specparam_declaration_instance8074();
    specparam_declaration8075 specparam_declaration_instance8075();
    specparam_declaration8076 specparam_declaration_instance8076();
    specparam_declaration8077 specparam_declaration_instance8077();
    specparam_declaration8078 specparam_declaration_instance8078();
    specparam_declaration8079 specparam_declaration_instance8079();
    specparam_declaration8080 specparam_declaration_instance8080();
    specparam_declaration8081 specparam_declaration_instance8081();
    specparam_declaration8082 specparam_declaration_instance8082();
    specparam_declaration8083 specparam_declaration_instance8083();
    specparam_declaration8084 specparam_declaration_instance8084();
    specparam_declaration8085 specparam_declaration_instance8085();
    specparam_declaration8086 specparam_declaration_instance8086();
    specparam_declaration8087 specparam_declaration_instance8087();
    specparam_declaration8088 specparam_declaration_instance8088();
    specparam_declaration8089 specparam_declaration_instance8089();
    specparam_declaration8090 specparam_declaration_instance8090();
    specparam_declaration8091 specparam_declaration_instance8091();
    specparam_declaration8092 specparam_declaration_instance8092();
    specparam_declaration8093 specparam_declaration_instance8093();
    specparam_declaration8094 specparam_declaration_instance8094();
    specparam_declaration8095 specparam_declaration_instance8095();
    specparam_declaration8096 specparam_declaration_instance8096();
    specparam_declaration8097 specparam_declaration_instance8097();
    specparam_declaration8098 specparam_declaration_instance8098();
    specparam_declaration8099 specparam_declaration_instance8099();
    specparam_declaration8100 specparam_declaration_instance8100();
    specparam_declaration8101 specparam_declaration_instance8101();
    specparam_declaration8102 specparam_declaration_instance8102();
    specparam_declaration8103 specparam_declaration_instance8103();
    specparam_declaration8104 specparam_declaration_instance8104();
    specparam_declaration8105 specparam_declaration_instance8105();
    specparam_declaration8106 specparam_declaration_instance8106();
    specparam_declaration8107 specparam_declaration_instance8107();
    specparam_declaration8108 specparam_declaration_instance8108();
    specparam_declaration8109 specparam_declaration_instance8109();
    specparam_declaration8110 specparam_declaration_instance8110();
    specparam_declaration8111 specparam_declaration_instance8111();
    specparam_declaration8112 specparam_declaration_instance8112();
    specparam_declaration8113 specparam_declaration_instance8113();
    specparam_declaration8114 specparam_declaration_instance8114();
    specparam_declaration8115 specparam_declaration_instance8115();
    specparam_declaration8116 specparam_declaration_instance8116();
    specparam_declaration8117 specparam_declaration_instance8117();
    specparam_declaration8118 specparam_declaration_instance8118();
    specparam_declaration8119 specparam_declaration_instance8119();
    specparam_declaration8120 specparam_declaration_instance8120();
    specparam_declaration8121 specparam_declaration_instance8121();
    specparam_declaration8122 specparam_declaration_instance8122();
    specparam_declaration8123 specparam_declaration_instance8123();
    specparam_declaration8124 specparam_declaration_instance8124();
    specparam_declaration8125 specparam_declaration_instance8125();
    specparam_declaration8126 specparam_declaration_instance8126();
    specparam_declaration8127 specparam_declaration_instance8127();
    specparam_declaration8128 specparam_declaration_instance8128();
    specparam_declaration8129 specparam_declaration_instance8129();
    specparam_declaration8130 specparam_declaration_instance8130();
    specparam_declaration8131 specparam_declaration_instance8131();
    specparam_declaration8132 specparam_declaration_instance8132();
    specparam_declaration8133 specparam_declaration_instance8133();
    specparam_declaration8134 specparam_declaration_instance8134();
    specparam_declaration8135 specparam_declaration_instance8135();
    specparam_declaration8136 specparam_declaration_instance8136();
    specparam_declaration8137 specparam_declaration_instance8137();
    specparam_declaration8138 specparam_declaration_instance8138();
    specparam_declaration8139 specparam_declaration_instance8139();
    specparam_declaration8140 specparam_declaration_instance8140();
    specparam_declaration8141 specparam_declaration_instance8141();
    specparam_declaration8142 specparam_declaration_instance8142();
    specparam_declaration8143 specparam_declaration_instance8143();
    specparam_declaration8144 specparam_declaration_instance8144();
    specparam_declaration8145 specparam_declaration_instance8145();
    specparam_declaration8146 specparam_declaration_instance8146();
    specparam_declaration8147 specparam_declaration_instance8147();
    specparam_declaration8148 specparam_declaration_instance8148();
    specparam_declaration8149 specparam_declaration_instance8149();
    specparam_declaration8150 specparam_declaration_instance8150();
    specparam_declaration8151 specparam_declaration_instance8151();
    specparam_declaration8152 specparam_declaration_instance8152();
    specparam_declaration8153 specparam_declaration_instance8153();
    specparam_declaration8154 specparam_declaration_instance8154();
    specparam_declaration8155 specparam_declaration_instance8155();
    specparam_declaration8156 specparam_declaration_instance8156();
    specparam_declaration8157 specparam_declaration_instance8157();
    specparam_declaration8158 specparam_declaration_instance8158();
    specparam_declaration8159 specparam_declaration_instance8159();
    specparam_declaration8160 specparam_declaration_instance8160();
    specparam_declaration8161 specparam_declaration_instance8161();
    specparam_declaration8162 specparam_declaration_instance8162();
    specparam_declaration8163 specparam_declaration_instance8163();
    specparam_declaration8164 specparam_declaration_instance8164();
    specparam_declaration8165 specparam_declaration_instance8165();
    specparam_declaration8166 specparam_declaration_instance8166();
    specparam_declaration8167 specparam_declaration_instance8167();
    specparam_declaration8168 specparam_declaration_instance8168();
    specparam_declaration8169 specparam_declaration_instance8169();
    specparam_declaration8170 specparam_declaration_instance8170();
    specparam_declaration8171 specparam_declaration_instance8171();
    specparam_declaration8172 specparam_declaration_instance8172();
    specparam_declaration8173 specparam_declaration_instance8173();
    specparam_declaration8174 specparam_declaration_instance8174();
    specparam_declaration8175 specparam_declaration_instance8175();
    specparam_declaration8176 specparam_declaration_instance8176();
    specparam_declaration8177 specparam_declaration_instance8177();
    specparam_declaration8178 specparam_declaration_instance8178();
    specparam_declaration8179 specparam_declaration_instance8179();
    specparam_declaration8180 specparam_declaration_instance8180();
    specparam_declaration8181 specparam_declaration_instance8181();
    specparam_declaration8182 specparam_declaration_instance8182();
    specparam_declaration8183 specparam_declaration_instance8183();
    specparam_declaration8184 specparam_declaration_instance8184();
    specparam_declaration8185 specparam_declaration_instance8185();
    specparam_declaration8186 specparam_declaration_instance8186();
    specparam_declaration8187 specparam_declaration_instance8187();
    specparam_declaration8188 specparam_declaration_instance8188();
    specparam_declaration8189 specparam_declaration_instance8189();
    specparam_declaration8190 specparam_declaration_instance8190();
    specparam_declaration8191 specparam_declaration_instance8191();
    specparam_declaration8192 specparam_declaration_instance8192();
    specparam_declaration8193 specparam_declaration_instance8193();
    specparam_declaration8194 specparam_declaration_instance8194();
    specparam_declaration8195 specparam_declaration_instance8195();
    specparam_declaration8196 specparam_declaration_instance8196();
    specparam_declaration8197 specparam_declaration_instance8197();
    specparam_declaration8198 specparam_declaration_instance8198();
    specparam_declaration8199 specparam_declaration_instance8199();
    specparam_declaration8200 specparam_declaration_instance8200();
    specparam_declaration8201 specparam_declaration_instance8201();
    specparam_declaration8202 specparam_declaration_instance8202();
    specparam_declaration8203 specparam_declaration_instance8203();
    specparam_declaration8204 specparam_declaration_instance8204();
    specparam_declaration8205 specparam_declaration_instance8205();
    specparam_declaration8206 specparam_declaration_instance8206();
    specparam_declaration8207 specparam_declaration_instance8207();
    specparam_declaration8208 specparam_declaration_instance8208();
    specparam_declaration8209 specparam_declaration_instance8209();
    specparam_declaration8210 specparam_declaration_instance8210();
    specparam_declaration8211 specparam_declaration_instance8211();
    specparam_declaration8212 specparam_declaration_instance8212();
    specparam_declaration8213 specparam_declaration_instance8213();
    specparam_declaration8214 specparam_declaration_instance8214();
    specparam_declaration8215 specparam_declaration_instance8215();
    specparam_declaration8216 specparam_declaration_instance8216();
    specparam_declaration8217 specparam_declaration_instance8217();
    specparam_declaration8218 specparam_declaration_instance8218();
    specparam_declaration8219 specparam_declaration_instance8219();
    specparam_declaration8220 specparam_declaration_instance8220();
    specparam_declaration8221 specparam_declaration_instance8221();
    specparam_declaration8222 specparam_declaration_instance8222();
    specparam_declaration8223 specparam_declaration_instance8223();
    specparam_declaration8224 specparam_declaration_instance8224();
    specparam_declaration8225 specparam_declaration_instance8225();
    specparam_declaration8226 specparam_declaration_instance8226();
    specparam_declaration8227 specparam_declaration_instance8227();
    specparam_declaration8228 specparam_declaration_instance8228();
    specparam_declaration8229 specparam_declaration_instance8229();
    specparam_declaration8230 specparam_declaration_instance8230();
    specparam_declaration8231 specparam_declaration_instance8231();
    specparam_declaration8232 specparam_declaration_instance8232();
    specparam_declaration8233 specparam_declaration_instance8233();
    specparam_declaration8234 specparam_declaration_instance8234();
    specparam_declaration8235 specparam_declaration_instance8235();
    specparam_declaration8236 specparam_declaration_instance8236();
    specparam_declaration8237 specparam_declaration_instance8237();
    specparam_declaration8238 specparam_declaration_instance8238();
    specparam_declaration8239 specparam_declaration_instance8239();
    specparam_declaration8240 specparam_declaration_instance8240();
    specparam_declaration8241 specparam_declaration_instance8241();
    specparam_declaration8242 specparam_declaration_instance8242();
    specparam_declaration8243 specparam_declaration_instance8243();
    specparam_declaration8244 specparam_declaration_instance8244();
    specparam_declaration8245 specparam_declaration_instance8245();
    specparam_declaration8246 specparam_declaration_instance8246();
    specparam_declaration8247 specparam_declaration_instance8247();
    specparam_declaration8248 specparam_declaration_instance8248();
    specparam_declaration8249 specparam_declaration_instance8249();
    specparam_declaration8250 specparam_declaration_instance8250();
    specparam_declaration8251 specparam_declaration_instance8251();
    specparam_declaration8252 specparam_declaration_instance8252();
    specparam_declaration8253 specparam_declaration_instance8253();
    specparam_declaration8254 specparam_declaration_instance8254();
    specparam_declaration8255 specparam_declaration_instance8255();
    specparam_declaration8256 specparam_declaration_instance8256();
    specparam_declaration8257 specparam_declaration_instance8257();
    specparam_declaration8258 specparam_declaration_instance8258();
    specparam_declaration8259 specparam_declaration_instance8259();
    specparam_declaration8260 specparam_declaration_instance8260();
    specparam_declaration8261 specparam_declaration_instance8261();
    specparam_declaration8262 specparam_declaration_instance8262();
    specparam_declaration8263 specparam_declaration_instance8263();
    specparam_declaration8264 specparam_declaration_instance8264();
    specparam_declaration8265 specparam_declaration_instance8265();
    specparam_declaration8266 specparam_declaration_instance8266();
    specparam_declaration8267 specparam_declaration_instance8267();
    specparam_declaration8268 specparam_declaration_instance8268();
    specparam_declaration8269 specparam_declaration_instance8269();
    specparam_declaration8270 specparam_declaration_instance8270();
    specparam_declaration8271 specparam_declaration_instance8271();
    specparam_declaration8272 specparam_declaration_instance8272();
    specparam_declaration8273 specparam_declaration_instance8273();
    specparam_declaration8274 specparam_declaration_instance8274();
    specparam_declaration8275 specparam_declaration_instance8275();
    specparam_declaration8276 specparam_declaration_instance8276();
    specparam_declaration8277 specparam_declaration_instance8277();
    specparam_declaration8278 specparam_declaration_instance8278();
    specparam_declaration8279 specparam_declaration_instance8279();
    specparam_declaration8280 specparam_declaration_instance8280();
    specparam_declaration8281 specparam_declaration_instance8281();
    specparam_declaration8282 specparam_declaration_instance8282();
    specparam_declaration8283 specparam_declaration_instance8283();
    specparam_declaration8284 specparam_declaration_instance8284();
    specparam_declaration8285 specparam_declaration_instance8285();
    specparam_declaration8286 specparam_declaration_instance8286();
    specparam_declaration8287 specparam_declaration_instance8287();
    specparam_declaration8288 specparam_declaration_instance8288();
    specparam_declaration8289 specparam_declaration_instance8289();
    specparam_declaration8290 specparam_declaration_instance8290();
    specparam_declaration8291 specparam_declaration_instance8291();
    specparam_declaration8292 specparam_declaration_instance8292();
    specparam_declaration8293 specparam_declaration_instance8293();
    specparam_declaration8294 specparam_declaration_instance8294();
    specparam_declaration8295 specparam_declaration_instance8295();
    specparam_declaration8296 specparam_declaration_instance8296();
    specparam_declaration8297 specparam_declaration_instance8297();
    specparam_declaration8298 specparam_declaration_instance8298();
    specparam_declaration8299 specparam_declaration_instance8299();
    specparam_declaration8300 specparam_declaration_instance8300();
    specparam_declaration8301 specparam_declaration_instance8301();
    specparam_declaration8302 specparam_declaration_instance8302();
    specparam_declaration8303 specparam_declaration_instance8303();
    specparam_declaration8304 specparam_declaration_instance8304();
    specparam_declaration8305 specparam_declaration_instance8305();
    specparam_declaration8306 specparam_declaration_instance8306();
    specparam_declaration8307 specparam_declaration_instance8307();
    specparam_declaration8308 specparam_declaration_instance8308();
    specparam_declaration8309 specparam_declaration_instance8309();
    specparam_declaration8310 specparam_declaration_instance8310();
    specparam_declaration8311 specparam_declaration_instance8311();
    specparam_declaration8312 specparam_declaration_instance8312();
    specparam_declaration8313 specparam_declaration_instance8313();
    specparam_declaration8314 specparam_declaration_instance8314();
    specparam_declaration8315 specparam_declaration_instance8315();
    specparam_declaration8316 specparam_declaration_instance8316();
    specparam_declaration8317 specparam_declaration_instance8317();
    specparam_declaration8318 specparam_declaration_instance8318();
    specparam_declaration8319 specparam_declaration_instance8319();
    specparam_declaration8320 specparam_declaration_instance8320();
    specparam_declaration8321 specparam_declaration_instance8321();
    specparam_declaration8322 specparam_declaration_instance8322();
    specparam_declaration8323 specparam_declaration_instance8323();
    specparam_declaration8324 specparam_declaration_instance8324();
    specparam_declaration8325 specparam_declaration_instance8325();
    specparam_declaration8326 specparam_declaration_instance8326();
    specparam_declaration8327 specparam_declaration_instance8327();
    specparam_declaration8328 specparam_declaration_instance8328();
    specparam_declaration8329 specparam_declaration_instance8329();
    specparam_declaration8330 specparam_declaration_instance8330();
    specparam_declaration8331 specparam_declaration_instance8331();
    specparam_declaration8332 specparam_declaration_instance8332();
    specparam_declaration8333 specparam_declaration_instance8333();
    specparam_declaration8334 specparam_declaration_instance8334();
    specparam_declaration8335 specparam_declaration_instance8335();
    specparam_declaration8336 specparam_declaration_instance8336();
    specparam_declaration8337 specparam_declaration_instance8337();
    specparam_declaration8338 specparam_declaration_instance8338();
    specparam_declaration8339 specparam_declaration_instance8339();
    specparam_declaration8340 specparam_declaration_instance8340();
    specparam_declaration8341 specparam_declaration_instance8341();
    specparam_declaration8342 specparam_declaration_instance8342();
    specparam_declaration8343 specparam_declaration_instance8343();
    specparam_declaration8344 specparam_declaration_instance8344();
    specparam_declaration8345 specparam_declaration_instance8345();
    specparam_declaration8346 specparam_declaration_instance8346();
    specparam_declaration8347 specparam_declaration_instance8347();
    specparam_declaration8348 specparam_declaration_instance8348();
    specparam_declaration8349 specparam_declaration_instance8349();
    specparam_declaration8350 specparam_declaration_instance8350();
    specparam_declaration8351 specparam_declaration_instance8351();
    specparam_declaration8352 specparam_declaration_instance8352();
    specparam_declaration8353 specparam_declaration_instance8353();
    specparam_declaration8354 specparam_declaration_instance8354();
    specparam_declaration8355 specparam_declaration_instance8355();
    specparam_declaration8356 specparam_declaration_instance8356();
    specparam_declaration8357 specparam_declaration_instance8357();
    specparam_declaration8358 specparam_declaration_instance8358();
    specparam_declaration8359 specparam_declaration_instance8359();
    specparam_declaration8360 specparam_declaration_instance8360();
    specparam_declaration8361 specparam_declaration_instance8361();
    specparam_declaration8362 specparam_declaration_instance8362();
    specparam_declaration8363 specparam_declaration_instance8363();
    specparam_declaration8364 specparam_declaration_instance8364();
    specparam_declaration8365 specparam_declaration_instance8365();
    specparam_declaration8366 specparam_declaration_instance8366();
    specparam_declaration8367 specparam_declaration_instance8367();
    specparam_declaration8368 specparam_declaration_instance8368();
    specparam_declaration8369 specparam_declaration_instance8369();
    specparam_declaration8370 specparam_declaration_instance8370();
    specparam_declaration8371 specparam_declaration_instance8371();
    specparam_declaration8372 specparam_declaration_instance8372();
    specparam_declaration8373 specparam_declaration_instance8373();
    specparam_declaration8374 specparam_declaration_instance8374();
    specparam_declaration8375 specparam_declaration_instance8375();
    specparam_declaration8376 specparam_declaration_instance8376();
    specparam_declaration8377 specparam_declaration_instance8377();
    specparam_declaration8378 specparam_declaration_instance8378();
    specparam_declaration8379 specparam_declaration_instance8379();
    specparam_declaration8380 specparam_declaration_instance8380();
    specparam_declaration8381 specparam_declaration_instance8381();
    specparam_declaration8382 specparam_declaration_instance8382();
    specparam_declaration8383 specparam_declaration_instance8383();
    specparam_declaration8384 specparam_declaration_instance8384();
    specparam_declaration8385 specparam_declaration_instance8385();
    specparam_declaration8386 specparam_declaration_instance8386();
    specparam_declaration8387 specparam_declaration_instance8387();
    specparam_declaration8388 specparam_declaration_instance8388();
    specparam_declaration8389 specparam_declaration_instance8389();
    specparam_declaration8390 specparam_declaration_instance8390();
    specparam_declaration8391 specparam_declaration_instance8391();
    specparam_declaration8392 specparam_declaration_instance8392();
    specparam_declaration8393 specparam_declaration_instance8393();
    specparam_declaration8394 specparam_declaration_instance8394();
    specparam_declaration8395 specparam_declaration_instance8395();
    specparam_declaration8396 specparam_declaration_instance8396();
    specparam_declaration8397 specparam_declaration_instance8397();
    specparam_declaration8398 specparam_declaration_instance8398();
    specparam_declaration8399 specparam_declaration_instance8399();
    specparam_declaration8400 specparam_declaration_instance8400();
    specparam_declaration8401 specparam_declaration_instance8401();
    specparam_declaration8402 specparam_declaration_instance8402();
    specparam_declaration8403 specparam_declaration_instance8403();
    specparam_declaration8404 specparam_declaration_instance8404();
    specparam_declaration8405 specparam_declaration_instance8405();
    specparam_declaration8406 specparam_declaration_instance8406();
    specparam_declaration8407 specparam_declaration_instance8407();
    specparam_declaration8408 specparam_declaration_instance8408();
    specparam_declaration8409 specparam_declaration_instance8409();
    specparam_declaration8410 specparam_declaration_instance8410();
    specparam_declaration8411 specparam_declaration_instance8411();
    specparam_declaration8412 specparam_declaration_instance8412();
    specparam_declaration8413 specparam_declaration_instance8413();
    specparam_declaration8414 specparam_declaration_instance8414();
    specparam_declaration8415 specparam_declaration_instance8415();
    specparam_declaration8416 specparam_declaration_instance8416();
    specparam_declaration8417 specparam_declaration_instance8417();
    specparam_declaration8418 specparam_declaration_instance8418();
    specparam_declaration8419 specparam_declaration_instance8419();
    specparam_declaration8420 specparam_declaration_instance8420();
    specparam_declaration8421 specparam_declaration_instance8421();
    specparam_declaration8422 specparam_declaration_instance8422();
    specparam_declaration8423 specparam_declaration_instance8423();
    specparam_declaration8424 specparam_declaration_instance8424();
    specparam_declaration8425 specparam_declaration_instance8425();
    specparam_declaration8426 specparam_declaration_instance8426();
    specparam_declaration8427 specparam_declaration_instance8427();
    specparam_declaration8428 specparam_declaration_instance8428();
    specparam_declaration8429 specparam_declaration_instance8429();
    specparam_declaration8430 specparam_declaration_instance8430();
    specparam_declaration8431 specparam_declaration_instance8431();
    specparam_declaration8432 specparam_declaration_instance8432();
    specparam_declaration8433 specparam_declaration_instance8433();
    specparam_declaration8434 specparam_declaration_instance8434();
    specparam_declaration8435 specparam_declaration_instance8435();
    specparam_declaration8436 specparam_declaration_instance8436();
    specparam_declaration8437 specparam_declaration_instance8437();
    specparam_declaration8438 specparam_declaration_instance8438();
    specparam_declaration8439 specparam_declaration_instance8439();
    specparam_declaration8440 specparam_declaration_instance8440();
    specparam_declaration8441 specparam_declaration_instance8441();
    specparam_declaration8442 specparam_declaration_instance8442();
    specparam_declaration8443 specparam_declaration_instance8443();
    specparam_declaration8444 specparam_declaration_instance8444();
    specparam_declaration8445 specparam_declaration_instance8445();
    specparam_declaration8446 specparam_declaration_instance8446();
    specparam_declaration8447 specparam_declaration_instance8447();
    specparam_declaration8448 specparam_declaration_instance8448();
    specparam_declaration8449 specparam_declaration_instance8449();
    specparam_declaration8450 specparam_declaration_instance8450();
    specparam_declaration8451 specparam_declaration_instance8451();
    specparam_declaration8452 specparam_declaration_instance8452();
    specparam_declaration8453 specparam_declaration_instance8453();
    specparam_declaration8454 specparam_declaration_instance8454();
    specparam_declaration8455 specparam_declaration_instance8455();
    specparam_declaration8456 specparam_declaration_instance8456();
    specparam_declaration8457 specparam_declaration_instance8457();
    specparam_declaration8458 specparam_declaration_instance8458();
    specparam_declaration8459 specparam_declaration_instance8459();
    specparam_declaration8460 specparam_declaration_instance8460();
    specparam_declaration8461 specparam_declaration_instance8461();
    specparam_declaration8462 specparam_declaration_instance8462();
    specparam_declaration8463 specparam_declaration_instance8463();
    specparam_declaration8464 specparam_declaration_instance8464();
    specparam_declaration8465 specparam_declaration_instance8465();
    specparam_declaration8466 specparam_declaration_instance8466();
    specparam_declaration8467 specparam_declaration_instance8467();
    specparam_declaration8468 specparam_declaration_instance8468();
    specparam_declaration8469 specparam_declaration_instance8469();
    specparam_declaration8470 specparam_declaration_instance8470();
    specparam_declaration8471 specparam_declaration_instance8471();
    specparam_declaration8472 specparam_declaration_instance8472();
    specparam_declaration8473 specparam_declaration_instance8473();
    specparam_declaration8474 specparam_declaration_instance8474();
    specparam_declaration8475 specparam_declaration_instance8475();
    specparam_declaration8476 specparam_declaration_instance8476();
    specparam_declaration8477 specparam_declaration_instance8477();
    specparam_declaration8478 specparam_declaration_instance8478();
    specparam_declaration8479 specparam_declaration_instance8479();
    specparam_declaration8480 specparam_declaration_instance8480();
    specparam_declaration8481 specparam_declaration_instance8481();
    specparam_declaration8482 specparam_declaration_instance8482();
    specparam_declaration8483 specparam_declaration_instance8483();
    specparam_declaration8484 specparam_declaration_instance8484();
    specparam_declaration8485 specparam_declaration_instance8485();
    specparam_declaration8486 specparam_declaration_instance8486();
    specparam_declaration8487 specparam_declaration_instance8487();
    specparam_declaration8488 specparam_declaration_instance8488();
    specparam_declaration8489 specparam_declaration_instance8489();
    specparam_declaration8490 specparam_declaration_instance8490();
    specparam_declaration8491 specparam_declaration_instance8491();
    specparam_declaration8492 specparam_declaration_instance8492();
    specparam_declaration8493 specparam_declaration_instance8493();
    specparam_declaration8494 specparam_declaration_instance8494();
    specparam_declaration8495 specparam_declaration_instance8495();
    specparam_declaration8496 specparam_declaration_instance8496();
    specparam_declaration8497 specparam_declaration_instance8497();
    specparam_declaration8498 specparam_declaration_instance8498();
    specparam_declaration8499 specparam_declaration_instance8499();
    specparam_declaration8500 specparam_declaration_instance8500();
    specparam_declaration8501 specparam_declaration_instance8501();
    specparam_declaration8502 specparam_declaration_instance8502();
    specparam_declaration8503 specparam_declaration_instance8503();
    specparam_declaration8504 specparam_declaration_instance8504();
    specparam_declaration8505 specparam_declaration_instance8505();
    specparam_declaration8506 specparam_declaration_instance8506();
    specparam_declaration8507 specparam_declaration_instance8507();
    specparam_declaration8508 specparam_declaration_instance8508();
    specparam_declaration8509 specparam_declaration_instance8509();
    specparam_declaration8510 specparam_declaration_instance8510();
    specparam_declaration8511 specparam_declaration_instance8511();
    specparam_declaration8512 specparam_declaration_instance8512();
    specparam_declaration8513 specparam_declaration_instance8513();
    specparam_declaration8514 specparam_declaration_instance8514();
    specparam_declaration8515 specparam_declaration_instance8515();
    specparam_declaration8516 specparam_declaration_instance8516();
    specparam_declaration8517 specparam_declaration_instance8517();
    specparam_declaration8518 specparam_declaration_instance8518();
    specparam_declaration8519 specparam_declaration_instance8519();
    specparam_declaration8520 specparam_declaration_instance8520();
    specparam_declaration8521 specparam_declaration_instance8521();
    specparam_declaration8522 specparam_declaration_instance8522();
    specparam_declaration8523 specparam_declaration_instance8523();
    specparam_declaration8524 specparam_declaration_instance8524();
    specparam_declaration8525 specparam_declaration_instance8525();
    specparam_declaration8526 specparam_declaration_instance8526();
    specparam_declaration8527 specparam_declaration_instance8527();
    specparam_declaration8528 specparam_declaration_instance8528();
    specparam_declaration8529 specparam_declaration_instance8529();
    specparam_declaration8530 specparam_declaration_instance8530();
    specparam_declaration8531 specparam_declaration_instance8531();
    specparam_declaration8532 specparam_declaration_instance8532();
    specparam_declaration8533 specparam_declaration_instance8533();
    specparam_declaration8534 specparam_declaration_instance8534();
    specparam_declaration8535 specparam_declaration_instance8535();
    specparam_declaration8536 specparam_declaration_instance8536();
    specparam_declaration8537 specparam_declaration_instance8537();
    specparam_declaration8538 specparam_declaration_instance8538();
    specparam_declaration8539 specparam_declaration_instance8539();
    specparam_declaration8540 specparam_declaration_instance8540();
    specparam_declaration8541 specparam_declaration_instance8541();
    specparam_declaration8542 specparam_declaration_instance8542();
    specparam_declaration8543 specparam_declaration_instance8543();
    specparam_declaration8544 specparam_declaration_instance8544();
    specparam_declaration8545 specparam_declaration_instance8545();
    specparam_declaration8546 specparam_declaration_instance8546();
    specparam_declaration8547 specparam_declaration_instance8547();
    specparam_declaration8548 specparam_declaration_instance8548();
    specparam_declaration8549 specparam_declaration_instance8549();
    specparam_declaration8550 specparam_declaration_instance8550();
    specparam_declaration8551 specparam_declaration_instance8551();
    specparam_declaration8552 specparam_declaration_instance8552();
    specparam_declaration8553 specparam_declaration_instance8553();
    specparam_declaration8554 specparam_declaration_instance8554();
    specparam_declaration8555 specparam_declaration_instance8555();
    specparam_declaration8556 specparam_declaration_instance8556();
    specparam_declaration8557 specparam_declaration_instance8557();
    specparam_declaration8558 specparam_declaration_instance8558();
    specparam_declaration8559 specparam_declaration_instance8559();
    specparam_declaration8560 specparam_declaration_instance8560();
    specparam_declaration8561 specparam_declaration_instance8561();
    specparam_declaration8562 specparam_declaration_instance8562();
    specparam_declaration8563 specparam_declaration_instance8563();
    specparam_declaration8564 specparam_declaration_instance8564();
    specparam_declaration8565 specparam_declaration_instance8565();
    specparam_declaration8566 specparam_declaration_instance8566();
    specparam_declaration8567 specparam_declaration_instance8567();
    specparam_declaration8568 specparam_declaration_instance8568();
    specparam_declaration8569 specparam_declaration_instance8569();
    specparam_declaration8570 specparam_declaration_instance8570();
    specparam_declaration8571 specparam_declaration_instance8571();
    specparam_declaration8572 specparam_declaration_instance8572();
    specparam_declaration8573 specparam_declaration_instance8573();
    specparam_declaration8574 specparam_declaration_instance8574();
    specparam_declaration8575 specparam_declaration_instance8575();
    specparam_declaration8576 specparam_declaration_instance8576();
    specparam_declaration8577 specparam_declaration_instance8577();
    specparam_declaration8578 specparam_declaration_instance8578();
    specparam_declaration8579 specparam_declaration_instance8579();
    specparam_declaration8580 specparam_declaration_instance8580();
    specparam_declaration8581 specparam_declaration_instance8581();
    specparam_declaration8582 specparam_declaration_instance8582();
    specparam_declaration8583 specparam_declaration_instance8583();
    specparam_declaration8584 specparam_declaration_instance8584();
    specparam_declaration8585 specparam_declaration_instance8585();
    specparam_declaration8586 specparam_declaration_instance8586();
    specparam_declaration8587 specparam_declaration_instance8587();
    specparam_declaration8588 specparam_declaration_instance8588();
    specparam_declaration8589 specparam_declaration_instance8589();
    specparam_declaration8590 specparam_declaration_instance8590();
    specparam_declaration8591 specparam_declaration_instance8591();
    specparam_declaration8592 specparam_declaration_instance8592();
    specparam_declaration8593 specparam_declaration_instance8593();
    specparam_declaration8594 specparam_declaration_instance8594();
    specparam_declaration8595 specparam_declaration_instance8595();
    specparam_declaration8596 specparam_declaration_instance8596();
    specparam_declaration8597 specparam_declaration_instance8597();
    specparam_declaration8598 specparam_declaration_instance8598();
    specparam_declaration8599 specparam_declaration_instance8599();
    specparam_declaration8600 specparam_declaration_instance8600();
    specparam_declaration8601 specparam_declaration_instance8601();
    specparam_declaration8602 specparam_declaration_instance8602();
    specparam_declaration8603 specparam_declaration_instance8603();
    specparam_declaration8604 specparam_declaration_instance8604();
    specparam_declaration8605 specparam_declaration_instance8605();
    specparam_declaration8606 specparam_declaration_instance8606();
    specparam_declaration8607 specparam_declaration_instance8607();
    specparam_declaration8608 specparam_declaration_instance8608();
    specparam_declaration8609 specparam_declaration_instance8609();
    specparam_declaration8610 specparam_declaration_instance8610();
    specparam_declaration8611 specparam_declaration_instance8611();
    specparam_declaration8612 specparam_declaration_instance8612();
    specparam_declaration8613 specparam_declaration_instance8613();
    specparam_declaration8614 specparam_declaration_instance8614();
    specparam_declaration8615 specparam_declaration_instance8615();
    specparam_declaration8616 specparam_declaration_instance8616();
    specparam_declaration8617 specparam_declaration_instance8617();
    specparam_declaration8618 specparam_declaration_instance8618();
    specparam_declaration8619 specparam_declaration_instance8619();
    specparam_declaration8620 specparam_declaration_instance8620();
    specparam_declaration8621 specparam_declaration_instance8621();
    specparam_declaration8622 specparam_declaration_instance8622();
    specparam_declaration8623 specparam_declaration_instance8623();
    specparam_declaration8624 specparam_declaration_instance8624();
    specparam_declaration8625 specparam_declaration_instance8625();
    specparam_declaration8626 specparam_declaration_instance8626();
    specparam_declaration8627 specparam_declaration_instance8627();
    specparam_declaration8628 specparam_declaration_instance8628();
    specparam_declaration8629 specparam_declaration_instance8629();
    specparam_declaration8630 specparam_declaration_instance8630();
    specparam_declaration8631 specparam_declaration_instance8631();
    specparam_declaration8632 specparam_declaration_instance8632();
    specparam_declaration8633 specparam_declaration_instance8633();
    specparam_declaration8634 specparam_declaration_instance8634();
    specparam_declaration8635 specparam_declaration_instance8635();
    specparam_declaration8636 specparam_declaration_instance8636();
    specparam_declaration8637 specparam_declaration_instance8637();
    specparam_declaration8638 specparam_declaration_instance8638();
    specparam_declaration8639 specparam_declaration_instance8639();
    specparam_declaration8640 specparam_declaration_instance8640();
    specparam_declaration8641 specparam_declaration_instance8641();
    specparam_declaration8642 specparam_declaration_instance8642();
    specparam_declaration8643 specparam_declaration_instance8643();
    specparam_declaration8644 specparam_declaration_instance8644();
    specparam_declaration8645 specparam_declaration_instance8645();
    specparam_declaration8646 specparam_declaration_instance8646();
    specparam_declaration8647 specparam_declaration_instance8647();
    specparam_declaration8648 specparam_declaration_instance8648();
    specparam_declaration8649 specparam_declaration_instance8649();
    specparam_declaration8650 specparam_declaration_instance8650();
    specparam_declaration8651 specparam_declaration_instance8651();
    specparam_declaration8652 specparam_declaration_instance8652();
    specparam_declaration8653 specparam_declaration_instance8653();
    specparam_declaration8654 specparam_declaration_instance8654();
    specparam_declaration8655 specparam_declaration_instance8655();
    specparam_declaration8656 specparam_declaration_instance8656();
    specparam_declaration8657 specparam_declaration_instance8657();
    specparam_declaration8658 specparam_declaration_instance8658();
    specparam_declaration8659 specparam_declaration_instance8659();
    specparam_declaration8660 specparam_declaration_instance8660();
    specparam_declaration8661 specparam_declaration_instance8661();
    specparam_declaration8662 specparam_declaration_instance8662();
    specparam_declaration8663 specparam_declaration_instance8663();
    specparam_declaration8664 specparam_declaration_instance8664();
    specparam_declaration8665 specparam_declaration_instance8665();
    specparam_declaration8666 specparam_declaration_instance8666();
    specparam_declaration8667 specparam_declaration_instance8667();
    specparam_declaration8668 specparam_declaration_instance8668();
    specparam_declaration8669 specparam_declaration_instance8669();
    specparam_declaration8670 specparam_declaration_instance8670();
    specparam_declaration8671 specparam_declaration_instance8671();
    specparam_declaration8672 specparam_declaration_instance8672();
    specparam_declaration8673 specparam_declaration_instance8673();
    specparam_declaration8674 specparam_declaration_instance8674();
    specparam_declaration8675 specparam_declaration_instance8675();
    specparam_declaration8676 specparam_declaration_instance8676();
    specparam_declaration8677 specparam_declaration_instance8677();
    specparam_declaration8678 specparam_declaration_instance8678();
    specparam_declaration8679 specparam_declaration_instance8679();
    specparam_declaration8680 specparam_declaration_instance8680();
    specparam_declaration8681 specparam_declaration_instance8681();
    specparam_declaration8682 specparam_declaration_instance8682();
    specparam_declaration8683 specparam_declaration_instance8683();
    specparam_declaration8684 specparam_declaration_instance8684();
    specparam_declaration8685 specparam_declaration_instance8685();
    specparam_declaration8686 specparam_declaration_instance8686();
    specparam_declaration8687 specparam_declaration_instance8687();
    specparam_declaration8688 specparam_declaration_instance8688();
    specparam_declaration8689 specparam_declaration_instance8689();
    specparam_declaration8690 specparam_declaration_instance8690();
    specparam_declaration8691 specparam_declaration_instance8691();
    specparam_declaration8692 specparam_declaration_instance8692();
    specparam_declaration8693 specparam_declaration_instance8693();
    specparam_declaration8694 specparam_declaration_instance8694();
    specparam_declaration8695 specparam_declaration_instance8695();
    specparam_declaration8696 specparam_declaration_instance8696();
    specparam_declaration8697 specparam_declaration_instance8697();
    specparam_declaration8698 specparam_declaration_instance8698();
    specparam_declaration8699 specparam_declaration_instance8699();
    specparam_declaration8700 specparam_declaration_instance8700();
    specparam_declaration8701 specparam_declaration_instance8701();
    specparam_declaration8702 specparam_declaration_instance8702();
    specparam_declaration8703 specparam_declaration_instance8703();
    specparam_declaration8704 specparam_declaration_instance8704();
    specparam_declaration8705 specparam_declaration_instance8705();
    specparam_declaration8706 specparam_declaration_instance8706();
    specparam_declaration8707 specparam_declaration_instance8707();
    specparam_declaration8708 specparam_declaration_instance8708();
    specparam_declaration8709 specparam_declaration_instance8709();
    specparam_declaration8710 specparam_declaration_instance8710();
    specparam_declaration8711 specparam_declaration_instance8711();
    specparam_declaration8712 specparam_declaration_instance8712();
    specparam_declaration8713 specparam_declaration_instance8713();
    specparam_declaration8714 specparam_declaration_instance8714();
    specparam_declaration8715 specparam_declaration_instance8715();
    specparam_declaration8716 specparam_declaration_instance8716();
    specparam_declaration8717 specparam_declaration_instance8717();
    specparam_declaration8718 specparam_declaration_instance8718();
    specparam_declaration8719 specparam_declaration_instance8719();
    specparam_declaration8720 specparam_declaration_instance8720();
    specparam_declaration8721 specparam_declaration_instance8721();
    specparam_declaration8722 specparam_declaration_instance8722();
    specparam_declaration8723 specparam_declaration_instance8723();
    specparam_declaration8724 specparam_declaration_instance8724();
    specparam_declaration8725 specparam_declaration_instance8725();
    specparam_declaration8726 specparam_declaration_instance8726();
    specparam_declaration8727 specparam_declaration_instance8727();
    specparam_declaration8728 specparam_declaration_instance8728();
    specparam_declaration8729 specparam_declaration_instance8729();
    specparam_declaration8730 specparam_declaration_instance8730();
    specparam_declaration8731 specparam_declaration_instance8731();
    specparam_declaration8732 specparam_declaration_instance8732();
    specparam_declaration8733 specparam_declaration_instance8733();
    specparam_declaration8734 specparam_declaration_instance8734();
    specparam_declaration8735 specparam_declaration_instance8735();
    specparam_declaration8736 specparam_declaration_instance8736();
    specparam_declaration8737 specparam_declaration_instance8737();
    specparam_declaration8738 specparam_declaration_instance8738();
    specparam_declaration8739 specparam_declaration_instance8739();
    specparam_declaration8740 specparam_declaration_instance8740();
    specparam_declaration8741 specparam_declaration_instance8741();
    specparam_declaration8742 specparam_declaration_instance8742();
    specparam_declaration8743 specparam_declaration_instance8743();
    specparam_declaration8744 specparam_declaration_instance8744();
    specparam_declaration8745 specparam_declaration_instance8745();
    specparam_declaration8746 specparam_declaration_instance8746();
    specparam_declaration8747 specparam_declaration_instance8747();
    specparam_declaration8748 specparam_declaration_instance8748();
    specparam_declaration8749 specparam_declaration_instance8749();
    specparam_declaration8750 specparam_declaration_instance8750();
    specparam_declaration8751 specparam_declaration_instance8751();
    specparam_declaration8752 specparam_declaration_instance8752();
    specparam_declaration8753 specparam_declaration_instance8753();
    specparam_declaration8754 specparam_declaration_instance8754();
    specparam_declaration8755 specparam_declaration_instance8755();
    specparam_declaration8756 specparam_declaration_instance8756();
    specparam_declaration8757 specparam_declaration_instance8757();
    specparam_declaration8758 specparam_declaration_instance8758();
    specparam_declaration8759 specparam_declaration_instance8759();
    specparam_declaration8760 specparam_declaration_instance8760();
    specparam_declaration8761 specparam_declaration_instance8761();
    specparam_declaration8762 specparam_declaration_instance8762();
    specparam_declaration8763 specparam_declaration_instance8763();
    specparam_declaration8764 specparam_declaration_instance8764();
    specparam_declaration8765 specparam_declaration_instance8765();
    specparam_declaration8766 specparam_declaration_instance8766();
    specparam_declaration8767 specparam_declaration_instance8767();
    specparam_declaration8768 specparam_declaration_instance8768();
    specparam_declaration8769 specparam_declaration_instance8769();
    specparam_declaration8770 specparam_declaration_instance8770();
    specparam_declaration8771 specparam_declaration_instance8771();
    specparam_declaration8772 specparam_declaration_instance8772();
    specparam_declaration8773 specparam_declaration_instance8773();
    specparam_declaration8774 specparam_declaration_instance8774();
    specparam_declaration8775 specparam_declaration_instance8775();
    specparam_declaration8776 specparam_declaration_instance8776();
    specparam_declaration8777 specparam_declaration_instance8777();
    specparam_declaration8778 specparam_declaration_instance8778();
    specparam_declaration8779 specparam_declaration_instance8779();
    specparam_declaration8780 specparam_declaration_instance8780();
    specparam_declaration8781 specparam_declaration_instance8781();
    specparam_declaration8782 specparam_declaration_instance8782();
    specparam_declaration8783 specparam_declaration_instance8783();
    specparam_declaration8784 specparam_declaration_instance8784();
    specparam_declaration8785 specparam_declaration_instance8785();
    specparam_declaration8786 specparam_declaration_instance8786();
    specparam_declaration8787 specparam_declaration_instance8787();
    specparam_declaration8788 specparam_declaration_instance8788();
    specparam_declaration8789 specparam_declaration_instance8789();
    specparam_declaration8790 specparam_declaration_instance8790();
    specparam_declaration8791 specparam_declaration_instance8791();
    specparam_declaration8792 specparam_declaration_instance8792();
    specparam_declaration8793 specparam_declaration_instance8793();
    specparam_declaration8794 specparam_declaration_instance8794();
    specparam_declaration8795 specparam_declaration_instance8795();
    specparam_declaration8796 specparam_declaration_instance8796();
    specparam_declaration8797 specparam_declaration_instance8797();
    specparam_declaration8798 specparam_declaration_instance8798();
    specparam_declaration8799 specparam_declaration_instance8799();
    specparam_declaration8800 specparam_declaration_instance8800();
    specparam_declaration8801 specparam_declaration_instance8801();
    specparam_declaration8802 specparam_declaration_instance8802();
    specparam_declaration8803 specparam_declaration_instance8803();
    specparam_declaration8804 specparam_declaration_instance8804();
    specparam_declaration8805 specparam_declaration_instance8805();
    specparam_declaration8806 specparam_declaration_instance8806();
    specparam_declaration8807 specparam_declaration_instance8807();
    specparam_declaration8808 specparam_declaration_instance8808();
    specparam_declaration8809 specparam_declaration_instance8809();
    specparam_declaration8810 specparam_declaration_instance8810();
    specparam_declaration8811 specparam_declaration_instance8811();
    specparam_declaration8812 specparam_declaration_instance8812();
    specparam_declaration8813 specparam_declaration_instance8813();
    specparam_declaration8814 specparam_declaration_instance8814();
    specparam_declaration8815 specparam_declaration_instance8815();
    specparam_declaration8816 specparam_declaration_instance8816();
    specparam_declaration8817 specparam_declaration_instance8817();
    specparam_declaration8818 specparam_declaration_instance8818();
    specparam_declaration8819 specparam_declaration_instance8819();
    specparam_declaration8820 specparam_declaration_instance8820();
    specparam_declaration8821 specparam_declaration_instance8821();
    specparam_declaration8822 specparam_declaration_instance8822();
    specparam_declaration8823 specparam_declaration_instance8823();
    specparam_declaration8824 specparam_declaration_instance8824();
    specparam_declaration8825 specparam_declaration_instance8825();
    specparam_declaration8826 specparam_declaration_instance8826();
    specparam_declaration8827 specparam_declaration_instance8827();
    specparam_declaration8828 specparam_declaration_instance8828();
    specparam_declaration8829 specparam_declaration_instance8829();
    specparam_declaration8830 specparam_declaration_instance8830();
    specparam_declaration8831 specparam_declaration_instance8831();
    specparam_declaration8832 specparam_declaration_instance8832();
    specparam_declaration8833 specparam_declaration_instance8833();
    specparam_declaration8834 specparam_declaration_instance8834();
    specparam_declaration8835 specparam_declaration_instance8835();
    specparam_declaration8836 specparam_declaration_instance8836();
    specparam_declaration8837 specparam_declaration_instance8837();
    specparam_declaration8838 specparam_declaration_instance8838();
    specparam_declaration8839 specparam_declaration_instance8839();
    specparam_declaration8840 specparam_declaration_instance8840();
    specparam_declaration8841 specparam_declaration_instance8841();
    specparam_declaration8842 specparam_declaration_instance8842();
    specparam_declaration8843 specparam_declaration_instance8843();
    specparam_declaration8844 specparam_declaration_instance8844();
    specparam_declaration8845 specparam_declaration_instance8845();
    specparam_declaration8846 specparam_declaration_instance8846();
    specparam_declaration8847 specparam_declaration_instance8847();
    specparam_declaration8848 specparam_declaration_instance8848();
    specparam_declaration8849 specparam_declaration_instance8849();
    specparam_declaration8850 specparam_declaration_instance8850();
    specparam_declaration8851 specparam_declaration_instance8851();
    specparam_declaration8852 specparam_declaration_instance8852();
    specparam_declaration8853 specparam_declaration_instance8853();
    specparam_declaration8854 specparam_declaration_instance8854();
    specparam_declaration8855 specparam_declaration_instance8855();
    specparam_declaration8856 specparam_declaration_instance8856();
    specparam_declaration8857 specparam_declaration_instance8857();
    specparam_declaration8858 specparam_declaration_instance8858();
    specparam_declaration8859 specparam_declaration_instance8859();
    specparam_declaration8860 specparam_declaration_instance8860();
    specparam_declaration8861 specparam_declaration_instance8861();
    specparam_declaration8862 specparam_declaration_instance8862();
    specparam_declaration8863 specparam_declaration_instance8863();
    specparam_declaration8864 specparam_declaration_instance8864();
    specparam_declaration8865 specparam_declaration_instance8865();
    specparam_declaration8866 specparam_declaration_instance8866();
    specparam_declaration8867 specparam_declaration_instance8867();
    specparam_declaration8868 specparam_declaration_instance8868();
    specparam_declaration8869 specparam_declaration_instance8869();
    specparam_declaration8870 specparam_declaration_instance8870();
    specparam_declaration8871 specparam_declaration_instance8871();
    specparam_declaration8872 specparam_declaration_instance8872();
    specparam_declaration8873 specparam_declaration_instance8873();
    specparam_declaration8874 specparam_declaration_instance8874();
    specparam_declaration8875 specparam_declaration_instance8875();
    specparam_declaration8876 specparam_declaration_instance8876();
    specparam_declaration8877 specparam_declaration_instance8877();
    specparam_declaration8878 specparam_declaration_instance8878();
    specparam_declaration8879 specparam_declaration_instance8879();
    specparam_declaration8880 specparam_declaration_instance8880();
    specparam_declaration8881 specparam_declaration_instance8881();
    specparam_declaration8882 specparam_declaration_instance8882();
    specparam_declaration8883 specparam_declaration_instance8883();
    specparam_declaration8884 specparam_declaration_instance8884();
    specparam_declaration8885 specparam_declaration_instance8885();
    specparam_declaration8886 specparam_declaration_instance8886();
    specparam_declaration8887 specparam_declaration_instance8887();
    specparam_declaration8888 specparam_declaration_instance8888();
    specparam_declaration8889 specparam_declaration_instance8889();
    specparam_declaration8890 specparam_declaration_instance8890();
    specparam_declaration8891 specparam_declaration_instance8891();
    specparam_declaration8892 specparam_declaration_instance8892();
    specparam_declaration8893 specparam_declaration_instance8893();
    specparam_declaration8894 specparam_declaration_instance8894();
    specparam_declaration8895 specparam_declaration_instance8895();
    specparam_declaration8896 specparam_declaration_instance8896();
    specparam_declaration8897 specparam_declaration_instance8897();
    specparam_declaration8898 specparam_declaration_instance8898();
    specparam_declaration8899 specparam_declaration_instance8899();
    specparam_declaration8900 specparam_declaration_instance8900();
    specparam_declaration8901 specparam_declaration_instance8901();
    specparam_declaration8902 specparam_declaration_instance8902();
    specparam_declaration8903 specparam_declaration_instance8903();
    specparam_declaration8904 specparam_declaration_instance8904();
    specparam_declaration8905 specparam_declaration_instance8905();
    specparam_declaration8906 specparam_declaration_instance8906();
    specparam_declaration8907 specparam_declaration_instance8907();
    specparam_declaration8908 specparam_declaration_instance8908();
    specparam_declaration8909 specparam_declaration_instance8909();
    specparam_declaration8910 specparam_declaration_instance8910();
    specparam_declaration8911 specparam_declaration_instance8911();
    specparam_declaration8912 specparam_declaration_instance8912();
    specparam_declaration8913 specparam_declaration_instance8913();
    specparam_declaration8914 specparam_declaration_instance8914();
    specparam_declaration8915 specparam_declaration_instance8915();
    specparam_declaration8916 specparam_declaration_instance8916();
    specparam_declaration8917 specparam_declaration_instance8917();
    specparam_declaration8918 specparam_declaration_instance8918();
    specparam_declaration8919 specparam_declaration_instance8919();
    specparam_declaration8920 specparam_declaration_instance8920();
    specparam_declaration8921 specparam_declaration_instance8921();
    specparam_declaration8922 specparam_declaration_instance8922();
    specparam_declaration8923 specparam_declaration_instance8923();
    specparam_declaration8924 specparam_declaration_instance8924();
    specparam_declaration8925 specparam_declaration_instance8925();
    specparam_declaration8926 specparam_declaration_instance8926();
    specparam_declaration8927 specparam_declaration_instance8927();
    specparam_declaration8928 specparam_declaration_instance8928();
    specparam_declaration8929 specparam_declaration_instance8929();
    specparam_declaration8930 specparam_declaration_instance8930();
    specparam_declaration8931 specparam_declaration_instance8931();
    specparam_declaration8932 specparam_declaration_instance8932();
    specparam_declaration8933 specparam_declaration_instance8933();
    specparam_declaration8934 specparam_declaration_instance8934();
    specparam_declaration8935 specparam_declaration_instance8935();
    specparam_declaration8936 specparam_declaration_instance8936();
    specparam_declaration8937 specparam_declaration_instance8937();
    specparam_declaration8938 specparam_declaration_instance8938();
    specparam_declaration8939 specparam_declaration_instance8939();
    specparam_declaration8940 specparam_declaration_instance8940();
    specparam_declaration8941 specparam_declaration_instance8941();
    specparam_declaration8942 specparam_declaration_instance8942();
    specparam_declaration8943 specparam_declaration_instance8943();
    specparam_declaration8944 specparam_declaration_instance8944();
    specparam_declaration8945 specparam_declaration_instance8945();
    specparam_declaration8946 specparam_declaration_instance8946();
    specparam_declaration8947 specparam_declaration_instance8947();
    specparam_declaration8948 specparam_declaration_instance8948();
    specparam_declaration8949 specparam_declaration_instance8949();
    specparam_declaration8950 specparam_declaration_instance8950();
    specparam_declaration8951 specparam_declaration_instance8951();
    specparam_declaration8952 specparam_declaration_instance8952();
    specparam_declaration8953 specparam_declaration_instance8953();
    specparam_declaration8954 specparam_declaration_instance8954();
    specparam_declaration8955 specparam_declaration_instance8955();
    specparam_declaration8956 specparam_declaration_instance8956();
    specparam_declaration8957 specparam_declaration_instance8957();
    specparam_declaration8958 specparam_declaration_instance8958();
    specparam_declaration8959 specparam_declaration_instance8959();
    specparam_declaration8960 specparam_declaration_instance8960();
    specparam_declaration8961 specparam_declaration_instance8961();
    specparam_declaration8962 specparam_declaration_instance8962();
    specparam_declaration8963 specparam_declaration_instance8963();
    specparam_declaration8964 specparam_declaration_instance8964();
    specparam_declaration8965 specparam_declaration_instance8965();
    specparam_declaration8966 specparam_declaration_instance8966();
    specparam_declaration8967 specparam_declaration_instance8967();
    specparam_declaration8968 specparam_declaration_instance8968();
    specparam_declaration8969 specparam_declaration_instance8969();
    specparam_declaration8970 specparam_declaration_instance8970();
    specparam_declaration8971 specparam_declaration_instance8971();
    specparam_declaration8972 specparam_declaration_instance8972();
    specparam_declaration8973 specparam_declaration_instance8973();
    specparam_declaration8974 specparam_declaration_instance8974();
    specparam_declaration8975 specparam_declaration_instance8975();
    specparam_declaration8976 specparam_declaration_instance8976();
    specparam_declaration8977 specparam_declaration_instance8977();
    specparam_declaration8978 specparam_declaration_instance8978();
    specparam_declaration8979 specparam_declaration_instance8979();
    specparam_declaration8980 specparam_declaration_instance8980();
    specparam_declaration8981 specparam_declaration_instance8981();
    specparam_declaration8982 specparam_declaration_instance8982();
    specparam_declaration8983 specparam_declaration_instance8983();
    specparam_declaration8984 specparam_declaration_instance8984();
    specparam_declaration8985 specparam_declaration_instance8985();
    specparam_declaration8986 specparam_declaration_instance8986();
    specparam_declaration8987 specparam_declaration_instance8987();
    specparam_declaration8988 specparam_declaration_instance8988();
    specparam_declaration8989 specparam_declaration_instance8989();
    specparam_declaration8990 specparam_declaration_instance8990();
    specparam_declaration8991 specparam_declaration_instance8991();
    specparam_declaration8992 specparam_declaration_instance8992();
    specparam_declaration8993 specparam_declaration_instance8993();
    specparam_declaration8994 specparam_declaration_instance8994();
    specparam_declaration8995 specparam_declaration_instance8995();
    specparam_declaration8996 specparam_declaration_instance8996();
    specparam_declaration8997 specparam_declaration_instance8997();
    specparam_declaration8998 specparam_declaration_instance8998();
    specparam_declaration8999 specparam_declaration_instance8999();
    specparam_declaration9000 specparam_declaration_instance9000();
    specparam_declaration9001 specparam_declaration_instance9001();
    specparam_declaration9002 specparam_declaration_instance9002();
    specparam_declaration9003 specparam_declaration_instance9003();
    specparam_declaration9004 specparam_declaration_instance9004();
    specparam_declaration9005 specparam_declaration_instance9005();
    specparam_declaration9006 specparam_declaration_instance9006();
    specparam_declaration9007 specparam_declaration_instance9007();
    specparam_declaration9008 specparam_declaration_instance9008();
    specparam_declaration9009 specparam_declaration_instance9009();
    specparam_declaration9010 specparam_declaration_instance9010();
    specparam_declaration9011 specparam_declaration_instance9011();
    specparam_declaration9012 specparam_declaration_instance9012();
    specparam_declaration9013 specparam_declaration_instance9013();
    specparam_declaration9014 specparam_declaration_instance9014();
    specparam_declaration9015 specparam_declaration_instance9015();
    specparam_declaration9016 specparam_declaration_instance9016();
    specparam_declaration9017 specparam_declaration_instance9017();
    specparam_declaration9018 specparam_declaration_instance9018();
    specparam_declaration9019 specparam_declaration_instance9019();
    specparam_declaration9020 specparam_declaration_instance9020();
    specparam_declaration9021 specparam_declaration_instance9021();
    specparam_declaration9022 specparam_declaration_instance9022();
    specparam_declaration9023 specparam_declaration_instance9023();
    specparam_declaration9024 specparam_declaration_instance9024();
    specparam_declaration9025 specparam_declaration_instance9025();
    specparam_declaration9026 specparam_declaration_instance9026();
    specparam_declaration9027 specparam_declaration_instance9027();
    specparam_declaration9028 specparam_declaration_instance9028();
    specparam_declaration9029 specparam_declaration_instance9029();
    specparam_declaration9030 specparam_declaration_instance9030();
    specparam_declaration9031 specparam_declaration_instance9031();
    specparam_declaration9032 specparam_declaration_instance9032();
    specparam_declaration9033 specparam_declaration_instance9033();
    specparam_declaration9034 specparam_declaration_instance9034();
    specparam_declaration9035 specparam_declaration_instance9035();
    specparam_declaration9036 specparam_declaration_instance9036();
    specparam_declaration9037 specparam_declaration_instance9037();
    specparam_declaration9038 specparam_declaration_instance9038();
    specparam_declaration9039 specparam_declaration_instance9039();
    specparam_declaration9040 specparam_declaration_instance9040();
    specparam_declaration9041 specparam_declaration_instance9041();
    specparam_declaration9042 specparam_declaration_instance9042();
    specparam_declaration9043 specparam_declaration_instance9043();
    specparam_declaration9044 specparam_declaration_instance9044();
    specparam_declaration9045 specparam_declaration_instance9045();
    specparam_declaration9046 specparam_declaration_instance9046();
    specparam_declaration9047 specparam_declaration_instance9047();
    specparam_declaration9048 specparam_declaration_instance9048();
    specparam_declaration9049 specparam_declaration_instance9049();
    specparam_declaration9050 specparam_declaration_instance9050();
    specparam_declaration9051 specparam_declaration_instance9051();
    specparam_declaration9052 specparam_declaration_instance9052();
    specparam_declaration9053 specparam_declaration_instance9053();
    specparam_declaration9054 specparam_declaration_instance9054();
    specparam_declaration9055 specparam_declaration_instance9055();
    specparam_declaration9056 specparam_declaration_instance9056();
    specparam_declaration9057 specparam_declaration_instance9057();
    specparam_declaration9058 specparam_declaration_instance9058();
    specparam_declaration9059 specparam_declaration_instance9059();
    specparam_declaration9060 specparam_declaration_instance9060();
    specparam_declaration9061 specparam_declaration_instance9061();
    specparam_declaration9062 specparam_declaration_instance9062();
    specparam_declaration9063 specparam_declaration_instance9063();
    specparam_declaration9064 specparam_declaration_instance9064();
    specparam_declaration9065 specparam_declaration_instance9065();
    specparam_declaration9066 specparam_declaration_instance9066();
    specparam_declaration9067 specparam_declaration_instance9067();
    specparam_declaration9068 specparam_declaration_instance9068();
    specparam_declaration9069 specparam_declaration_instance9069();
    specparam_declaration9070 specparam_declaration_instance9070();
    specparam_declaration9071 specparam_declaration_instance9071();
    specparam_declaration9072 specparam_declaration_instance9072();
    specparam_declaration9073 specparam_declaration_instance9073();
    specparam_declaration9074 specparam_declaration_instance9074();
    specparam_declaration9075 specparam_declaration_instance9075();
    specparam_declaration9076 specparam_declaration_instance9076();
    specparam_declaration9077 specparam_declaration_instance9077();
    specparam_declaration9078 specparam_declaration_instance9078();
    specparam_declaration9079 specparam_declaration_instance9079();
    specparam_declaration9080 specparam_declaration_instance9080();
    specparam_declaration9081 specparam_declaration_instance9081();
    specparam_declaration9082 specparam_declaration_instance9082();
    specparam_declaration9083 specparam_declaration_instance9083();
    specparam_declaration9084 specparam_declaration_instance9084();
    specparam_declaration9085 specparam_declaration_instance9085();
    specparam_declaration9086 specparam_declaration_instance9086();
    specparam_declaration9087 specparam_declaration_instance9087();
    specparam_declaration9088 specparam_declaration_instance9088();
    specparam_declaration9089 specparam_declaration_instance9089();
    specparam_declaration9090 specparam_declaration_instance9090();
    specparam_declaration9091 specparam_declaration_instance9091();
    specparam_declaration9092 specparam_declaration_instance9092();
    specparam_declaration9093 specparam_declaration_instance9093();
    specparam_declaration9094 specparam_declaration_instance9094();
    specparam_declaration9095 specparam_declaration_instance9095();
    specparam_declaration9096 specparam_declaration_instance9096();
    specparam_declaration9097 specparam_declaration_instance9097();
    specparam_declaration9098 specparam_declaration_instance9098();
    specparam_declaration9099 specparam_declaration_instance9099();
    specparam_declaration9100 specparam_declaration_instance9100();
    specparam_declaration9101 specparam_declaration_instance9101();
    specparam_declaration9102 specparam_declaration_instance9102();
    specparam_declaration9103 specparam_declaration_instance9103();
    specparam_declaration9104 specparam_declaration_instance9104();
    specparam_declaration9105 specparam_declaration_instance9105();
    specparam_declaration9106 specparam_declaration_instance9106();
    specparam_declaration9107 specparam_declaration_instance9107();
    specparam_declaration9108 specparam_declaration_instance9108();
    specparam_declaration9109 specparam_declaration_instance9109();
    specparam_declaration9110 specparam_declaration_instance9110();
    specparam_declaration9111 specparam_declaration_instance9111();
    specparam_declaration9112 specparam_declaration_instance9112();
    specparam_declaration9113 specparam_declaration_instance9113();
    specparam_declaration9114 specparam_declaration_instance9114();
    specparam_declaration9115 specparam_declaration_instance9115();
    specparam_declaration9116 specparam_declaration_instance9116();
    specparam_declaration9117 specparam_declaration_instance9117();
    specparam_declaration9118 specparam_declaration_instance9118();
    specparam_declaration9119 specparam_declaration_instance9119();
    specparam_declaration9120 specparam_declaration_instance9120();
    specparam_declaration9121 specparam_declaration_instance9121();
    specparam_declaration9122 specparam_declaration_instance9122();
    specparam_declaration9123 specparam_declaration_instance9123();
    specparam_declaration9124 specparam_declaration_instance9124();
    specparam_declaration9125 specparam_declaration_instance9125();
    specparam_declaration9126 specparam_declaration_instance9126();
    specparam_declaration9127 specparam_declaration_instance9127();
    specparam_declaration9128 specparam_declaration_instance9128();
    specparam_declaration9129 specparam_declaration_instance9129();
    specparam_declaration9130 specparam_declaration_instance9130();
    specparam_declaration9131 specparam_declaration_instance9131();
    specparam_declaration9132 specparam_declaration_instance9132();
    specparam_declaration9133 specparam_declaration_instance9133();
    specparam_declaration9134 specparam_declaration_instance9134();
    specparam_declaration9135 specparam_declaration_instance9135();
    specparam_declaration9136 specparam_declaration_instance9136();
    specparam_declaration9137 specparam_declaration_instance9137();
    specparam_declaration9138 specparam_declaration_instance9138();
    specparam_declaration9139 specparam_declaration_instance9139();
    specparam_declaration9140 specparam_declaration_instance9140();
    specparam_declaration9141 specparam_declaration_instance9141();
    specparam_declaration9142 specparam_declaration_instance9142();
    specparam_declaration9143 specparam_declaration_instance9143();
    specparam_declaration9144 specparam_declaration_instance9144();
    specparam_declaration9145 specparam_declaration_instance9145();
    specparam_declaration9146 specparam_declaration_instance9146();
    specparam_declaration9147 specparam_declaration_instance9147();
    specparam_declaration9148 specparam_declaration_instance9148();
    specparam_declaration9149 specparam_declaration_instance9149();
    specparam_declaration9150 specparam_declaration_instance9150();
    specparam_declaration9151 specparam_declaration_instance9151();
    specparam_declaration9152 specparam_declaration_instance9152();
    specparam_declaration9153 specparam_declaration_instance9153();
    specparam_declaration9154 specparam_declaration_instance9154();
    specparam_declaration9155 specparam_declaration_instance9155();
    specparam_declaration9156 specparam_declaration_instance9156();
    specparam_declaration9157 specparam_declaration_instance9157();
    specparam_declaration9158 specparam_declaration_instance9158();
    specparam_declaration9159 specparam_declaration_instance9159();
    specparam_declaration9160 specparam_declaration_instance9160();
    specparam_declaration9161 specparam_declaration_instance9161();
    specparam_declaration9162 specparam_declaration_instance9162();
    specparam_declaration9163 specparam_declaration_instance9163();
    specparam_declaration9164 specparam_declaration_instance9164();
    specparam_declaration9165 specparam_declaration_instance9165();
    specparam_declaration9166 specparam_declaration_instance9166();
    specparam_declaration9167 specparam_declaration_instance9167();
    specparam_declaration9168 specparam_declaration_instance9168();
    specparam_declaration9169 specparam_declaration_instance9169();
    specparam_declaration9170 specparam_declaration_instance9170();
    specparam_declaration9171 specparam_declaration_instance9171();
    specparam_declaration9172 specparam_declaration_instance9172();
    specparam_declaration9173 specparam_declaration_instance9173();
    specparam_declaration9174 specparam_declaration_instance9174();
    specparam_declaration9175 specparam_declaration_instance9175();
    specparam_declaration9176 specparam_declaration_instance9176();
    specparam_declaration9177 specparam_declaration_instance9177();
    specparam_declaration9178 specparam_declaration_instance9178();
    specparam_declaration9179 specparam_declaration_instance9179();
    specparam_declaration9180 specparam_declaration_instance9180();
    specparam_declaration9181 specparam_declaration_instance9181();
    specparam_declaration9182 specparam_declaration_instance9182();
    specparam_declaration9183 specparam_declaration_instance9183();
    specparam_declaration9184 specparam_declaration_instance9184();
    specparam_declaration9185 specparam_declaration_instance9185();
    specparam_declaration9186 specparam_declaration_instance9186();
    specparam_declaration9187 specparam_declaration_instance9187();
    specparam_declaration9188 specparam_declaration_instance9188();
    specparam_declaration9189 specparam_declaration_instance9189();
    specparam_declaration9190 specparam_declaration_instance9190();
    specparam_declaration9191 specparam_declaration_instance9191();
    specparam_declaration9192 specparam_declaration_instance9192();
    specparam_declaration9193 specparam_declaration_instance9193();
    specparam_declaration9194 specparam_declaration_instance9194();
    specparam_declaration9195 specparam_declaration_instance9195();
    specparam_declaration9196 specparam_declaration_instance9196();
    specparam_declaration9197 specparam_declaration_instance9197();
    specparam_declaration9198 specparam_declaration_instance9198();
    specparam_declaration9199 specparam_declaration_instance9199();
    specparam_declaration9200 specparam_declaration_instance9200();
    specparam_declaration9201 specparam_declaration_instance9201();
    specparam_declaration9202 specparam_declaration_instance9202();
    specparam_declaration9203 specparam_declaration_instance9203();
    specparam_declaration9204 specparam_declaration_instance9204();
    specparam_declaration9205 specparam_declaration_instance9205();
    specparam_declaration9206 specparam_declaration_instance9206();
    specparam_declaration9207 specparam_declaration_instance9207();
    specparam_declaration9208 specparam_declaration_instance9208();
    specparam_declaration9209 specparam_declaration_instance9209();
    specparam_declaration9210 specparam_declaration_instance9210();
    specparam_declaration9211 specparam_declaration_instance9211();
    specparam_declaration9212 specparam_declaration_instance9212();
    specparam_declaration9213 specparam_declaration_instance9213();
    specparam_declaration9214 specparam_declaration_instance9214();
    specparam_declaration9215 specparam_declaration_instance9215();
    specparam_declaration9216 specparam_declaration_instance9216();
    specparam_declaration9217 specparam_declaration_instance9217();
    specparam_declaration9218 specparam_declaration_instance9218();
    specparam_declaration9219 specparam_declaration_instance9219();
    specparam_declaration9220 specparam_declaration_instance9220();
    specparam_declaration9221 specparam_declaration_instance9221();
    specparam_declaration9222 specparam_declaration_instance9222();
    specparam_declaration9223 specparam_declaration_instance9223();
    specparam_declaration9224 specparam_declaration_instance9224();
    specparam_declaration9225 specparam_declaration_instance9225();
    specparam_declaration9226 specparam_declaration_instance9226();
    specparam_declaration9227 specparam_declaration_instance9227();
    specparam_declaration9228 specparam_declaration_instance9228();
    specparam_declaration9229 specparam_declaration_instance9229();
    specparam_declaration9230 specparam_declaration_instance9230();
    specparam_declaration9231 specparam_declaration_instance9231();
    specparam_declaration9232 specparam_declaration_instance9232();
    specparam_declaration9233 specparam_declaration_instance9233();
    specparam_declaration9234 specparam_declaration_instance9234();
    specparam_declaration9235 specparam_declaration_instance9235();
    specparam_declaration9236 specparam_declaration_instance9236();
    specparam_declaration9237 specparam_declaration_instance9237();
    specparam_declaration9238 specparam_declaration_instance9238();
    specparam_declaration9239 specparam_declaration_instance9239();
    specparam_declaration9240 specparam_declaration_instance9240();
    specparam_declaration9241 specparam_declaration_instance9241();
    specparam_declaration9242 specparam_declaration_instance9242();
    specparam_declaration9243 specparam_declaration_instance9243();
    specparam_declaration9244 specparam_declaration_instance9244();
    specparam_declaration9245 specparam_declaration_instance9245();
    specparam_declaration9246 specparam_declaration_instance9246();
    specparam_declaration9247 specparam_declaration_instance9247();
    specparam_declaration9248 specparam_declaration_instance9248();
    specparam_declaration9249 specparam_declaration_instance9249();
    specparam_declaration9250 specparam_declaration_instance9250();
    specparam_declaration9251 specparam_declaration_instance9251();
    specparam_declaration9252 specparam_declaration_instance9252();
    specparam_declaration9253 specparam_declaration_instance9253();
    specparam_declaration9254 specparam_declaration_instance9254();
    specparam_declaration9255 specparam_declaration_instance9255();
    specparam_declaration9256 specparam_declaration_instance9256();
    specparam_declaration9257 specparam_declaration_instance9257();
    specparam_declaration9258 specparam_declaration_instance9258();
    specparam_declaration9259 specparam_declaration_instance9259();
    specparam_declaration9260 specparam_declaration_instance9260();
    specparam_declaration9261 specparam_declaration_instance9261();
    specparam_declaration9262 specparam_declaration_instance9262();
    specparam_declaration9263 specparam_declaration_instance9263();
    specparam_declaration9264 specparam_declaration_instance9264();
    specparam_declaration9265 specparam_declaration_instance9265();
    specparam_declaration9266 specparam_declaration_instance9266();
    specparam_declaration9267 specparam_declaration_instance9267();
    specparam_declaration9268 specparam_declaration_instance9268();
    specparam_declaration9269 specparam_declaration_instance9269();
    specparam_declaration9270 specparam_declaration_instance9270();
    specparam_declaration9271 specparam_declaration_instance9271();
    specparam_declaration9272 specparam_declaration_instance9272();
    specparam_declaration9273 specparam_declaration_instance9273();
    specparam_declaration9274 specparam_declaration_instance9274();
    specparam_declaration9275 specparam_declaration_instance9275();
    specparam_declaration9276 specparam_declaration_instance9276();
    specparam_declaration9277 specparam_declaration_instance9277();
    specparam_declaration9278 specparam_declaration_instance9278();
    specparam_declaration9279 specparam_declaration_instance9279();
    specparam_declaration9280 specparam_declaration_instance9280();
    specparam_declaration9281 specparam_declaration_instance9281();
    specparam_declaration9282 specparam_declaration_instance9282();
    specparam_declaration9283 specparam_declaration_instance9283();
    specparam_declaration9284 specparam_declaration_instance9284();
    specparam_declaration9285 specparam_declaration_instance9285();
    specparam_declaration9286 specparam_declaration_instance9286();
    specparam_declaration9287 specparam_declaration_instance9287();
    specparam_declaration9288 specparam_declaration_instance9288();
    specparam_declaration9289 specparam_declaration_instance9289();
    specparam_declaration9290 specparam_declaration_instance9290();
    specparam_declaration9291 specparam_declaration_instance9291();
    specparam_declaration9292 specparam_declaration_instance9292();
    specparam_declaration9293 specparam_declaration_instance9293();
    specparam_declaration9294 specparam_declaration_instance9294();
    specparam_declaration9295 specparam_declaration_instance9295();
    specparam_declaration9296 specparam_declaration_instance9296();
    specparam_declaration9297 specparam_declaration_instance9297();
    specparam_declaration9298 specparam_declaration_instance9298();
    specparam_declaration9299 specparam_declaration_instance9299();
    specparam_declaration9300 specparam_declaration_instance9300();
    specparam_declaration9301 specparam_declaration_instance9301();
    specparam_declaration9302 specparam_declaration_instance9302();
    specparam_declaration9303 specparam_declaration_instance9303();
    specparam_declaration9304 specparam_declaration_instance9304();
    specparam_declaration9305 specparam_declaration_instance9305();
    specparam_declaration9306 specparam_declaration_instance9306();
    specparam_declaration9307 specparam_declaration_instance9307();
    specparam_declaration9308 specparam_declaration_instance9308();
    specparam_declaration9309 specparam_declaration_instance9309();
    specparam_declaration9310 specparam_declaration_instance9310();
    specparam_declaration9311 specparam_declaration_instance9311();
    specparam_declaration9312 specparam_declaration_instance9312();
    specparam_declaration9313 specparam_declaration_instance9313();
    specparam_declaration9314 specparam_declaration_instance9314();
    specparam_declaration9315 specparam_declaration_instance9315();
    specparam_declaration9316 specparam_declaration_instance9316();
    specparam_declaration9317 specparam_declaration_instance9317();
    specparam_declaration9318 specparam_declaration_instance9318();
    specparam_declaration9319 specparam_declaration_instance9319();
    specparam_declaration9320 specparam_declaration_instance9320();
    specparam_declaration9321 specparam_declaration_instance9321();
    specparam_declaration9322 specparam_declaration_instance9322();
    specparam_declaration9323 specparam_declaration_instance9323();
    specparam_declaration9324 specparam_declaration_instance9324();
    specparam_declaration9325 specparam_declaration_instance9325();
    specparam_declaration9326 specparam_declaration_instance9326();
    specparam_declaration9327 specparam_declaration_instance9327();
    specparam_declaration9328 specparam_declaration_instance9328();
    specparam_declaration9329 specparam_declaration_instance9329();
    specparam_declaration9330 specparam_declaration_instance9330();
    specparam_declaration9331 specparam_declaration_instance9331();
    specparam_declaration9332 specparam_declaration_instance9332();
    specparam_declaration9333 specparam_declaration_instance9333();
    specparam_declaration9334 specparam_declaration_instance9334();
    specparam_declaration9335 specparam_declaration_instance9335();
    specparam_declaration9336 specparam_declaration_instance9336();
    specparam_declaration9337 specparam_declaration_instance9337();
    specparam_declaration9338 specparam_declaration_instance9338();
    specparam_declaration9339 specparam_declaration_instance9339();
    specparam_declaration9340 specparam_declaration_instance9340();
    specparam_declaration9341 specparam_declaration_instance9341();
    specparam_declaration9342 specparam_declaration_instance9342();
    specparam_declaration9343 specparam_declaration_instance9343();
    specparam_declaration9344 specparam_declaration_instance9344();
    specparam_declaration9345 specparam_declaration_instance9345();
    specparam_declaration9346 specparam_declaration_instance9346();
    specparam_declaration9347 specparam_declaration_instance9347();
    specparam_declaration9348 specparam_declaration_instance9348();
    specparam_declaration9349 specparam_declaration_instance9349();
    specparam_declaration9350 specparam_declaration_instance9350();
    specparam_declaration9351 specparam_declaration_instance9351();
    specparam_declaration9352 specparam_declaration_instance9352();
    specparam_declaration9353 specparam_declaration_instance9353();
    specparam_declaration9354 specparam_declaration_instance9354();
    specparam_declaration9355 specparam_declaration_instance9355();
    specparam_declaration9356 specparam_declaration_instance9356();
    specparam_declaration9357 specparam_declaration_instance9357();
    specparam_declaration9358 specparam_declaration_instance9358();
    specparam_declaration9359 specparam_declaration_instance9359();
    specparam_declaration9360 specparam_declaration_instance9360();
    specparam_declaration9361 specparam_declaration_instance9361();
    specparam_declaration9362 specparam_declaration_instance9362();
    specparam_declaration9363 specparam_declaration_instance9363();
    specparam_declaration9364 specparam_declaration_instance9364();
    specparam_declaration9365 specparam_declaration_instance9365();
    specparam_declaration9366 specparam_declaration_instance9366();
    specparam_declaration9367 specparam_declaration_instance9367();
    specparam_declaration9368 specparam_declaration_instance9368();
    specparam_declaration9369 specparam_declaration_instance9369();
    specparam_declaration9370 specparam_declaration_instance9370();
    specparam_declaration9371 specparam_declaration_instance9371();
    specparam_declaration9372 specparam_declaration_instance9372();
    specparam_declaration9373 specparam_declaration_instance9373();
    specparam_declaration9374 specparam_declaration_instance9374();
    specparam_declaration9375 specparam_declaration_instance9375();
    specparam_declaration9376 specparam_declaration_instance9376();
    specparam_declaration9377 specparam_declaration_instance9377();
    specparam_declaration9378 specparam_declaration_instance9378();
    specparam_declaration9379 specparam_declaration_instance9379();
    specparam_declaration9380 specparam_declaration_instance9380();
    specparam_declaration9381 specparam_declaration_instance9381();
    specparam_declaration9382 specparam_declaration_instance9382();
    specparam_declaration9383 specparam_declaration_instance9383();
    specparam_declaration9384 specparam_declaration_instance9384();
    specparam_declaration9385 specparam_declaration_instance9385();
    specparam_declaration9386 specparam_declaration_instance9386();
    specparam_declaration9387 specparam_declaration_instance9387();
    specparam_declaration9388 specparam_declaration_instance9388();
    specparam_declaration9389 specparam_declaration_instance9389();
    specparam_declaration9390 specparam_declaration_instance9390();
    specparam_declaration9391 specparam_declaration_instance9391();
    specparam_declaration9392 specparam_declaration_instance9392();
    specparam_declaration9393 specparam_declaration_instance9393();
    specparam_declaration9394 specparam_declaration_instance9394();
    specparam_declaration9395 specparam_declaration_instance9395();
    specparam_declaration9396 specparam_declaration_instance9396();
    specparam_declaration9397 specparam_declaration_instance9397();
    specparam_declaration9398 specparam_declaration_instance9398();
    specparam_declaration9399 specparam_declaration_instance9399();
    specparam_declaration9400 specparam_declaration_instance9400();
    specparam_declaration9401 specparam_declaration_instance9401();
    specparam_declaration9402 specparam_declaration_instance9402();
    specparam_declaration9403 specparam_declaration_instance9403();
    specparam_declaration9404 specparam_declaration_instance9404();
    specparam_declaration9405 specparam_declaration_instance9405();
    specparam_declaration9406 specparam_declaration_instance9406();
    specparam_declaration9407 specparam_declaration_instance9407();
    specparam_declaration9408 specparam_declaration_instance9408();
    specparam_declaration9409 specparam_declaration_instance9409();
    specparam_declaration9410 specparam_declaration_instance9410();
    specparam_declaration9411 specparam_declaration_instance9411();
    specparam_declaration9412 specparam_declaration_instance9412();
    specparam_declaration9413 specparam_declaration_instance9413();
    specparam_declaration9414 specparam_declaration_instance9414();
    specparam_declaration9415 specparam_declaration_instance9415();
    specparam_declaration9416 specparam_declaration_instance9416();
    specparam_declaration9417 specparam_declaration_instance9417();
    specparam_declaration9418 specparam_declaration_instance9418();
    specparam_declaration9419 specparam_declaration_instance9419();
    specparam_declaration9420 specparam_declaration_instance9420();
    specparam_declaration9421 specparam_declaration_instance9421();
    specparam_declaration9422 specparam_declaration_instance9422();
    specparam_declaration9423 specparam_declaration_instance9423();
    specparam_declaration9424 specparam_declaration_instance9424();
    specparam_declaration9425 specparam_declaration_instance9425();
    specparam_declaration9426 specparam_declaration_instance9426();
    specparam_declaration9427 specparam_declaration_instance9427();
    specparam_declaration9428 specparam_declaration_instance9428();
    specparam_declaration9429 specparam_declaration_instance9429();
    specparam_declaration9430 specparam_declaration_instance9430();
    specparam_declaration9431 specparam_declaration_instance9431();
    specparam_declaration9432 specparam_declaration_instance9432();
    specparam_declaration9433 specparam_declaration_instance9433();
    specparam_declaration9434 specparam_declaration_instance9434();
    specparam_declaration9435 specparam_declaration_instance9435();
    specparam_declaration9436 specparam_declaration_instance9436();
    specparam_declaration9437 specparam_declaration_instance9437();
    specparam_declaration9438 specparam_declaration_instance9438();
    specparam_declaration9439 specparam_declaration_instance9439();
    specparam_declaration9440 specparam_declaration_instance9440();
    specparam_declaration9441 specparam_declaration_instance9441();
    specparam_declaration9442 specparam_declaration_instance9442();
    specparam_declaration9443 specparam_declaration_instance9443();
    specparam_declaration9444 specparam_declaration_instance9444();
    specparam_declaration9445 specparam_declaration_instance9445();
    specparam_declaration9446 specparam_declaration_instance9446();
    specparam_declaration9447 specparam_declaration_instance9447();
    specparam_declaration9448 specparam_declaration_instance9448();
    specparam_declaration9449 specparam_declaration_instance9449();
    specparam_declaration9450 specparam_declaration_instance9450();
    specparam_declaration9451 specparam_declaration_instance9451();
    specparam_declaration9452 specparam_declaration_instance9452();
    specparam_declaration9453 specparam_declaration_instance9453();
    specparam_declaration9454 specparam_declaration_instance9454();
    specparam_declaration9455 specparam_declaration_instance9455();
    specparam_declaration9456 specparam_declaration_instance9456();
    specparam_declaration9457 specparam_declaration_instance9457();
    specparam_declaration9458 specparam_declaration_instance9458();
    specparam_declaration9459 specparam_declaration_instance9459();
    specparam_declaration9460 specparam_declaration_instance9460();
    specparam_declaration9461 specparam_declaration_instance9461();
    specparam_declaration9462 specparam_declaration_instance9462();
    specparam_declaration9463 specparam_declaration_instance9463();
    specparam_declaration9464 specparam_declaration_instance9464();
    specparam_declaration9465 specparam_declaration_instance9465();
    specparam_declaration9466 specparam_declaration_instance9466();
    specparam_declaration9467 specparam_declaration_instance9467();
    specparam_declaration9468 specparam_declaration_instance9468();
    specparam_declaration9469 specparam_declaration_instance9469();
    specparam_declaration9470 specparam_declaration_instance9470();
    specparam_declaration9471 specparam_declaration_instance9471();
    specparam_declaration9472 specparam_declaration_instance9472();
    specparam_declaration9473 specparam_declaration_instance9473();
    specparam_declaration9474 specparam_declaration_instance9474();
    specparam_declaration9475 specparam_declaration_instance9475();
    specparam_declaration9476 specparam_declaration_instance9476();
    specparam_declaration9477 specparam_declaration_instance9477();
    specparam_declaration9478 specparam_declaration_instance9478();
    specparam_declaration9479 specparam_declaration_instance9479();
    specparam_declaration9480 specparam_declaration_instance9480();
    specparam_declaration9481 specparam_declaration_instance9481();
    specparam_declaration9482 specparam_declaration_instance9482();
    specparam_declaration9483 specparam_declaration_instance9483();
    specparam_declaration9484 specparam_declaration_instance9484();
    specparam_declaration9485 specparam_declaration_instance9485();
    specparam_declaration9486 specparam_declaration_instance9486();
    specparam_declaration9487 specparam_declaration_instance9487();
    specparam_declaration9488 specparam_declaration_instance9488();
    specparam_declaration9489 specparam_declaration_instance9489();
    specparam_declaration9490 specparam_declaration_instance9490();
    specparam_declaration9491 specparam_declaration_instance9491();
    specparam_declaration9492 specparam_declaration_instance9492();
    specparam_declaration9493 specparam_declaration_instance9493();
    specparam_declaration9494 specparam_declaration_instance9494();
    specparam_declaration9495 specparam_declaration_instance9495();
    specparam_declaration9496 specparam_declaration_instance9496();
    specparam_declaration9497 specparam_declaration_instance9497();
    specparam_declaration9498 specparam_declaration_instance9498();
    specparam_declaration9499 specparam_declaration_instance9499();
    specparam_declaration9500 specparam_declaration_instance9500();
    specparam_declaration9501 specparam_declaration_instance9501();
    specparam_declaration9502 specparam_declaration_instance9502();
    specparam_declaration9503 specparam_declaration_instance9503();
    specparam_declaration9504 specparam_declaration_instance9504();
    specparam_declaration9505 specparam_declaration_instance9505();
    specparam_declaration9506 specparam_declaration_instance9506();
    specparam_declaration9507 specparam_declaration_instance9507();
    specparam_declaration9508 specparam_declaration_instance9508();
    specparam_declaration9509 specparam_declaration_instance9509();
    specparam_declaration9510 specparam_declaration_instance9510();
    specparam_declaration9511 specparam_declaration_instance9511();
    specparam_declaration9512 specparam_declaration_instance9512();
    specparam_declaration9513 specparam_declaration_instance9513();
    specparam_declaration9514 specparam_declaration_instance9514();
    specparam_declaration9515 specparam_declaration_instance9515();
    specparam_declaration9516 specparam_declaration_instance9516();
    specparam_declaration9517 specparam_declaration_instance9517();
    specparam_declaration9518 specparam_declaration_instance9518();
    specparam_declaration9519 specparam_declaration_instance9519();
    specparam_declaration9520 specparam_declaration_instance9520();
    specparam_declaration9521 specparam_declaration_instance9521();
    specparam_declaration9522 specparam_declaration_instance9522();
    specparam_declaration9523 specparam_declaration_instance9523();
    specparam_declaration9524 specparam_declaration_instance9524();
    specparam_declaration9525 specparam_declaration_instance9525();
    specparam_declaration9526 specparam_declaration_instance9526();
    specparam_declaration9527 specparam_declaration_instance9527();
    specparam_declaration9528 specparam_declaration_instance9528();
    specparam_declaration9529 specparam_declaration_instance9529();
    specparam_declaration9530 specparam_declaration_instance9530();
    specparam_declaration9531 specparam_declaration_instance9531();
    specparam_declaration9532 specparam_declaration_instance9532();
    specparam_declaration9533 specparam_declaration_instance9533();
    specparam_declaration9534 specparam_declaration_instance9534();
    specparam_declaration9535 specparam_declaration_instance9535();
    specparam_declaration9536 specparam_declaration_instance9536();
    specparam_declaration9537 specparam_declaration_instance9537();
    specparam_declaration9538 specparam_declaration_instance9538();
    specparam_declaration9539 specparam_declaration_instance9539();
    specparam_declaration9540 specparam_declaration_instance9540();
    specparam_declaration9541 specparam_declaration_instance9541();
    specparam_declaration9542 specparam_declaration_instance9542();
    specparam_declaration9543 specparam_declaration_instance9543();
    specparam_declaration9544 specparam_declaration_instance9544();
    specparam_declaration9545 specparam_declaration_instance9545();
    specparam_declaration9546 specparam_declaration_instance9546();
    specparam_declaration9547 specparam_declaration_instance9547();
    specparam_declaration9548 specparam_declaration_instance9548();
    specparam_declaration9549 specparam_declaration_instance9549();
    specparam_declaration9550 specparam_declaration_instance9550();
    specparam_declaration9551 specparam_declaration_instance9551();
    specparam_declaration9552 specparam_declaration_instance9552();
    specparam_declaration9553 specparam_declaration_instance9553();
    specparam_declaration9554 specparam_declaration_instance9554();
    specparam_declaration9555 specparam_declaration_instance9555();
    specparam_declaration9556 specparam_declaration_instance9556();
    specparam_declaration9557 specparam_declaration_instance9557();
    specparam_declaration9558 specparam_declaration_instance9558();
    specparam_declaration9559 specparam_declaration_instance9559();
    specparam_declaration9560 specparam_declaration_instance9560();
    specparam_declaration9561 specparam_declaration_instance9561();
    specparam_declaration9562 specparam_declaration_instance9562();
    specparam_declaration9563 specparam_declaration_instance9563();
    specparam_declaration9564 specparam_declaration_instance9564();
    specparam_declaration9565 specparam_declaration_instance9565();
    specparam_declaration9566 specparam_declaration_instance9566();
    specparam_declaration9567 specparam_declaration_instance9567();
    specparam_declaration9568 specparam_declaration_instance9568();
    specparam_declaration9569 specparam_declaration_instance9569();
    specparam_declaration9570 specparam_declaration_instance9570();
    specparam_declaration9571 specparam_declaration_instance9571();
    specparam_declaration9572 specparam_declaration_instance9572();
    specparam_declaration9573 specparam_declaration_instance9573();
    specparam_declaration9574 specparam_declaration_instance9574();
    specparam_declaration9575 specparam_declaration_instance9575();
    specparam_declaration9576 specparam_declaration_instance9576();
    specparam_declaration9577 specparam_declaration_instance9577();
    specparam_declaration9578 specparam_declaration_instance9578();
    specparam_declaration9579 specparam_declaration_instance9579();
    specparam_declaration9580 specparam_declaration_instance9580();
    specparam_declaration9581 specparam_declaration_instance9581();
    specparam_declaration9582 specparam_declaration_instance9582();
    specparam_declaration9583 specparam_declaration_instance9583();
    specparam_declaration9584 specparam_declaration_instance9584();
    specparam_declaration9585 specparam_declaration_instance9585();
    specparam_declaration9586 specparam_declaration_instance9586();
    specparam_declaration9587 specparam_declaration_instance9587();
    specparam_declaration9588 specparam_declaration_instance9588();
    specparam_declaration9589 specparam_declaration_instance9589();
    specparam_declaration9590 specparam_declaration_instance9590();
    specparam_declaration9591 specparam_declaration_instance9591();
    specparam_declaration9592 specparam_declaration_instance9592();
    specparam_declaration9593 specparam_declaration_instance9593();
    specparam_declaration9594 specparam_declaration_instance9594();
    specparam_declaration9595 specparam_declaration_instance9595();
    specparam_declaration9596 specparam_declaration_instance9596();
    specparam_declaration9597 specparam_declaration_instance9597();
    specparam_declaration9598 specparam_declaration_instance9598();
    specparam_declaration9599 specparam_declaration_instance9599();
    specparam_declaration9600 specparam_declaration_instance9600();
    specparam_declaration9601 specparam_declaration_instance9601();
    specparam_declaration9602 specparam_declaration_instance9602();
    specparam_declaration9603 specparam_declaration_instance9603();
    specparam_declaration9604 specparam_declaration_instance9604();
    specparam_declaration9605 specparam_declaration_instance9605();
    specparam_declaration9606 specparam_declaration_instance9606();
    specparam_declaration9607 specparam_declaration_instance9607();
    specparam_declaration9608 specparam_declaration_instance9608();
    specparam_declaration9609 specparam_declaration_instance9609();
    specparam_declaration9610 specparam_declaration_instance9610();
    specparam_declaration9611 specparam_declaration_instance9611();
    specparam_declaration9612 specparam_declaration_instance9612();
    specparam_declaration9613 specparam_declaration_instance9613();
    specparam_declaration9614 specparam_declaration_instance9614();
    specparam_declaration9615 specparam_declaration_instance9615();
    specparam_declaration9616 specparam_declaration_instance9616();
    specparam_declaration9617 specparam_declaration_instance9617();
    specparam_declaration9618 specparam_declaration_instance9618();
    specparam_declaration9619 specparam_declaration_instance9619();
    specparam_declaration9620 specparam_declaration_instance9620();
    specparam_declaration9621 specparam_declaration_instance9621();
    specparam_declaration9622 specparam_declaration_instance9622();
    specparam_declaration9623 specparam_declaration_instance9623();
    specparam_declaration9624 specparam_declaration_instance9624();
    specparam_declaration9625 specparam_declaration_instance9625();
    specparam_declaration9626 specparam_declaration_instance9626();
    specparam_declaration9627 specparam_declaration_instance9627();
    specparam_declaration9628 specparam_declaration_instance9628();
    specparam_declaration9629 specparam_declaration_instance9629();
    specparam_declaration9630 specparam_declaration_instance9630();
    specparam_declaration9631 specparam_declaration_instance9631();
    specparam_declaration9632 specparam_declaration_instance9632();
    specparam_declaration9633 specparam_declaration_instance9633();
    specparam_declaration9634 specparam_declaration_instance9634();
    specparam_declaration9635 specparam_declaration_instance9635();
    specparam_declaration9636 specparam_declaration_instance9636();
    specparam_declaration9637 specparam_declaration_instance9637();
    specparam_declaration9638 specparam_declaration_instance9638();
    specparam_declaration9639 specparam_declaration_instance9639();
    specparam_declaration9640 specparam_declaration_instance9640();
    specparam_declaration9641 specparam_declaration_instance9641();
    specparam_declaration9642 specparam_declaration_instance9642();
    specparam_declaration9643 specparam_declaration_instance9643();
    specparam_declaration9644 specparam_declaration_instance9644();
    specparam_declaration9645 specparam_declaration_instance9645();
    specparam_declaration9646 specparam_declaration_instance9646();
    specparam_declaration9647 specparam_declaration_instance9647();
    specparam_declaration9648 specparam_declaration_instance9648();
    specparam_declaration9649 specparam_declaration_instance9649();
    specparam_declaration9650 specparam_declaration_instance9650();
    specparam_declaration9651 specparam_declaration_instance9651();
    specparam_declaration9652 specparam_declaration_instance9652();
    specparam_declaration9653 specparam_declaration_instance9653();
    specparam_declaration9654 specparam_declaration_instance9654();
    specparam_declaration9655 specparam_declaration_instance9655();
    specparam_declaration9656 specparam_declaration_instance9656();
    specparam_declaration9657 specparam_declaration_instance9657();
    specparam_declaration9658 specparam_declaration_instance9658();
    specparam_declaration9659 specparam_declaration_instance9659();
    specparam_declaration9660 specparam_declaration_instance9660();
    specparam_declaration9661 specparam_declaration_instance9661();
    specparam_declaration9662 specparam_declaration_instance9662();
    specparam_declaration9663 specparam_declaration_instance9663();
    specparam_declaration9664 specparam_declaration_instance9664();
    specparam_declaration9665 specparam_declaration_instance9665();
    specparam_declaration9666 specparam_declaration_instance9666();
    specparam_declaration9667 specparam_declaration_instance9667();
    specparam_declaration9668 specparam_declaration_instance9668();
    specparam_declaration9669 specparam_declaration_instance9669();
    specparam_declaration9670 specparam_declaration_instance9670();
    specparam_declaration9671 specparam_declaration_instance9671();
    specparam_declaration9672 specparam_declaration_instance9672();
    specparam_declaration9673 specparam_declaration_instance9673();
    specparam_declaration9674 specparam_declaration_instance9674();
    specparam_declaration9675 specparam_declaration_instance9675();
    specparam_declaration9676 specparam_declaration_instance9676();
    specparam_declaration9677 specparam_declaration_instance9677();
    specparam_declaration9678 specparam_declaration_instance9678();
    specparam_declaration9679 specparam_declaration_instance9679();
    specparam_declaration9680 specparam_declaration_instance9680();
    specparam_declaration9681 specparam_declaration_instance9681();
    specparam_declaration9682 specparam_declaration_instance9682();
    specparam_declaration9683 specparam_declaration_instance9683();
    specparam_declaration9684 specparam_declaration_instance9684();
    specparam_declaration9685 specparam_declaration_instance9685();
    specparam_declaration9686 specparam_declaration_instance9686();
    specparam_declaration9687 specparam_declaration_instance9687();
    specparam_declaration9688 specparam_declaration_instance9688();
    specparam_declaration9689 specparam_declaration_instance9689();
    specparam_declaration9690 specparam_declaration_instance9690();
    specparam_declaration9691 specparam_declaration_instance9691();
    specparam_declaration9692 specparam_declaration_instance9692();
    specparam_declaration9693 specparam_declaration_instance9693();
    specparam_declaration9694 specparam_declaration_instance9694();
    specparam_declaration9695 specparam_declaration_instance9695();
    specparam_declaration9696 specparam_declaration_instance9696();
    specparam_declaration9697 specparam_declaration_instance9697();
    specparam_declaration9698 specparam_declaration_instance9698();
    specparam_declaration9699 specparam_declaration_instance9699();
    specparam_declaration9700 specparam_declaration_instance9700();
    specparam_declaration9701 specparam_declaration_instance9701();
    specparam_declaration9702 specparam_declaration_instance9702();
    specparam_declaration9703 specparam_declaration_instance9703();
    specparam_declaration9704 specparam_declaration_instance9704();
    specparam_declaration9705 specparam_declaration_instance9705();
    specparam_declaration9706 specparam_declaration_instance9706();
    specparam_declaration9707 specparam_declaration_instance9707();
    specparam_declaration9708 specparam_declaration_instance9708();
    specparam_declaration9709 specparam_declaration_instance9709();
    specparam_declaration9710 specparam_declaration_instance9710();
    specparam_declaration9711 specparam_declaration_instance9711();
    specparam_declaration9712 specparam_declaration_instance9712();
    specparam_declaration9713 specparam_declaration_instance9713();
    specparam_declaration9714 specparam_declaration_instance9714();
    specparam_declaration9715 specparam_declaration_instance9715();
    specparam_declaration9716 specparam_declaration_instance9716();
    specparam_declaration9717 specparam_declaration_instance9717();
    specparam_declaration9718 specparam_declaration_instance9718();
    specparam_declaration9719 specparam_declaration_instance9719();
    specparam_declaration9720 specparam_declaration_instance9720();
    specparam_declaration9721 specparam_declaration_instance9721();
    specparam_declaration9722 specparam_declaration_instance9722();
    specparam_declaration9723 specparam_declaration_instance9723();
    specparam_declaration9724 specparam_declaration_instance9724();
    specparam_declaration9725 specparam_declaration_instance9725();
    specparam_declaration9726 specparam_declaration_instance9726();
    specparam_declaration9727 specparam_declaration_instance9727();
    specparam_declaration9728 specparam_declaration_instance9728();
    specparam_declaration9729 specparam_declaration_instance9729();
    specparam_declaration9730 specparam_declaration_instance9730();
    specparam_declaration9731 specparam_declaration_instance9731();
    specparam_declaration9732 specparam_declaration_instance9732();
    specparam_declaration9733 specparam_declaration_instance9733();
    specparam_declaration9734 specparam_declaration_instance9734();
    specparam_declaration9735 specparam_declaration_instance9735();
    specparam_declaration9736 specparam_declaration_instance9736();
    specparam_declaration9737 specparam_declaration_instance9737();
    specparam_declaration9738 specparam_declaration_instance9738();
    specparam_declaration9739 specparam_declaration_instance9739();
    specparam_declaration9740 specparam_declaration_instance9740();
    specparam_declaration9741 specparam_declaration_instance9741();
    specparam_declaration9742 specparam_declaration_instance9742();
    specparam_declaration9743 specparam_declaration_instance9743();
    specparam_declaration9744 specparam_declaration_instance9744();
    specparam_declaration9745 specparam_declaration_instance9745();
    specparam_declaration9746 specparam_declaration_instance9746();
    specparam_declaration9747 specparam_declaration_instance9747();
    specparam_declaration9748 specparam_declaration_instance9748();
    specparam_declaration9749 specparam_declaration_instance9749();
    specparam_declaration9750 specparam_declaration_instance9750();
    specparam_declaration9751 specparam_declaration_instance9751();
    specparam_declaration9752 specparam_declaration_instance9752();
    specparam_declaration9753 specparam_declaration_instance9753();
    specparam_declaration9754 specparam_declaration_instance9754();
    specparam_declaration9755 specparam_declaration_instance9755();
    specparam_declaration9756 specparam_declaration_instance9756();
    specparam_declaration9757 specparam_declaration_instance9757();
    specparam_declaration9758 specparam_declaration_instance9758();
    specparam_declaration9759 specparam_declaration_instance9759();
    specparam_declaration9760 specparam_declaration_instance9760();
    specparam_declaration9761 specparam_declaration_instance9761();
    specparam_declaration9762 specparam_declaration_instance9762();
    specparam_declaration9763 specparam_declaration_instance9763();
    specparam_declaration9764 specparam_declaration_instance9764();
    specparam_declaration9765 specparam_declaration_instance9765();
    specparam_declaration9766 specparam_declaration_instance9766();
    specparam_declaration9767 specparam_declaration_instance9767();
    specparam_declaration9768 specparam_declaration_instance9768();
    specparam_declaration9769 specparam_declaration_instance9769();
    specparam_declaration9770 specparam_declaration_instance9770();
    specparam_declaration9771 specparam_declaration_instance9771();
    specparam_declaration9772 specparam_declaration_instance9772();
    specparam_declaration9773 specparam_declaration_instance9773();
    specparam_declaration9774 specparam_declaration_instance9774();
    specparam_declaration9775 specparam_declaration_instance9775();
    specparam_declaration9776 specparam_declaration_instance9776();
    specparam_declaration9777 specparam_declaration_instance9777();
    specparam_declaration9778 specparam_declaration_instance9778();
    specparam_declaration9779 specparam_declaration_instance9779();
    specparam_declaration9780 specparam_declaration_instance9780();
    specparam_declaration9781 specparam_declaration_instance9781();
    specparam_declaration9782 specparam_declaration_instance9782();
    specparam_declaration9783 specparam_declaration_instance9783();
    specparam_declaration9784 specparam_declaration_instance9784();
    specparam_declaration9785 specparam_declaration_instance9785();
    specparam_declaration9786 specparam_declaration_instance9786();
    specparam_declaration9787 specparam_declaration_instance9787();
    specparam_declaration9788 specparam_declaration_instance9788();
    specparam_declaration9789 specparam_declaration_instance9789();
    specparam_declaration9790 specparam_declaration_instance9790();
    specparam_declaration9791 specparam_declaration_instance9791();
    specparam_declaration9792 specparam_declaration_instance9792();
    specparam_declaration9793 specparam_declaration_instance9793();
    specparam_declaration9794 specparam_declaration_instance9794();
    specparam_declaration9795 specparam_declaration_instance9795();
    specparam_declaration9796 specparam_declaration_instance9796();
    specparam_declaration9797 specparam_declaration_instance9797();
    specparam_declaration9798 specparam_declaration_instance9798();
    specparam_declaration9799 specparam_declaration_instance9799();
    specparam_declaration9800 specparam_declaration_instance9800();
    specparam_declaration9801 specparam_declaration_instance9801();
    specparam_declaration9802 specparam_declaration_instance9802();
    specparam_declaration9803 specparam_declaration_instance9803();
    specparam_declaration9804 specparam_declaration_instance9804();
    specparam_declaration9805 specparam_declaration_instance9805();
    specparam_declaration9806 specparam_declaration_instance9806();
    specparam_declaration9807 specparam_declaration_instance9807();
    specparam_declaration9808 specparam_declaration_instance9808();
    specparam_declaration9809 specparam_declaration_instance9809();
    specparam_declaration9810 specparam_declaration_instance9810();
    specparam_declaration9811 specparam_declaration_instance9811();
    specparam_declaration9812 specparam_declaration_instance9812();
    specparam_declaration9813 specparam_declaration_instance9813();
    specparam_declaration9814 specparam_declaration_instance9814();
    specparam_declaration9815 specparam_declaration_instance9815();
    specparam_declaration9816 specparam_declaration_instance9816();
    specparam_declaration9817 specparam_declaration_instance9817();
    specparam_declaration9818 specparam_declaration_instance9818();
    specparam_declaration9819 specparam_declaration_instance9819();
    specparam_declaration9820 specparam_declaration_instance9820();
    specparam_declaration9821 specparam_declaration_instance9821();
    specparam_declaration9822 specparam_declaration_instance9822();
    specparam_declaration9823 specparam_declaration_instance9823();
    specparam_declaration9824 specparam_declaration_instance9824();
    specparam_declaration9825 specparam_declaration_instance9825();
    specparam_declaration9826 specparam_declaration_instance9826();
    specparam_declaration9827 specparam_declaration_instance9827();
    specparam_declaration9828 specparam_declaration_instance9828();
    specparam_declaration9829 specparam_declaration_instance9829();
    specparam_declaration9830 specparam_declaration_instance9830();
    specparam_declaration9831 specparam_declaration_instance9831();
    specparam_declaration9832 specparam_declaration_instance9832();
    specparam_declaration9833 specparam_declaration_instance9833();
    specparam_declaration9834 specparam_declaration_instance9834();
    specparam_declaration9835 specparam_declaration_instance9835();
    specparam_declaration9836 specparam_declaration_instance9836();
    specparam_declaration9837 specparam_declaration_instance9837();
    specparam_declaration9838 specparam_declaration_instance9838();
    specparam_declaration9839 specparam_declaration_instance9839();
    specparam_declaration9840 specparam_declaration_instance9840();
    specparam_declaration9841 specparam_declaration_instance9841();
    specparam_declaration9842 specparam_declaration_instance9842();
    specparam_declaration9843 specparam_declaration_instance9843();
    specparam_declaration9844 specparam_declaration_instance9844();
    specparam_declaration9845 specparam_declaration_instance9845();
    specparam_declaration9846 specparam_declaration_instance9846();
    specparam_declaration9847 specparam_declaration_instance9847();
    specparam_declaration9848 specparam_declaration_instance9848();
    specparam_declaration9849 specparam_declaration_instance9849();
    specparam_declaration9850 specparam_declaration_instance9850();
    specparam_declaration9851 specparam_declaration_instance9851();
    specparam_declaration9852 specparam_declaration_instance9852();
    specparam_declaration9853 specparam_declaration_instance9853();
    specparam_declaration9854 specparam_declaration_instance9854();
    specparam_declaration9855 specparam_declaration_instance9855();
    specparam_declaration9856 specparam_declaration_instance9856();
    specparam_declaration9857 specparam_declaration_instance9857();
    specparam_declaration9858 specparam_declaration_instance9858();
    specparam_declaration9859 specparam_declaration_instance9859();
    specparam_declaration9860 specparam_declaration_instance9860();
    specparam_declaration9861 specparam_declaration_instance9861();
    specparam_declaration9862 specparam_declaration_instance9862();
    specparam_declaration9863 specparam_declaration_instance9863();
    specparam_declaration9864 specparam_declaration_instance9864();
    specparam_declaration9865 specparam_declaration_instance9865();
    specparam_declaration9866 specparam_declaration_instance9866();
    specparam_declaration9867 specparam_declaration_instance9867();
    specparam_declaration9868 specparam_declaration_instance9868();
    specparam_declaration9869 specparam_declaration_instance9869();
    specparam_declaration9870 specparam_declaration_instance9870();
    specparam_declaration9871 specparam_declaration_instance9871();
    specparam_declaration9872 specparam_declaration_instance9872();
    specparam_declaration9873 specparam_declaration_instance9873();
    specparam_declaration9874 specparam_declaration_instance9874();
    specparam_declaration9875 specparam_declaration_instance9875();
    specparam_declaration9876 specparam_declaration_instance9876();
    specparam_declaration9877 specparam_declaration_instance9877();
    specparam_declaration9878 specparam_declaration_instance9878();
    specparam_declaration9879 specparam_declaration_instance9879();
    specparam_declaration9880 specparam_declaration_instance9880();
    specparam_declaration9881 specparam_declaration_instance9881();
    specparam_declaration9882 specparam_declaration_instance9882();
    specparam_declaration9883 specparam_declaration_instance9883();
    specparam_declaration9884 specparam_declaration_instance9884();
    specparam_declaration9885 specparam_declaration_instance9885();
    specparam_declaration9886 specparam_declaration_instance9886();
    specparam_declaration9887 specparam_declaration_instance9887();
    specparam_declaration9888 specparam_declaration_instance9888();
    specparam_declaration9889 specparam_declaration_instance9889();
    specparam_declaration9890 specparam_declaration_instance9890();
    specparam_declaration9891 specparam_declaration_instance9891();
    specparam_declaration9892 specparam_declaration_instance9892();
    specparam_declaration9893 specparam_declaration_instance9893();
    specparam_declaration9894 specparam_declaration_instance9894();
    specparam_declaration9895 specparam_declaration_instance9895();
    specparam_declaration9896 specparam_declaration_instance9896();
    specparam_declaration9897 specparam_declaration_instance9897();
    specparam_declaration9898 specparam_declaration_instance9898();
    specparam_declaration9899 specparam_declaration_instance9899();
    specparam_declaration9900 specparam_declaration_instance9900();
    specparam_declaration9901 specparam_declaration_instance9901();
    specparam_declaration9902 specparam_declaration_instance9902();
    specparam_declaration9903 specparam_declaration_instance9903();
    specparam_declaration9904 specparam_declaration_instance9904();
    specparam_declaration9905 specparam_declaration_instance9905();
    specparam_declaration9906 specparam_declaration_instance9906();
    specparam_declaration9907 specparam_declaration_instance9907();
    specparam_declaration9908 specparam_declaration_instance9908();
    specparam_declaration9909 specparam_declaration_instance9909();
    specparam_declaration9910 specparam_declaration_instance9910();
    specparam_declaration9911 specparam_declaration_instance9911();
    specparam_declaration9912 specparam_declaration_instance9912();
    specparam_declaration9913 specparam_declaration_instance9913();
    specparam_declaration9914 specparam_declaration_instance9914();
    specparam_declaration9915 specparam_declaration_instance9915();
    specparam_declaration9916 specparam_declaration_instance9916();
    specparam_declaration9917 specparam_declaration_instance9917();
    specparam_declaration9918 specparam_declaration_instance9918();
    specparam_declaration9919 specparam_declaration_instance9919();
    specparam_declaration9920 specparam_declaration_instance9920();
    specparam_declaration9921 specparam_declaration_instance9921();
    specparam_declaration9922 specparam_declaration_instance9922();
    specparam_declaration9923 specparam_declaration_instance9923();
    specparam_declaration9924 specparam_declaration_instance9924();
    specparam_declaration9925 specparam_declaration_instance9925();
    specparam_declaration9926 specparam_declaration_instance9926();
    specparam_declaration9927 specparam_declaration_instance9927();
    specparam_declaration9928 specparam_declaration_instance9928();
    specparam_declaration9929 specparam_declaration_instance9929();
    specparam_declaration9930 specparam_declaration_instance9930();
    specparam_declaration9931 specparam_declaration_instance9931();
    specparam_declaration9932 specparam_declaration_instance9932();
    specparam_declaration9933 specparam_declaration_instance9933();
    specparam_declaration9934 specparam_declaration_instance9934();
    specparam_declaration9935 specparam_declaration_instance9935();
    specparam_declaration9936 specparam_declaration_instance9936();
    specparam_declaration9937 specparam_declaration_instance9937();
    specparam_declaration9938 specparam_declaration_instance9938();
    specparam_declaration9939 specparam_declaration_instance9939();
    specparam_declaration9940 specparam_declaration_instance9940();
    specparam_declaration9941 specparam_declaration_instance9941();
    specparam_declaration9942 specparam_declaration_instance9942();
    specparam_declaration9943 specparam_declaration_instance9943();
    specparam_declaration9944 specparam_declaration_instance9944();
    specparam_declaration9945 specparam_declaration_instance9945();
    specparam_declaration9946 specparam_declaration_instance9946();
    specparam_declaration9947 specparam_declaration_instance9947();
    specparam_declaration9948 specparam_declaration_instance9948();
    specparam_declaration9949 specparam_declaration_instance9949();
    specparam_declaration9950 specparam_declaration_instance9950();
    specparam_declaration9951 specparam_declaration_instance9951();
    specparam_declaration9952 specparam_declaration_instance9952();
    specparam_declaration9953 specparam_declaration_instance9953();
    specparam_declaration9954 specparam_declaration_instance9954();
    specparam_declaration9955 specparam_declaration_instance9955();
    specparam_declaration9956 specparam_declaration_instance9956();
    specparam_declaration9957 specparam_declaration_instance9957();
    specparam_declaration9958 specparam_declaration_instance9958();
    specparam_declaration9959 specparam_declaration_instance9959();
    specparam_declaration9960 specparam_declaration_instance9960();
    specparam_declaration9961 specparam_declaration_instance9961();
    specparam_declaration9962 specparam_declaration_instance9962();
    specparam_declaration9963 specparam_declaration_instance9963();
    specparam_declaration9964 specparam_declaration_instance9964();
    specparam_declaration9965 specparam_declaration_instance9965();
    specparam_declaration9966 specparam_declaration_instance9966();
    specparam_declaration9967 specparam_declaration_instance9967();
    specparam_declaration9968 specparam_declaration_instance9968();
    specparam_declaration9969 specparam_declaration_instance9969();
    specparam_declaration9970 specparam_declaration_instance9970();
    specparam_declaration9971 specparam_declaration_instance9971();
    specparam_declaration9972 specparam_declaration_instance9972();
    specparam_declaration9973 specparam_declaration_instance9973();
    specparam_declaration9974 specparam_declaration_instance9974();
    specparam_declaration9975 specparam_declaration_instance9975();
    specparam_declaration9976 specparam_declaration_instance9976();
    specparam_declaration9977 specparam_declaration_instance9977();
    specparam_declaration9978 specparam_declaration_instance9978();
    specparam_declaration9979 specparam_declaration_instance9979();
    specparam_declaration9980 specparam_declaration_instance9980();
    specparam_declaration9981 specparam_declaration_instance9981();
    specparam_declaration9982 specparam_declaration_instance9982();
    specparam_declaration9983 specparam_declaration_instance9983();
    specparam_declaration9984 specparam_declaration_instance9984();
    specparam_declaration9985 specparam_declaration_instance9985();
    specparam_declaration9986 specparam_declaration_instance9986();
    specparam_declaration9987 specparam_declaration_instance9987();
    specparam_declaration9988 specparam_declaration_instance9988();
    specparam_declaration9989 specparam_declaration_instance9989();
    specparam_declaration9990 specparam_declaration_instance9990();
    specparam_declaration9991 specparam_declaration_instance9991();
    specparam_declaration9992 specparam_declaration_instance9992();
    specparam_declaration9993 specparam_declaration_instance9993();
    specparam_declaration9994 specparam_declaration_instance9994();
    specparam_declaration9995 specparam_declaration_instance9995();
    specparam_declaration9996 specparam_declaration_instance9996();
    specparam_declaration9997 specparam_declaration_instance9997();
    specparam_declaration9998 specparam_declaration_instance9998();
    specparam_declaration9999 specparam_declaration_instance9999();
    specparam_declaration10000 specparam_declaration_instance10000();
    specparam_declaration10001 specparam_declaration_instance10001();
    specparam_declaration10002 specparam_declaration_instance10002();
    specparam_declaration10003 specparam_declaration_instance10003();
    specparam_declaration10004 specparam_declaration_instance10004();
    specparam_declaration10005 specparam_declaration_instance10005();
    specparam_declaration10006 specparam_declaration_instance10006();
    specparam_declaration10007 specparam_declaration_instance10007();
    specparam_declaration10008 specparam_declaration_instance10008();
    specparam_declaration10009 specparam_declaration_instance10009();
    specparam_declaration10010 specparam_declaration_instance10010();
    specparam_declaration10011 specparam_declaration_instance10011();
    specparam_declaration10012 specparam_declaration_instance10012();
    specparam_declaration10013 specparam_declaration_instance10013();
    specparam_declaration10014 specparam_declaration_instance10014();
    specparam_declaration10015 specparam_declaration_instance10015();
    specparam_declaration10016 specparam_declaration_instance10016();
    specparam_declaration10017 specparam_declaration_instance10017();
    specparam_declaration10018 specparam_declaration_instance10018();
    specparam_declaration10019 specparam_declaration_instance10019();
    specparam_declaration10020 specparam_declaration_instance10020();
    specparam_declaration10021 specparam_declaration_instance10021();
    specparam_declaration10022 specparam_declaration_instance10022();
    specparam_declaration10023 specparam_declaration_instance10023();
    specparam_declaration10024 specparam_declaration_instance10024();
    specparam_declaration10025 specparam_declaration_instance10025();
    specparam_declaration10026 specparam_declaration_instance10026();
    specparam_declaration10027 specparam_declaration_instance10027();
    specparam_declaration10028 specparam_declaration_instance10028();
    specparam_declaration10029 specparam_declaration_instance10029();
    specparam_declaration10030 specparam_declaration_instance10030();
    specparam_declaration10031 specparam_declaration_instance10031();
    specparam_declaration10032 specparam_declaration_instance10032();
    specparam_declaration10033 specparam_declaration_instance10033();
    specparam_declaration10034 specparam_declaration_instance10034();
    specparam_declaration10035 specparam_declaration_instance10035();
    specparam_declaration10036 specparam_declaration_instance10036();
    specparam_declaration10037 specparam_declaration_instance10037();
    specparam_declaration10038 specparam_declaration_instance10038();
    specparam_declaration10039 specparam_declaration_instance10039();
    specparam_declaration10040 specparam_declaration_instance10040();
    specparam_declaration10041 specparam_declaration_instance10041();
    specparam_declaration10042 specparam_declaration_instance10042();
    specparam_declaration10043 specparam_declaration_instance10043();
    specparam_declaration10044 specparam_declaration_instance10044();
    specparam_declaration10045 specparam_declaration_instance10045();
    specparam_declaration10046 specparam_declaration_instance10046();
    specparam_declaration10047 specparam_declaration_instance10047();
    specparam_declaration10048 specparam_declaration_instance10048();
    specparam_declaration10049 specparam_declaration_instance10049();
    specparam_declaration10050 specparam_declaration_instance10050();
    specparam_declaration10051 specparam_declaration_instance10051();
    specparam_declaration10052 specparam_declaration_instance10052();
    specparam_declaration10053 specparam_declaration_instance10053();
    specparam_declaration10054 specparam_declaration_instance10054();
    specparam_declaration10055 specparam_declaration_instance10055();
    specparam_declaration10056 specparam_declaration_instance10056();
    specparam_declaration10057 specparam_declaration_instance10057();
    specparam_declaration10058 specparam_declaration_instance10058();
    specparam_declaration10059 specparam_declaration_instance10059();
    specparam_declaration10060 specparam_declaration_instance10060();
    specparam_declaration10061 specparam_declaration_instance10061();
    specparam_declaration10062 specparam_declaration_instance10062();
    specparam_declaration10063 specparam_declaration_instance10063();
    specparam_declaration10064 specparam_declaration_instance10064();
    specparam_declaration10065 specparam_declaration_instance10065();
    specparam_declaration10066 specparam_declaration_instance10066();
    specparam_declaration10067 specparam_declaration_instance10067();
    specparam_declaration10068 specparam_declaration_instance10068();
    specparam_declaration10069 specparam_declaration_instance10069();
    specparam_declaration10070 specparam_declaration_instance10070();
    specparam_declaration10071 specparam_declaration_instance10071();
    specparam_declaration10072 specparam_declaration_instance10072();
    specparam_declaration10073 specparam_declaration_instance10073();
    specparam_declaration10074 specparam_declaration_instance10074();
    specparam_declaration10075 specparam_declaration_instance10075();
    specparam_declaration10076 specparam_declaration_instance10076();
    specparam_declaration10077 specparam_declaration_instance10077();
    specparam_declaration10078 specparam_declaration_instance10078();
    specparam_declaration10079 specparam_declaration_instance10079();
    specparam_declaration10080 specparam_declaration_instance10080();
    specparam_declaration10081 specparam_declaration_instance10081();
    specparam_declaration10082 specparam_declaration_instance10082();
    specparam_declaration10083 specparam_declaration_instance10083();
    specparam_declaration10084 specparam_declaration_instance10084();
    specparam_declaration10085 specparam_declaration_instance10085();
    specparam_declaration10086 specparam_declaration_instance10086();
    specparam_declaration10087 specparam_declaration_instance10087();
    specparam_declaration10088 specparam_declaration_instance10088();
    specparam_declaration10089 specparam_declaration_instance10089();
    specparam_declaration10090 specparam_declaration_instance10090();
    specparam_declaration10091 specparam_declaration_instance10091();
    specparam_declaration10092 specparam_declaration_instance10092();
    specparam_declaration10093 specparam_declaration_instance10093();
    specparam_declaration10094 specparam_declaration_instance10094();
    specparam_declaration10095 specparam_declaration_instance10095();
    specparam_declaration10096 specparam_declaration_instance10096();
    specparam_declaration10097 specparam_declaration_instance10097();
    specparam_declaration10098 specparam_declaration_instance10098();
    specparam_declaration10099 specparam_declaration_instance10099();
    specparam_declaration10100 specparam_declaration_instance10100();
    specparam_declaration10101 specparam_declaration_instance10101();
    specparam_declaration10102 specparam_declaration_instance10102();
    specparam_declaration10103 specparam_declaration_instance10103();
    specparam_declaration10104 specparam_declaration_instance10104();
    specparam_declaration10105 specparam_declaration_instance10105();
    specparam_declaration10106 specparam_declaration_instance10106();
    specparam_declaration10107 specparam_declaration_instance10107();
    specparam_declaration10108 specparam_declaration_instance10108();
    specparam_declaration10109 specparam_declaration_instance10109();
    specparam_declaration10110 specparam_declaration_instance10110();
    specparam_declaration10111 specparam_declaration_instance10111();
    specparam_declaration10112 specparam_declaration_instance10112();
    specparam_declaration10113 specparam_declaration_instance10113();
    specparam_declaration10114 specparam_declaration_instance10114();
    specparam_declaration10115 specparam_declaration_instance10115();
    specparam_declaration10116 specparam_declaration_instance10116();
    specparam_declaration10117 specparam_declaration_instance10117();
    specparam_declaration10118 specparam_declaration_instance10118();
    specparam_declaration10119 specparam_declaration_instance10119();
    specparam_declaration10120 specparam_declaration_instance10120();
    specparam_declaration10121 specparam_declaration_instance10121();
    specparam_declaration10122 specparam_declaration_instance10122();
    specparam_declaration10123 specparam_declaration_instance10123();
    specparam_declaration10124 specparam_declaration_instance10124();
    specparam_declaration10125 specparam_declaration_instance10125();
    specparam_declaration10126 specparam_declaration_instance10126();
    specparam_declaration10127 specparam_declaration_instance10127();
    specparam_declaration10128 specparam_declaration_instance10128();
    specparam_declaration10129 specparam_declaration_instance10129();
    specparam_declaration10130 specparam_declaration_instance10130();
    specparam_declaration10131 specparam_declaration_instance10131();
    specparam_declaration10132 specparam_declaration_instance10132();
    specparam_declaration10133 specparam_declaration_instance10133();
    specparam_declaration10134 specparam_declaration_instance10134();
    specparam_declaration10135 specparam_declaration_instance10135();
    specparam_declaration10136 specparam_declaration_instance10136();
    specparam_declaration10137 specparam_declaration_instance10137();
    specparam_declaration10138 specparam_declaration_instance10138();
    specparam_declaration10139 specparam_declaration_instance10139();
    specparam_declaration10140 specparam_declaration_instance10140();
    specparam_declaration10141 specparam_declaration_instance10141();
    specparam_declaration10142 specparam_declaration_instance10142();
    specparam_declaration10143 specparam_declaration_instance10143();
    specparam_declaration10144 specparam_declaration_instance10144();
    specparam_declaration10145 specparam_declaration_instance10145();
    specparam_declaration10146 specparam_declaration_instance10146();
    specparam_declaration10147 specparam_declaration_instance10147();
    specparam_declaration10148 specparam_declaration_instance10148();
    specparam_declaration10149 specparam_declaration_instance10149();
    specparam_declaration10150 specparam_declaration_instance10150();
    specparam_declaration10151 specparam_declaration_instance10151();
    specparam_declaration10152 specparam_declaration_instance10152();
    specparam_declaration10153 specparam_declaration_instance10153();
    specparam_declaration10154 specparam_declaration_instance10154();
    specparam_declaration10155 specparam_declaration_instance10155();
    specparam_declaration10156 specparam_declaration_instance10156();
    specparam_declaration10157 specparam_declaration_instance10157();
    specparam_declaration10158 specparam_declaration_instance10158();
    specparam_declaration10159 specparam_declaration_instance10159();
    specparam_declaration10160 specparam_declaration_instance10160();
    specparam_declaration10161 specparam_declaration_instance10161();
    specparam_declaration10162 specparam_declaration_instance10162();
    specparam_declaration10163 specparam_declaration_instance10163();
    specparam_declaration10164 specparam_declaration_instance10164();
    specparam_declaration10165 specparam_declaration_instance10165();
    specparam_declaration10166 specparam_declaration_instance10166();
    specparam_declaration10167 specparam_declaration_instance10167();
    specparam_declaration10168 specparam_declaration_instance10168();
    specparam_declaration10169 specparam_declaration_instance10169();
    specparam_declaration10170 specparam_declaration_instance10170();
    specparam_declaration10171 specparam_declaration_instance10171();
    specparam_declaration10172 specparam_declaration_instance10172();
    specparam_declaration10173 specparam_declaration_instance10173();
    specparam_declaration10174 specparam_declaration_instance10174();
    specparam_declaration10175 specparam_declaration_instance10175();
    specparam_declaration10176 specparam_declaration_instance10176();
    specparam_declaration10177 specparam_declaration_instance10177();
    specparam_declaration10178 specparam_declaration_instance10178();
    specparam_declaration10179 specparam_declaration_instance10179();
    specparam_declaration10180 specparam_declaration_instance10180();
    specparam_declaration10181 specparam_declaration_instance10181();
    specparam_declaration10182 specparam_declaration_instance10182();
    specparam_declaration10183 specparam_declaration_instance10183();
    specparam_declaration10184 specparam_declaration_instance10184();
    specparam_declaration10185 specparam_declaration_instance10185();
    specparam_declaration10186 specparam_declaration_instance10186();
    specparam_declaration10187 specparam_declaration_instance10187();
    specparam_declaration10188 specparam_declaration_instance10188();
    specparam_declaration10189 specparam_declaration_instance10189();
    specparam_declaration10190 specparam_declaration_instance10190();
    specparam_declaration10191 specparam_declaration_instance10191();
    specparam_declaration10192 specparam_declaration_instance10192();
    specparam_declaration10193 specparam_declaration_instance10193();
    specparam_declaration10194 specparam_declaration_instance10194();
    specparam_declaration10195 specparam_declaration_instance10195();
    specparam_declaration10196 specparam_declaration_instance10196();
    specparam_declaration10197 specparam_declaration_instance10197();
    specparam_declaration10198 specparam_declaration_instance10198();
    specparam_declaration10199 specparam_declaration_instance10199();
    specparam_declaration10200 specparam_declaration_instance10200();
    specparam_declaration10201 specparam_declaration_instance10201();
    specparam_declaration10202 specparam_declaration_instance10202();
    specparam_declaration10203 specparam_declaration_instance10203();
    specparam_declaration10204 specparam_declaration_instance10204();
    specparam_declaration10205 specparam_declaration_instance10205();
    specparam_declaration10206 specparam_declaration_instance10206();
    specparam_declaration10207 specparam_declaration_instance10207();
    specparam_declaration10208 specparam_declaration_instance10208();
    specparam_declaration10209 specparam_declaration_instance10209();
    specparam_declaration10210 specparam_declaration_instance10210();
    specparam_declaration10211 specparam_declaration_instance10211();
    specparam_declaration10212 specparam_declaration_instance10212();
    specparam_declaration10213 specparam_declaration_instance10213();
    specparam_declaration10214 specparam_declaration_instance10214();
    specparam_declaration10215 specparam_declaration_instance10215();
    specparam_declaration10216 specparam_declaration_instance10216();
    specparam_declaration10217 specparam_declaration_instance10217();
    specparam_declaration10218 specparam_declaration_instance10218();
    specparam_declaration10219 specparam_declaration_instance10219();
    specparam_declaration10220 specparam_declaration_instance10220();
    specparam_declaration10221 specparam_declaration_instance10221();
    specparam_declaration10222 specparam_declaration_instance10222();
    specparam_declaration10223 specparam_declaration_instance10223();
    specparam_declaration10224 specparam_declaration_instance10224();
    specparam_declaration10225 specparam_declaration_instance10225();
    specparam_declaration10226 specparam_declaration_instance10226();
    specparam_declaration10227 specparam_declaration_instance10227();
    specparam_declaration10228 specparam_declaration_instance10228();
    specparam_declaration10229 specparam_declaration_instance10229();
    specparam_declaration10230 specparam_declaration_instance10230();
    specparam_declaration10231 specparam_declaration_instance10231();
    specparam_declaration10232 specparam_declaration_instance10232();
    specparam_declaration10233 specparam_declaration_instance10233();
    specparam_declaration10234 specparam_declaration_instance10234();
    specparam_declaration10235 specparam_declaration_instance10235();
    specparam_declaration10236 specparam_declaration_instance10236();
    specparam_declaration10237 specparam_declaration_instance10237();
    specparam_declaration10238 specparam_declaration_instance10238();
    specparam_declaration10239 specparam_declaration_instance10239();
    specparam_declaration10240 specparam_declaration_instance10240();
    specparam_declaration10241 specparam_declaration_instance10241();
    specparam_declaration10242 specparam_declaration_instance10242();
    specparam_declaration10243 specparam_declaration_instance10243();
    specparam_declaration10244 specparam_declaration_instance10244();
    specparam_declaration10245 specparam_declaration_instance10245();
    specparam_declaration10246 specparam_declaration_instance10246();
    specparam_declaration10247 specparam_declaration_instance10247();
    specparam_declaration10248 specparam_declaration_instance10248();
    specparam_declaration10249 specparam_declaration_instance10249();
    specparam_declaration10250 specparam_declaration_instance10250();
    specparam_declaration10251 specparam_declaration_instance10251();
    specparam_declaration10252 specparam_declaration_instance10252();
    specparam_declaration10253 specparam_declaration_instance10253();
    specparam_declaration10254 specparam_declaration_instance10254();
    specparam_declaration10255 specparam_declaration_instance10255();
    specparam_declaration10256 specparam_declaration_instance10256();
    specparam_declaration10257 specparam_declaration_instance10257();
    specparam_declaration10258 specparam_declaration_instance10258();
    specparam_declaration10259 specparam_declaration_instance10259();
    specparam_declaration10260 specparam_declaration_instance10260();
    specparam_declaration10261 specparam_declaration_instance10261();
    specparam_declaration10262 specparam_declaration_instance10262();
    specparam_declaration10263 specparam_declaration_instance10263();
    specparam_declaration10264 specparam_declaration_instance10264();
    specparam_declaration10265 specparam_declaration_instance10265();
    specparam_declaration10266 specparam_declaration_instance10266();
    specparam_declaration10267 specparam_declaration_instance10267();
    specparam_declaration10268 specparam_declaration_instance10268();
    specparam_declaration10269 specparam_declaration_instance10269();
    specparam_declaration10270 specparam_declaration_instance10270();
    specparam_declaration10271 specparam_declaration_instance10271();
    specparam_declaration10272 specparam_declaration_instance10272();
    specparam_declaration10273 specparam_declaration_instance10273();
    specparam_declaration10274 specparam_declaration_instance10274();
    specparam_declaration10275 specparam_declaration_instance10275();
    specparam_declaration10276 specparam_declaration_instance10276();
    specparam_declaration10277 specparam_declaration_instance10277();
    specparam_declaration10278 specparam_declaration_instance10278();
    specparam_declaration10279 specparam_declaration_instance10279();
    specparam_declaration10280 specparam_declaration_instance10280();
    specparam_declaration10281 specparam_declaration_instance10281();
    specparam_declaration10282 specparam_declaration_instance10282();
    specparam_declaration10283 specparam_declaration_instance10283();
    specparam_declaration10284 specparam_declaration_instance10284();
    specparam_declaration10285 specparam_declaration_instance10285();
    specparam_declaration10286 specparam_declaration_instance10286();
    specparam_declaration10287 specparam_declaration_instance10287();
    specparam_declaration10288 specparam_declaration_instance10288();
    specparam_declaration10289 specparam_declaration_instance10289();
    specparam_declaration10290 specparam_declaration_instance10290();
    specparam_declaration10291 specparam_declaration_instance10291();
    specparam_declaration10292 specparam_declaration_instance10292();
    specparam_declaration10293 specparam_declaration_instance10293();
    specparam_declaration10294 specparam_declaration_instance10294();
    specparam_declaration10295 specparam_declaration_instance10295();
    specparam_declaration10296 specparam_declaration_instance10296();
    specparam_declaration10297 specparam_declaration_instance10297();
    specparam_declaration10298 specparam_declaration_instance10298();
    specparam_declaration10299 specparam_declaration_instance10299();
    specparam_declaration10300 specparam_declaration_instance10300();
    specparam_declaration10301 specparam_declaration_instance10301();
    specparam_declaration10302 specparam_declaration_instance10302();
    specparam_declaration10303 specparam_declaration_instance10303();
    specparam_declaration10304 specparam_declaration_instance10304();
    specparam_declaration10305 specparam_declaration_instance10305();
    specparam_declaration10306 specparam_declaration_instance10306();
    specparam_declaration10307 specparam_declaration_instance10307();
    specparam_declaration10308 specparam_declaration_instance10308();
    specparam_declaration10309 specparam_declaration_instance10309();
    specparam_declaration10310 specparam_declaration_instance10310();
    specparam_declaration10311 specparam_declaration_instance10311();
    specparam_declaration10312 specparam_declaration_instance10312();
    specparam_declaration10313 specparam_declaration_instance10313();
    specparam_declaration10314 specparam_declaration_instance10314();
    specparam_declaration10315 specparam_declaration_instance10315();
    specparam_declaration10316 specparam_declaration_instance10316();
    specparam_declaration10317 specparam_declaration_instance10317();
    specparam_declaration10318 specparam_declaration_instance10318();
    specparam_declaration10319 specparam_declaration_instance10319();
    specparam_declaration10320 specparam_declaration_instance10320();
    specparam_declaration10321 specparam_declaration_instance10321();
    specparam_declaration10322 specparam_declaration_instance10322();
    specparam_declaration10323 specparam_declaration_instance10323();
    specparam_declaration10324 specparam_declaration_instance10324();
    specparam_declaration10325 specparam_declaration_instance10325();
    specparam_declaration10326 specparam_declaration_instance10326();
    specparam_declaration10327 specparam_declaration_instance10327();
    specparam_declaration10328 specparam_declaration_instance10328();
    specparam_declaration10329 specparam_declaration_instance10329();
    specparam_declaration10330 specparam_declaration_instance10330();
    specparam_declaration10331 specparam_declaration_instance10331();
    specparam_declaration10332 specparam_declaration_instance10332();
    specparam_declaration10333 specparam_declaration_instance10333();
    specparam_declaration10334 specparam_declaration_instance10334();
    specparam_declaration10335 specparam_declaration_instance10335();
    specparam_declaration10336 specparam_declaration_instance10336();
    specparam_declaration10337 specparam_declaration_instance10337();
    specparam_declaration10338 specparam_declaration_instance10338();
    specparam_declaration10339 specparam_declaration_instance10339();
    specparam_declaration10340 specparam_declaration_instance10340();
    specparam_declaration10341 specparam_declaration_instance10341();
    specparam_declaration10342 specparam_declaration_instance10342();
    specparam_declaration10343 specparam_declaration_instance10343();
    specparam_declaration10344 specparam_declaration_instance10344();
    specparam_declaration10345 specparam_declaration_instance10345();
    specparam_declaration10346 specparam_declaration_instance10346();
    specparam_declaration10347 specparam_declaration_instance10347();
    specparam_declaration10348 specparam_declaration_instance10348();
    specparam_declaration10349 specparam_declaration_instance10349();
    specparam_declaration10350 specparam_declaration_instance10350();
    specparam_declaration10351 specparam_declaration_instance10351();
    specparam_declaration10352 specparam_declaration_instance10352();
    specparam_declaration10353 specparam_declaration_instance10353();
    specparam_declaration10354 specparam_declaration_instance10354();
    specparam_declaration10355 specparam_declaration_instance10355();
    specparam_declaration10356 specparam_declaration_instance10356();
    specparam_declaration10357 specparam_declaration_instance10357();
    specparam_declaration10358 specparam_declaration_instance10358();
    specparam_declaration10359 specparam_declaration_instance10359();
    specparam_declaration10360 specparam_declaration_instance10360();
    specparam_declaration10361 specparam_declaration_instance10361();
    specparam_declaration10362 specparam_declaration_instance10362();
    specparam_declaration10363 specparam_declaration_instance10363();
    specparam_declaration10364 specparam_declaration_instance10364();
    specparam_declaration10365 specparam_declaration_instance10365();
    specparam_declaration10366 specparam_declaration_instance10366();
    specparam_declaration10367 specparam_declaration_instance10367();
    specparam_declaration10368 specparam_declaration_instance10368();
    specparam_declaration10369 specparam_declaration_instance10369();
    specparam_declaration10370 specparam_declaration_instance10370();
    specparam_declaration10371 specparam_declaration_instance10371();
    specparam_declaration10372 specparam_declaration_instance10372();
    specparam_declaration10373 specparam_declaration_instance10373();
    specparam_declaration10374 specparam_declaration_instance10374();
    specparam_declaration10375 specparam_declaration_instance10375();
    specparam_declaration10376 specparam_declaration_instance10376();
    specparam_declaration10377 specparam_declaration_instance10377();
    specparam_declaration10378 specparam_declaration_instance10378();
    specparam_declaration10379 specparam_declaration_instance10379();
    specparam_declaration10380 specparam_declaration_instance10380();
    specparam_declaration10381 specparam_declaration_instance10381();
    specparam_declaration10382 specparam_declaration_instance10382();
    specparam_declaration10383 specparam_declaration_instance10383();
    specparam_declaration10384 specparam_declaration_instance10384();
    specparam_declaration10385 specparam_declaration_instance10385();
    specparam_declaration10386 specparam_declaration_instance10386();
    specparam_declaration10387 specparam_declaration_instance10387();
    specparam_declaration10388 specparam_declaration_instance10388();
    specparam_declaration10389 specparam_declaration_instance10389();
    specparam_declaration10390 specparam_declaration_instance10390();
    specparam_declaration10391 specparam_declaration_instance10391();
    specparam_declaration10392 specparam_declaration_instance10392();
    specparam_declaration10393 specparam_declaration_instance10393();
    specparam_declaration10394 specparam_declaration_instance10394();
    specparam_declaration10395 specparam_declaration_instance10395();
    specparam_declaration10396 specparam_declaration_instance10396();
    specparam_declaration10397 specparam_declaration_instance10397();
    specparam_declaration10398 specparam_declaration_instance10398();
    specparam_declaration10399 specparam_declaration_instance10399();
    specparam_declaration10400 specparam_declaration_instance10400();
    specparam_declaration10401 specparam_declaration_instance10401();
    specparam_declaration10402 specparam_declaration_instance10402();
    specparam_declaration10403 specparam_declaration_instance10403();
    specparam_declaration10404 specparam_declaration_instance10404();
    specparam_declaration10405 specparam_declaration_instance10405();
    specparam_declaration10406 specparam_declaration_instance10406();
    specparam_declaration10407 specparam_declaration_instance10407();
    specparam_declaration10408 specparam_declaration_instance10408();
    specparam_declaration10409 specparam_declaration_instance10409();
    specparam_declaration10410 specparam_declaration_instance10410();
    specparam_declaration10411 specparam_declaration_instance10411();
    specparam_declaration10412 specparam_declaration_instance10412();
    specparam_declaration10413 specparam_declaration_instance10413();
    specparam_declaration10414 specparam_declaration_instance10414();
    specparam_declaration10415 specparam_declaration_instance10415();
    specparam_declaration10416 specparam_declaration_instance10416();
    specparam_declaration10417 specparam_declaration_instance10417();
    specparam_declaration10418 specparam_declaration_instance10418();
    specparam_declaration10419 specparam_declaration_instance10419();
    specparam_declaration10420 specparam_declaration_instance10420();
    specparam_declaration10421 specparam_declaration_instance10421();
    specparam_declaration10422 specparam_declaration_instance10422();
    specparam_declaration10423 specparam_declaration_instance10423();
    specparam_declaration10424 specparam_declaration_instance10424();
    specparam_declaration10425 specparam_declaration_instance10425();
    specparam_declaration10426 specparam_declaration_instance10426();
    specparam_declaration10427 specparam_declaration_instance10427();
    specparam_declaration10428 specparam_declaration_instance10428();
    specparam_declaration10429 specparam_declaration_instance10429();
    specparam_declaration10430 specparam_declaration_instance10430();
    specparam_declaration10431 specparam_declaration_instance10431();
    specparam_declaration10432 specparam_declaration_instance10432();
    specparam_declaration10433 specparam_declaration_instance10433();
    specparam_declaration10434 specparam_declaration_instance10434();
    specparam_declaration10435 specparam_declaration_instance10435();
    specparam_declaration10436 specparam_declaration_instance10436();
    specparam_declaration10437 specparam_declaration_instance10437();
    specparam_declaration10438 specparam_declaration_instance10438();
    specparam_declaration10439 specparam_declaration_instance10439();
    specparam_declaration10440 specparam_declaration_instance10440();
    specparam_declaration10441 specparam_declaration_instance10441();
    specparam_declaration10442 specparam_declaration_instance10442();
    specparam_declaration10443 specparam_declaration_instance10443();
    specparam_declaration10444 specparam_declaration_instance10444();
    specparam_declaration10445 specparam_declaration_instance10445();
    specparam_declaration10446 specparam_declaration_instance10446();
    specparam_declaration10447 specparam_declaration_instance10447();
    specparam_declaration10448 specparam_declaration_instance10448();
    specparam_declaration10449 specparam_declaration_instance10449();
    specparam_declaration10450 specparam_declaration_instance10450();
    specparam_declaration10451 specparam_declaration_instance10451();
    specparam_declaration10452 specparam_declaration_instance10452();
    specparam_declaration10453 specparam_declaration_instance10453();
    specparam_declaration10454 specparam_declaration_instance10454();
    specparam_declaration10455 specparam_declaration_instance10455();
    specparam_declaration10456 specparam_declaration_instance10456();
    specparam_declaration10457 specparam_declaration_instance10457();
    specparam_declaration10458 specparam_declaration_instance10458();
    specparam_declaration10459 specparam_declaration_instance10459();
    specparam_declaration10460 specparam_declaration_instance10460();
    specparam_declaration10461 specparam_declaration_instance10461();
    specparam_declaration10462 specparam_declaration_instance10462();
    specparam_declaration10463 specparam_declaration_instance10463();
    specparam_declaration10464 specparam_declaration_instance10464();
    specparam_declaration10465 specparam_declaration_instance10465();
    specparam_declaration10466 specparam_declaration_instance10466();
    specparam_declaration10467 specparam_declaration_instance10467();
    specparam_declaration10468 specparam_declaration_instance10468();
    specparam_declaration10469 specparam_declaration_instance10469();
    specparam_declaration10470 specparam_declaration_instance10470();
    specparam_declaration10471 specparam_declaration_instance10471();
    specparam_declaration10472 specparam_declaration_instance10472();
    specparam_declaration10473 specparam_declaration_instance10473();
    specparam_declaration10474 specparam_declaration_instance10474();
    specparam_declaration10475 specparam_declaration_instance10475();
    specparam_declaration10476 specparam_declaration_instance10476();
    specparam_declaration10477 specparam_declaration_instance10477();
    specparam_declaration10478 specparam_declaration_instance10478();
    specparam_declaration10479 specparam_declaration_instance10479();
    specparam_declaration10480 specparam_declaration_instance10480();
    specparam_declaration10481 specparam_declaration_instance10481();
    specparam_declaration10482 specparam_declaration_instance10482();
    specparam_declaration10483 specparam_declaration_instance10483();
    specparam_declaration10484 specparam_declaration_instance10484();
    specparam_declaration10485 specparam_declaration_instance10485();
    specparam_declaration10486 specparam_declaration_instance10486();
    specparam_declaration10487 specparam_declaration_instance10487();
    specparam_declaration10488 specparam_declaration_instance10488();
    specparam_declaration10489 specparam_declaration_instance10489();
    specparam_declaration10490 specparam_declaration_instance10490();
    specparam_declaration10491 specparam_declaration_instance10491();
    specparam_declaration10492 specparam_declaration_instance10492();
    specparam_declaration10493 specparam_declaration_instance10493();
    specparam_declaration10494 specparam_declaration_instance10494();
    specparam_declaration10495 specparam_declaration_instance10495();
    specparam_declaration10496 specparam_declaration_instance10496();
    specparam_declaration10497 specparam_declaration_instance10497();
    specparam_declaration10498 specparam_declaration_instance10498();
    specparam_declaration10499 specparam_declaration_instance10499();
    specparam_declaration10500 specparam_declaration_instance10500();
    specparam_declaration10501 specparam_declaration_instance10501();
    specparam_declaration10502 specparam_declaration_instance10502();
    specparam_declaration10503 specparam_declaration_instance10503();
    specparam_declaration10504 specparam_declaration_instance10504();
    specparam_declaration10505 specparam_declaration_instance10505();
    specparam_declaration10506 specparam_declaration_instance10506();
    specparam_declaration10507 specparam_declaration_instance10507();
    specparam_declaration10508 specparam_declaration_instance10508();
    specparam_declaration10509 specparam_declaration_instance10509();
    specparam_declaration10510 specparam_declaration_instance10510();
    specparam_declaration10511 specparam_declaration_instance10511();
    specparam_declaration10512 specparam_declaration_instance10512();
    specparam_declaration10513 specparam_declaration_instance10513();
    specparam_declaration10514 specparam_declaration_instance10514();
    specparam_declaration10515 specparam_declaration_instance10515();
    specparam_declaration10516 specparam_declaration_instance10516();
    specparam_declaration10517 specparam_declaration_instance10517();
    specparam_declaration10518 specparam_declaration_instance10518();
    specparam_declaration10519 specparam_declaration_instance10519();
    specparam_declaration10520 specparam_declaration_instance10520();
    specparam_declaration10521 specparam_declaration_instance10521();
    specparam_declaration10522 specparam_declaration_instance10522();
    specparam_declaration10523 specparam_declaration_instance10523();
    specparam_declaration10524 specparam_declaration_instance10524();
    specparam_declaration10525 specparam_declaration_instance10525();
    specparam_declaration10526 specparam_declaration_instance10526();
    specparam_declaration10527 specparam_declaration_instance10527();
    specparam_declaration10528 specparam_declaration_instance10528();
    specparam_declaration10529 specparam_declaration_instance10529();
    specparam_declaration10530 specparam_declaration_instance10530();
    specparam_declaration10531 specparam_declaration_instance10531();
    specparam_declaration10532 specparam_declaration_instance10532();
    specparam_declaration10533 specparam_declaration_instance10533();
    specparam_declaration10534 specparam_declaration_instance10534();
    specparam_declaration10535 specparam_declaration_instance10535();
    specparam_declaration10536 specparam_declaration_instance10536();
    specparam_declaration10537 specparam_declaration_instance10537();
    specparam_declaration10538 specparam_declaration_instance10538();
    specparam_declaration10539 specparam_declaration_instance10539();
    specparam_declaration10540 specparam_declaration_instance10540();
    specparam_declaration10541 specparam_declaration_instance10541();
    specparam_declaration10542 specparam_declaration_instance10542();
    specparam_declaration10543 specparam_declaration_instance10543();
    specparam_declaration10544 specparam_declaration_instance10544();
    specparam_declaration10545 specparam_declaration_instance10545();
    specparam_declaration10546 specparam_declaration_instance10546();
    specparam_declaration10547 specparam_declaration_instance10547();
    specparam_declaration10548 specparam_declaration_instance10548();
    specparam_declaration10549 specparam_declaration_instance10549();
    specparam_declaration10550 specparam_declaration_instance10550();
    specparam_declaration10551 specparam_declaration_instance10551();
    specparam_declaration10552 specparam_declaration_instance10552();
    specparam_declaration10553 specparam_declaration_instance10553();
    specparam_declaration10554 specparam_declaration_instance10554();
    specparam_declaration10555 specparam_declaration_instance10555();
    specparam_declaration10556 specparam_declaration_instance10556();
    specparam_declaration10557 specparam_declaration_instance10557();
    specparam_declaration10558 specparam_declaration_instance10558();
    specparam_declaration10559 specparam_declaration_instance10559();
    specparam_declaration10560 specparam_declaration_instance10560();
    specparam_declaration10561 specparam_declaration_instance10561();
    specparam_declaration10562 specparam_declaration_instance10562();
    specparam_declaration10563 specparam_declaration_instance10563();
    specparam_declaration10564 specparam_declaration_instance10564();
    specparam_declaration10565 specparam_declaration_instance10565();
    specparam_declaration10566 specparam_declaration_instance10566();
    specparam_declaration10567 specparam_declaration_instance10567();
    specparam_declaration10568 specparam_declaration_instance10568();
    specparam_declaration10569 specparam_declaration_instance10569();
    specparam_declaration10570 specparam_declaration_instance10570();
    specparam_declaration10571 specparam_declaration_instance10571();
    specparam_declaration10572 specparam_declaration_instance10572();
    specparam_declaration10573 specparam_declaration_instance10573();
    specparam_declaration10574 specparam_declaration_instance10574();
    specparam_declaration10575 specparam_declaration_instance10575();
    specparam_declaration10576 specparam_declaration_instance10576();
    specparam_declaration10577 specparam_declaration_instance10577();
    specparam_declaration10578 specparam_declaration_instance10578();
    specparam_declaration10579 specparam_declaration_instance10579();
    specparam_declaration10580 specparam_declaration_instance10580();
    specparam_declaration10581 specparam_declaration_instance10581();
    specparam_declaration10582 specparam_declaration_instance10582();
    specparam_declaration10583 specparam_declaration_instance10583();
    specparam_declaration10584 specparam_declaration_instance10584();
    specparam_declaration10585 specparam_declaration_instance10585();
    specparam_declaration10586 specparam_declaration_instance10586();
    specparam_declaration10587 specparam_declaration_instance10587();
    specparam_declaration10588 specparam_declaration_instance10588();
    specparam_declaration10589 specparam_declaration_instance10589();
    specparam_declaration10590 specparam_declaration_instance10590();
    specparam_declaration10591 specparam_declaration_instance10591();
    specparam_declaration10592 specparam_declaration_instance10592();
    specparam_declaration10593 specparam_declaration_instance10593();
    specparam_declaration10594 specparam_declaration_instance10594();
    specparam_declaration10595 specparam_declaration_instance10595();
    specparam_declaration10596 specparam_declaration_instance10596();
    specparam_declaration10597 specparam_declaration_instance10597();
    specparam_declaration10598 specparam_declaration_instance10598();
    specparam_declaration10599 specparam_declaration_instance10599();
    specparam_declaration10600 specparam_declaration_instance10600();
    specparam_declaration10601 specparam_declaration_instance10601();
    specparam_declaration10602 specparam_declaration_instance10602();
    specparam_declaration10603 specparam_declaration_instance10603();
    specparam_declaration10604 specparam_declaration_instance10604();
    specparam_declaration10605 specparam_declaration_instance10605();
    specparam_declaration10606 specparam_declaration_instance10606();
    specparam_declaration10607 specparam_declaration_instance10607();
    specparam_declaration10608 specparam_declaration_instance10608();
    specparam_declaration10609 specparam_declaration_instance10609();
    specparam_declaration10610 specparam_declaration_instance10610();
    specparam_declaration10611 specparam_declaration_instance10611();
    specparam_declaration10612 specparam_declaration_instance10612();
    specparam_declaration10613 specparam_declaration_instance10613();
    specparam_declaration10614 specparam_declaration_instance10614();
    specparam_declaration10615 specparam_declaration_instance10615();
    specparam_declaration10616 specparam_declaration_instance10616();
    specparam_declaration10617 specparam_declaration_instance10617();
    specparam_declaration10618 specparam_declaration_instance10618();
    specparam_declaration10619 specparam_declaration_instance10619();
    specparam_declaration10620 specparam_declaration_instance10620();
    specparam_declaration10621 specparam_declaration_instance10621();
    specparam_declaration10622 specparam_declaration_instance10622();
    specparam_declaration10623 specparam_declaration_instance10623();
    specparam_declaration10624 specparam_declaration_instance10624();
    specparam_declaration10625 specparam_declaration_instance10625();
    specparam_declaration10626 specparam_declaration_instance10626();
    specparam_declaration10627 specparam_declaration_instance10627();
    specparam_declaration10628 specparam_declaration_instance10628();
    specparam_declaration10629 specparam_declaration_instance10629();
    specparam_declaration10630 specparam_declaration_instance10630();
    specparam_declaration10631 specparam_declaration_instance10631();
    specparam_declaration10632 specparam_declaration_instance10632();
    specparam_declaration10633 specparam_declaration_instance10633();
    specparam_declaration10634 specparam_declaration_instance10634();
    specparam_declaration10635 specparam_declaration_instance10635();
    specparam_declaration10636 specparam_declaration_instance10636();
    specparam_declaration10637 specparam_declaration_instance10637();
    specparam_declaration10638 specparam_declaration_instance10638();
    specparam_declaration10639 specparam_declaration_instance10639();
    specparam_declaration10640 specparam_declaration_instance10640();
    specparam_declaration10641 specparam_declaration_instance10641();
    specparam_declaration10642 specparam_declaration_instance10642();
    specparam_declaration10643 specparam_declaration_instance10643();
    specparam_declaration10644 specparam_declaration_instance10644();
    specparam_declaration10645 specparam_declaration_instance10645();
    specparam_declaration10646 specparam_declaration_instance10646();
    specparam_declaration10647 specparam_declaration_instance10647();
    specparam_declaration10648 specparam_declaration_instance10648();
    specparam_declaration10649 specparam_declaration_instance10649();
    specparam_declaration10650 specparam_declaration_instance10650();
    specparam_declaration10651 specparam_declaration_instance10651();
    specparam_declaration10652 specparam_declaration_instance10652();
    specparam_declaration10653 specparam_declaration_instance10653();
    specparam_declaration10654 specparam_declaration_instance10654();
    specparam_declaration10655 specparam_declaration_instance10655();
    specparam_declaration10656 specparam_declaration_instance10656();
    specparam_declaration10657 specparam_declaration_instance10657();
    specparam_declaration10658 specparam_declaration_instance10658();
    specparam_declaration10659 specparam_declaration_instance10659();
    specparam_declaration10660 specparam_declaration_instance10660();
    specparam_declaration10661 specparam_declaration_instance10661();
    specparam_declaration10662 specparam_declaration_instance10662();
    specparam_declaration10663 specparam_declaration_instance10663();
    specparam_declaration10664 specparam_declaration_instance10664();
    specparam_declaration10665 specparam_declaration_instance10665();
    specparam_declaration10666 specparam_declaration_instance10666();
    specparam_declaration10667 specparam_declaration_instance10667();
    specparam_declaration10668 specparam_declaration_instance10668();
    specparam_declaration10669 specparam_declaration_instance10669();
    specparam_declaration10670 specparam_declaration_instance10670();
    specparam_declaration10671 specparam_declaration_instance10671();
    specparam_declaration10672 specparam_declaration_instance10672();
    specparam_declaration10673 specparam_declaration_instance10673();
    specparam_declaration10674 specparam_declaration_instance10674();
    specparam_declaration10675 specparam_declaration_instance10675();
    specparam_declaration10676 specparam_declaration_instance10676();
    specparam_declaration10677 specparam_declaration_instance10677();
    specparam_declaration10678 specparam_declaration_instance10678();
    specparam_declaration10679 specparam_declaration_instance10679();
    specparam_declaration10680 specparam_declaration_instance10680();
    specparam_declaration10681 specparam_declaration_instance10681();
    specparam_declaration10682 specparam_declaration_instance10682();
    specparam_declaration10683 specparam_declaration_instance10683();
    specparam_declaration10684 specparam_declaration_instance10684();
    specparam_declaration10685 specparam_declaration_instance10685();
    specparam_declaration10686 specparam_declaration_instance10686();
    specparam_declaration10687 specparam_declaration_instance10687();
    specparam_declaration10688 specparam_declaration_instance10688();
    specparam_declaration10689 specparam_declaration_instance10689();
    specparam_declaration10690 specparam_declaration_instance10690();
    specparam_declaration10691 specparam_declaration_instance10691();
    specparam_declaration10692 specparam_declaration_instance10692();
    specparam_declaration10693 specparam_declaration_instance10693();
    specparam_declaration10694 specparam_declaration_instance10694();
    specparam_declaration10695 specparam_declaration_instance10695();
    specparam_declaration10696 specparam_declaration_instance10696();
    specparam_declaration10697 specparam_declaration_instance10697();
    specparam_declaration10698 specparam_declaration_instance10698();
    specparam_declaration10699 specparam_declaration_instance10699();
    specparam_declaration10700 specparam_declaration_instance10700();
    specparam_declaration10701 specparam_declaration_instance10701();
    specparam_declaration10702 specparam_declaration_instance10702();
    specparam_declaration10703 specparam_declaration_instance10703();
    specparam_declaration10704 specparam_declaration_instance10704();
    specparam_declaration10705 specparam_declaration_instance10705();
    specparam_declaration10706 specparam_declaration_instance10706();
    specparam_declaration10707 specparam_declaration_instance10707();
    specparam_declaration10708 specparam_declaration_instance10708();
    specparam_declaration10709 specparam_declaration_instance10709();
    specparam_declaration10710 specparam_declaration_instance10710();
    specparam_declaration10711 specparam_declaration_instance10711();
    specparam_declaration10712 specparam_declaration_instance10712();
    specparam_declaration10713 specparam_declaration_instance10713();
    specparam_declaration10714 specparam_declaration_instance10714();
    specparam_declaration10715 specparam_declaration_instance10715();
    specparam_declaration10716 specparam_declaration_instance10716();
    specparam_declaration10717 specparam_declaration_instance10717();
    specparam_declaration10718 specparam_declaration_instance10718();
    specparam_declaration10719 specparam_declaration_instance10719();
    specparam_declaration10720 specparam_declaration_instance10720();
    specparam_declaration10721 specparam_declaration_instance10721();
    specparam_declaration10722 specparam_declaration_instance10722();
    specparam_declaration10723 specparam_declaration_instance10723();
    specparam_declaration10724 specparam_declaration_instance10724();
    specparam_declaration10725 specparam_declaration_instance10725();
    specparam_declaration10726 specparam_declaration_instance10726();
    specparam_declaration10727 specparam_declaration_instance10727();
    specparam_declaration10728 specparam_declaration_instance10728();
    specparam_declaration10729 specparam_declaration_instance10729();
    specparam_declaration10730 specparam_declaration_instance10730();
    specparam_declaration10731 specparam_declaration_instance10731();
    specparam_declaration10732 specparam_declaration_instance10732();
    specparam_declaration10733 specparam_declaration_instance10733();
    specparam_declaration10734 specparam_declaration_instance10734();
    specparam_declaration10735 specparam_declaration_instance10735();
    specparam_declaration10736 specparam_declaration_instance10736();
    specparam_declaration10737 specparam_declaration_instance10737();
    specparam_declaration10738 specparam_declaration_instance10738();
    specparam_declaration10739 specparam_declaration_instance10739();
    specparam_declaration10740 specparam_declaration_instance10740();
    specparam_declaration10741 specparam_declaration_instance10741();
    specparam_declaration10742 specparam_declaration_instance10742();
    specparam_declaration10743 specparam_declaration_instance10743();
    specparam_declaration10744 specparam_declaration_instance10744();
    specparam_declaration10745 specparam_declaration_instance10745();
    specparam_declaration10746 specparam_declaration_instance10746();
    specparam_declaration10747 specparam_declaration_instance10747();
    specparam_declaration10748 specparam_declaration_instance10748();
    specparam_declaration10749 specparam_declaration_instance10749();
    specparam_declaration10750 specparam_declaration_instance10750();
    specparam_declaration10751 specparam_declaration_instance10751();
    specparam_declaration10752 specparam_declaration_instance10752();
    specparam_declaration10753 specparam_declaration_instance10753();
    specparam_declaration10754 specparam_declaration_instance10754();
    specparam_declaration10755 specparam_declaration_instance10755();
    specparam_declaration10756 specparam_declaration_instance10756();
    specparam_declaration10757 specparam_declaration_instance10757();
    specparam_declaration10758 specparam_declaration_instance10758();
    specparam_declaration10759 specparam_declaration_instance10759();
    specparam_declaration10760 specparam_declaration_instance10760();
    specparam_declaration10761 specparam_declaration_instance10761();
    specparam_declaration10762 specparam_declaration_instance10762();
    specparam_declaration10763 specparam_declaration_instance10763();
    specparam_declaration10764 specparam_declaration_instance10764();
    specparam_declaration10765 specparam_declaration_instance10765();
    specparam_declaration10766 specparam_declaration_instance10766();
    specparam_declaration10767 specparam_declaration_instance10767();
    specparam_declaration10768 specparam_declaration_instance10768();
    specparam_declaration10769 specparam_declaration_instance10769();
    specparam_declaration10770 specparam_declaration_instance10770();
    specparam_declaration10771 specparam_declaration_instance10771();
    specparam_declaration10772 specparam_declaration_instance10772();
    specparam_declaration10773 specparam_declaration_instance10773();
    specparam_declaration10774 specparam_declaration_instance10774();
    specparam_declaration10775 specparam_declaration_instance10775();
    specparam_declaration10776 specparam_declaration_instance10776();
    specparam_declaration10777 specparam_declaration_instance10777();
    specparam_declaration10778 specparam_declaration_instance10778();
    specparam_declaration10779 specparam_declaration_instance10779();
    specparam_declaration10780 specparam_declaration_instance10780();
    specparam_declaration10781 specparam_declaration_instance10781();
    specparam_declaration10782 specparam_declaration_instance10782();
    specparam_declaration10783 specparam_declaration_instance10783();
    specparam_declaration10784 specparam_declaration_instance10784();
    specparam_declaration10785 specparam_declaration_instance10785();
    specparam_declaration10786 specparam_declaration_instance10786();
    specparam_declaration10787 specparam_declaration_instance10787();
    specparam_declaration10788 specparam_declaration_instance10788();
    specparam_declaration10789 specparam_declaration_instance10789();
    specparam_declaration10790 specparam_declaration_instance10790();
    specparam_declaration10791 specparam_declaration_instance10791();
    specparam_declaration10792 specparam_declaration_instance10792();
    specparam_declaration10793 specparam_declaration_instance10793();
    specparam_declaration10794 specparam_declaration_instance10794();
    specparam_declaration10795 specparam_declaration_instance10795();
    specparam_declaration10796 specparam_declaration_instance10796();
    specparam_declaration10797 specparam_declaration_instance10797();
    specparam_declaration10798 specparam_declaration_instance10798();
    specparam_declaration10799 specparam_declaration_instance10799();
    specparam_declaration10800 specparam_declaration_instance10800();
    specparam_declaration10801 specparam_declaration_instance10801();
    specparam_declaration10802 specparam_declaration_instance10802();
    specparam_declaration10803 specparam_declaration_instance10803();
    specparam_declaration10804 specparam_declaration_instance10804();
    specparam_declaration10805 specparam_declaration_instance10805();
    specparam_declaration10806 specparam_declaration_instance10806();
    specparam_declaration10807 specparam_declaration_instance10807();
    specparam_declaration10808 specparam_declaration_instance10808();
    specparam_declaration10809 specparam_declaration_instance10809();
    specparam_declaration10810 specparam_declaration_instance10810();
    specparam_declaration10811 specparam_declaration_instance10811();
    specparam_declaration10812 specparam_declaration_instance10812();
    specparam_declaration10813 specparam_declaration_instance10813();
    specparam_declaration10814 specparam_declaration_instance10814();
    specparam_declaration10815 specparam_declaration_instance10815();
    specparam_declaration10816 specparam_declaration_instance10816();
    specparam_declaration10817 specparam_declaration_instance10817();
    specparam_declaration10818 specparam_declaration_instance10818();
    specparam_declaration10819 specparam_declaration_instance10819();
    specparam_declaration10820 specparam_declaration_instance10820();
    specparam_declaration10821 specparam_declaration_instance10821();
    specparam_declaration10822 specparam_declaration_instance10822();
    specparam_declaration10823 specparam_declaration_instance10823();
    specparam_declaration10824 specparam_declaration_instance10824();
    specparam_declaration10825 specparam_declaration_instance10825();
    specparam_declaration10826 specparam_declaration_instance10826();
    specparam_declaration10827 specparam_declaration_instance10827();
    specparam_declaration10828 specparam_declaration_instance10828();
    specparam_declaration10829 specparam_declaration_instance10829();
    specparam_declaration10830 specparam_declaration_instance10830();
    specparam_declaration10831 specparam_declaration_instance10831();
    specparam_declaration10832 specparam_declaration_instance10832();
    specparam_declaration10833 specparam_declaration_instance10833();
    specparam_declaration10834 specparam_declaration_instance10834();
    specparam_declaration10835 specparam_declaration_instance10835();
    specparam_declaration10836 specparam_declaration_instance10836();
    specparam_declaration10837 specparam_declaration_instance10837();
    specparam_declaration10838 specparam_declaration_instance10838();
    specparam_declaration10839 specparam_declaration_instance10839();
    specparam_declaration10840 specparam_declaration_instance10840();
    specparam_declaration10841 specparam_declaration_instance10841();
    specparam_declaration10842 specparam_declaration_instance10842();
    specparam_declaration10843 specparam_declaration_instance10843();
    specparam_declaration10844 specparam_declaration_instance10844();
    specparam_declaration10845 specparam_declaration_instance10845();
    specparam_declaration10846 specparam_declaration_instance10846();
    specparam_declaration10847 specparam_declaration_instance10847();
    specparam_declaration10848 specparam_declaration_instance10848();
    specparam_declaration10849 specparam_declaration_instance10849();
    specparam_declaration10850 specparam_declaration_instance10850();
    specparam_declaration10851 specparam_declaration_instance10851();
    specparam_declaration10852 specparam_declaration_instance10852();
    specparam_declaration10853 specparam_declaration_instance10853();
    specparam_declaration10854 specparam_declaration_instance10854();
    specparam_declaration10855 specparam_declaration_instance10855();
    specparam_declaration10856 specparam_declaration_instance10856();
    specparam_declaration10857 specparam_declaration_instance10857();
    specparam_declaration10858 specparam_declaration_instance10858();
    specparam_declaration10859 specparam_declaration_instance10859();
    specparam_declaration10860 specparam_declaration_instance10860();
    specparam_declaration10861 specparam_declaration_instance10861();
    specparam_declaration10862 specparam_declaration_instance10862();
    specparam_declaration10863 specparam_declaration_instance10863();
    specparam_declaration10864 specparam_declaration_instance10864();
    specparam_declaration10865 specparam_declaration_instance10865();
    specparam_declaration10866 specparam_declaration_instance10866();
    specparam_declaration10867 specparam_declaration_instance10867();
    specparam_declaration10868 specparam_declaration_instance10868();
    specparam_declaration10869 specparam_declaration_instance10869();
    specparam_declaration10870 specparam_declaration_instance10870();
    specparam_declaration10871 specparam_declaration_instance10871();
    specparam_declaration10872 specparam_declaration_instance10872();
    specparam_declaration10873 specparam_declaration_instance10873();
    specparam_declaration10874 specparam_declaration_instance10874();
    specparam_declaration10875 specparam_declaration_instance10875();
    specparam_declaration10876 specparam_declaration_instance10876();
    specparam_declaration10877 specparam_declaration_instance10877();
    specparam_declaration10878 specparam_declaration_instance10878();
    specparam_declaration10879 specparam_declaration_instance10879();
    specparam_declaration10880 specparam_declaration_instance10880();
    specparam_declaration10881 specparam_declaration_instance10881();
    specparam_declaration10882 specparam_declaration_instance10882();
    specparam_declaration10883 specparam_declaration_instance10883();
    specparam_declaration10884 specparam_declaration_instance10884();
    specparam_declaration10885 specparam_declaration_instance10885();
    specparam_declaration10886 specparam_declaration_instance10886();
    specparam_declaration10887 specparam_declaration_instance10887();
    specparam_declaration10888 specparam_declaration_instance10888();
    specparam_declaration10889 specparam_declaration_instance10889();
    specparam_declaration10890 specparam_declaration_instance10890();
    specparam_declaration10891 specparam_declaration_instance10891();
    specparam_declaration10892 specparam_declaration_instance10892();
    specparam_declaration10893 specparam_declaration_instance10893();
    specparam_declaration10894 specparam_declaration_instance10894();
    specparam_declaration10895 specparam_declaration_instance10895();
    specparam_declaration10896 specparam_declaration_instance10896();
    specparam_declaration10897 specparam_declaration_instance10897();
    specparam_declaration10898 specparam_declaration_instance10898();
    specparam_declaration10899 specparam_declaration_instance10899();
    specparam_declaration10900 specparam_declaration_instance10900();
    specparam_declaration10901 specparam_declaration_instance10901();
    specparam_declaration10902 specparam_declaration_instance10902();
    specparam_declaration10903 specparam_declaration_instance10903();
    specparam_declaration10904 specparam_declaration_instance10904();
    specparam_declaration10905 specparam_declaration_instance10905();
    specparam_declaration10906 specparam_declaration_instance10906();
    specparam_declaration10907 specparam_declaration_instance10907();
    specparam_declaration10908 specparam_declaration_instance10908();
    specparam_declaration10909 specparam_declaration_instance10909();
    specparam_declaration10910 specparam_declaration_instance10910();
    specparam_declaration10911 specparam_declaration_instance10911();
    specparam_declaration10912 specparam_declaration_instance10912();
    specparam_declaration10913 specparam_declaration_instance10913();
    specparam_declaration10914 specparam_declaration_instance10914();
    specparam_declaration10915 specparam_declaration_instance10915();
    specparam_declaration10916 specparam_declaration_instance10916();
    specparam_declaration10917 specparam_declaration_instance10917();
    specparam_declaration10918 specparam_declaration_instance10918();
    specparam_declaration10919 specparam_declaration_instance10919();
    specparam_declaration10920 specparam_declaration_instance10920();
    specparam_declaration10921 specparam_declaration_instance10921();
    specparam_declaration10922 specparam_declaration_instance10922();
    specparam_declaration10923 specparam_declaration_instance10923();
    specparam_declaration10924 specparam_declaration_instance10924();
    specparam_declaration10925 specparam_declaration_instance10925();
    specparam_declaration10926 specparam_declaration_instance10926();
    specparam_declaration10927 specparam_declaration_instance10927();
    specparam_declaration10928 specparam_declaration_instance10928();
    specparam_declaration10929 specparam_declaration_instance10929();
    specparam_declaration10930 specparam_declaration_instance10930();
    specparam_declaration10931 specparam_declaration_instance10931();
    specparam_declaration10932 specparam_declaration_instance10932();
    specparam_declaration10933 specparam_declaration_instance10933();
    specparam_declaration10934 specparam_declaration_instance10934();
    specparam_declaration10935 specparam_declaration_instance10935();
    specparam_declaration10936 specparam_declaration_instance10936();
    specparam_declaration10937 specparam_declaration_instance10937();
    specparam_declaration10938 specparam_declaration_instance10938();
    specparam_declaration10939 specparam_declaration_instance10939();
    specparam_declaration10940 specparam_declaration_instance10940();
    specparam_declaration10941 specparam_declaration_instance10941();
    specparam_declaration10942 specparam_declaration_instance10942();
    specparam_declaration10943 specparam_declaration_instance10943();
    specparam_declaration10944 specparam_declaration_instance10944();
    specparam_declaration10945 specparam_declaration_instance10945();
    specparam_declaration10946 specparam_declaration_instance10946();
    specparam_declaration10947 specparam_declaration_instance10947();
    specparam_declaration10948 specparam_declaration_instance10948();
    specparam_declaration10949 specparam_declaration_instance10949();
    specparam_declaration10950 specparam_declaration_instance10950();
    specparam_declaration10951 specparam_declaration_instance10951();
    specparam_declaration10952 specparam_declaration_instance10952();
    specparam_declaration10953 specparam_declaration_instance10953();
    specparam_declaration10954 specparam_declaration_instance10954();
    specparam_declaration10955 specparam_declaration_instance10955();
    specparam_declaration10956 specparam_declaration_instance10956();
    specparam_declaration10957 specparam_declaration_instance10957();
    specparam_declaration10958 specparam_declaration_instance10958();
    specparam_declaration10959 specparam_declaration_instance10959();
    specparam_declaration10960 specparam_declaration_instance10960();
    specparam_declaration10961 specparam_declaration_instance10961();
    specparam_declaration10962 specparam_declaration_instance10962();
    specparam_declaration10963 specparam_declaration_instance10963();
    specparam_declaration10964 specparam_declaration_instance10964();
    specparam_declaration10965 specparam_declaration_instance10965();
    specparam_declaration10966 specparam_declaration_instance10966();
    specparam_declaration10967 specparam_declaration_instance10967();
    specparam_declaration10968 specparam_declaration_instance10968();
    specparam_declaration10969 specparam_declaration_instance10969();
    specparam_declaration10970 specparam_declaration_instance10970();
    specparam_declaration10971 specparam_declaration_instance10971();
    specparam_declaration10972 specparam_declaration_instance10972();
    specparam_declaration10973 specparam_declaration_instance10973();
    specparam_declaration10974 specparam_declaration_instance10974();
    specparam_declaration10975 specparam_declaration_instance10975();
    specparam_declaration10976 specparam_declaration_instance10976();
    specparam_declaration10977 specparam_declaration_instance10977();
    specparam_declaration10978 specparam_declaration_instance10978();
    specparam_declaration10979 specparam_declaration_instance10979();
    specparam_declaration10980 specparam_declaration_instance10980();
    specparam_declaration10981 specparam_declaration_instance10981();
    specparam_declaration10982 specparam_declaration_instance10982();
    specparam_declaration10983 specparam_declaration_instance10983();
    specparam_declaration10984 specparam_declaration_instance10984();
    specparam_declaration10985 specparam_declaration_instance10985();
    specparam_declaration10986 specparam_declaration_instance10986();
    specparam_declaration10987 specparam_declaration_instance10987();
    specparam_declaration10988 specparam_declaration_instance10988();
    specparam_declaration10989 specparam_declaration_instance10989();
    specparam_declaration10990 specparam_declaration_instance10990();
    specparam_declaration10991 specparam_declaration_instance10991();
    specparam_declaration10992 specparam_declaration_instance10992();
    specparam_declaration10993 specparam_declaration_instance10993();
    specparam_declaration10994 specparam_declaration_instance10994();
    specparam_declaration10995 specparam_declaration_instance10995();
    specparam_declaration10996 specparam_declaration_instance10996();
    specparam_declaration10997 specparam_declaration_instance10997();
    specparam_declaration10998 specparam_declaration_instance10998();
    specparam_declaration10999 specparam_declaration_instance10999();
    specparam_declaration11000 specparam_declaration_instance11000();
    specparam_declaration11001 specparam_declaration_instance11001();
    specparam_declaration11002 specparam_declaration_instance11002();
    specparam_declaration11003 specparam_declaration_instance11003();
    specparam_declaration11004 specparam_declaration_instance11004();
    specparam_declaration11005 specparam_declaration_instance11005();
    specparam_declaration11006 specparam_declaration_instance11006();
    specparam_declaration11007 specparam_declaration_instance11007();
    specparam_declaration11008 specparam_declaration_instance11008();
    specparam_declaration11009 specparam_declaration_instance11009();
    specparam_declaration11010 specparam_declaration_instance11010();
    specparam_declaration11011 specparam_declaration_instance11011();
    specparam_declaration11012 specparam_declaration_instance11012();
    specparam_declaration11013 specparam_declaration_instance11013();
    specparam_declaration11014 specparam_declaration_instance11014();
    specparam_declaration11015 specparam_declaration_instance11015();
    specparam_declaration11016 specparam_declaration_instance11016();
    specparam_declaration11017 specparam_declaration_instance11017();
    specparam_declaration11018 specparam_declaration_instance11018();
    specparam_declaration11019 specparam_declaration_instance11019();
    specparam_declaration11020 specparam_declaration_instance11020();
    specparam_declaration11021 specparam_declaration_instance11021();
    specparam_declaration11022 specparam_declaration_instance11022();
    specparam_declaration11023 specparam_declaration_instance11023();
    specparam_declaration11024 specparam_declaration_instance11024();
    specparam_declaration11025 specparam_declaration_instance11025();
    specparam_declaration11026 specparam_declaration_instance11026();
    specparam_declaration11027 specparam_declaration_instance11027();
    specparam_declaration11028 specparam_declaration_instance11028();
    specparam_declaration11029 specparam_declaration_instance11029();
    specparam_declaration11030 specparam_declaration_instance11030();
    specparam_declaration11031 specparam_declaration_instance11031();
    specparam_declaration11032 specparam_declaration_instance11032();
    specparam_declaration11033 specparam_declaration_instance11033();
    specparam_declaration11034 specparam_declaration_instance11034();
    specparam_declaration11035 specparam_declaration_instance11035();
    specparam_declaration11036 specparam_declaration_instance11036();
    specparam_declaration11037 specparam_declaration_instance11037();
    specparam_declaration11038 specparam_declaration_instance11038();
    specparam_declaration11039 specparam_declaration_instance11039();
    specparam_declaration11040 specparam_declaration_instance11040();
    specparam_declaration11041 specparam_declaration_instance11041();
    specparam_declaration11042 specparam_declaration_instance11042();
    specparam_declaration11043 specparam_declaration_instance11043();
    specparam_declaration11044 specparam_declaration_instance11044();
    specparam_declaration11045 specparam_declaration_instance11045();
    specparam_declaration11046 specparam_declaration_instance11046();
    specparam_declaration11047 specparam_declaration_instance11047();
    specparam_declaration11048 specparam_declaration_instance11048();
    specparam_declaration11049 specparam_declaration_instance11049();
    specparam_declaration11050 specparam_declaration_instance11050();
    specparam_declaration11051 specparam_declaration_instance11051();
    specparam_declaration11052 specparam_declaration_instance11052();
    specparam_declaration11053 specparam_declaration_instance11053();
    specparam_declaration11054 specparam_declaration_instance11054();
    specparam_declaration11055 specparam_declaration_instance11055();
    specparam_declaration11056 specparam_declaration_instance11056();
    specparam_declaration11057 specparam_declaration_instance11057();
    specparam_declaration11058 specparam_declaration_instance11058();
    specparam_declaration11059 specparam_declaration_instance11059();
    specparam_declaration11060 specparam_declaration_instance11060();
    specparam_declaration11061 specparam_declaration_instance11061();
    specparam_declaration11062 specparam_declaration_instance11062();
    specparam_declaration11063 specparam_declaration_instance11063();
    specparam_declaration11064 specparam_declaration_instance11064();
    specparam_declaration11065 specparam_declaration_instance11065();
    specparam_declaration11066 specparam_declaration_instance11066();
    specparam_declaration11067 specparam_declaration_instance11067();
    specparam_declaration11068 specparam_declaration_instance11068();
    specparam_declaration11069 specparam_declaration_instance11069();
    specparam_declaration11070 specparam_declaration_instance11070();
    specparam_declaration11071 specparam_declaration_instance11071();
    specparam_declaration11072 specparam_declaration_instance11072();
    specparam_declaration11073 specparam_declaration_instance11073();
    specparam_declaration11074 specparam_declaration_instance11074();
    specparam_declaration11075 specparam_declaration_instance11075();
    specparam_declaration11076 specparam_declaration_instance11076();
    specparam_declaration11077 specparam_declaration_instance11077();
    specparam_declaration11078 specparam_declaration_instance11078();
    specparam_declaration11079 specparam_declaration_instance11079();
    specparam_declaration11080 specparam_declaration_instance11080();
    specparam_declaration11081 specparam_declaration_instance11081();
    specparam_declaration11082 specparam_declaration_instance11082();
    specparam_declaration11083 specparam_declaration_instance11083();
    specparam_declaration11084 specparam_declaration_instance11084();
    specparam_declaration11085 specparam_declaration_instance11085();
    specparam_declaration11086 specparam_declaration_instance11086();
    specparam_declaration11087 specparam_declaration_instance11087();
    specparam_declaration11088 specparam_declaration_instance11088();
    specparam_declaration11089 specparam_declaration_instance11089();
    specparam_declaration11090 specparam_declaration_instance11090();
    specparam_declaration11091 specparam_declaration_instance11091();
    specparam_declaration11092 specparam_declaration_instance11092();
    specparam_declaration11093 specparam_declaration_instance11093();
    specparam_declaration11094 specparam_declaration_instance11094();
    specparam_declaration11095 specparam_declaration_instance11095();
    specparam_declaration11096 specparam_declaration_instance11096();
    specparam_declaration11097 specparam_declaration_instance11097();
    specparam_declaration11098 specparam_declaration_instance11098();
    specparam_declaration11099 specparam_declaration_instance11099();
    specparam_declaration11100 specparam_declaration_instance11100();
    specparam_declaration11101 specparam_declaration_instance11101();
    specparam_declaration11102 specparam_declaration_instance11102();
    specparam_declaration11103 specparam_declaration_instance11103();
    specparam_declaration11104 specparam_declaration_instance11104();
    specparam_declaration11105 specparam_declaration_instance11105();
    specparam_declaration11106 specparam_declaration_instance11106();
    specparam_declaration11107 specparam_declaration_instance11107();
    specparam_declaration11108 specparam_declaration_instance11108();
    specparam_declaration11109 specparam_declaration_instance11109();
    specparam_declaration11110 specparam_declaration_instance11110();
    specparam_declaration11111 specparam_declaration_instance11111();
    specparam_declaration11112 specparam_declaration_instance11112();
    specparam_declaration11113 specparam_declaration_instance11113();
    specparam_declaration11114 specparam_declaration_instance11114();
    specparam_declaration11115 specparam_declaration_instance11115();
    specparam_declaration11116 specparam_declaration_instance11116();
    specparam_declaration11117 specparam_declaration_instance11117();
    specparam_declaration11118 specparam_declaration_instance11118();
    specparam_declaration11119 specparam_declaration_instance11119();
    specparam_declaration11120 specparam_declaration_instance11120();
    specparam_declaration11121 specparam_declaration_instance11121();
    specparam_declaration11122 specparam_declaration_instance11122();
    specparam_declaration11123 specparam_declaration_instance11123();
    specparam_declaration11124 specparam_declaration_instance11124();
    specparam_declaration11125 specparam_declaration_instance11125();
    specparam_declaration11126 specparam_declaration_instance11126();
    specparam_declaration11127 specparam_declaration_instance11127();
    specparam_declaration11128 specparam_declaration_instance11128();
    specparam_declaration11129 specparam_declaration_instance11129();
    specparam_declaration11130 specparam_declaration_instance11130();
    specparam_declaration11131 specparam_declaration_instance11131();
    specparam_declaration11132 specparam_declaration_instance11132();
    specparam_declaration11133 specparam_declaration_instance11133();
    specparam_declaration11134 specparam_declaration_instance11134();
    specparam_declaration11135 specparam_declaration_instance11135();
    specparam_declaration11136 specparam_declaration_instance11136();
    specparam_declaration11137 specparam_declaration_instance11137();
    specparam_declaration11138 specparam_declaration_instance11138();
    specparam_declaration11139 specparam_declaration_instance11139();
    specparam_declaration11140 specparam_declaration_instance11140();
    specparam_declaration11141 specparam_declaration_instance11141();
    specparam_declaration11142 specparam_declaration_instance11142();
    specparam_declaration11143 specparam_declaration_instance11143();
    specparam_declaration11144 specparam_declaration_instance11144();
    specparam_declaration11145 specparam_declaration_instance11145();
    specparam_declaration11146 specparam_declaration_instance11146();
    specparam_declaration11147 specparam_declaration_instance11147();
    specparam_declaration11148 specparam_declaration_instance11148();
    specparam_declaration11149 specparam_declaration_instance11149();
    specparam_declaration11150 specparam_declaration_instance11150();
    specparam_declaration11151 specparam_declaration_instance11151();
    specparam_declaration11152 specparam_declaration_instance11152();
    specparam_declaration11153 specparam_declaration_instance11153();
    specparam_declaration11154 specparam_declaration_instance11154();
    specparam_declaration11155 specparam_declaration_instance11155();
    specparam_declaration11156 specparam_declaration_instance11156();
    specparam_declaration11157 specparam_declaration_instance11157();
    specparam_declaration11158 specparam_declaration_instance11158();
    specparam_declaration11159 specparam_declaration_instance11159();
    specparam_declaration11160 specparam_declaration_instance11160();
    specparam_declaration11161 specparam_declaration_instance11161();
    specparam_declaration11162 specparam_declaration_instance11162();
    specparam_declaration11163 specparam_declaration_instance11163();
    specparam_declaration11164 specparam_declaration_instance11164();
    specparam_declaration11165 specparam_declaration_instance11165();
    specparam_declaration11166 specparam_declaration_instance11166();
    specparam_declaration11167 specparam_declaration_instance11167();
    specparam_declaration11168 specparam_declaration_instance11168();
    specparam_declaration11169 specparam_declaration_instance11169();
    specparam_declaration11170 specparam_declaration_instance11170();
    specparam_declaration11171 specparam_declaration_instance11171();
    specparam_declaration11172 specparam_declaration_instance11172();
    specparam_declaration11173 specparam_declaration_instance11173();
    specparam_declaration11174 specparam_declaration_instance11174();
    specparam_declaration11175 specparam_declaration_instance11175();
    specparam_declaration11176 specparam_declaration_instance11176();
    specparam_declaration11177 specparam_declaration_instance11177();
    specparam_declaration11178 specparam_declaration_instance11178();
    specparam_declaration11179 specparam_declaration_instance11179();
    specparam_declaration11180 specparam_declaration_instance11180();
    specparam_declaration11181 specparam_declaration_instance11181();
    specparam_declaration11182 specparam_declaration_instance11182();
    specparam_declaration11183 specparam_declaration_instance11183();
    specparam_declaration11184 specparam_declaration_instance11184();
    specparam_declaration11185 specparam_declaration_instance11185();
    specparam_declaration11186 specparam_declaration_instance11186();
    specparam_declaration11187 specparam_declaration_instance11187();
    specparam_declaration11188 specparam_declaration_instance11188();
    specparam_declaration11189 specparam_declaration_instance11189();
    specparam_declaration11190 specparam_declaration_instance11190();
    specparam_declaration11191 specparam_declaration_instance11191();
    specparam_declaration11192 specparam_declaration_instance11192();
    specparam_declaration11193 specparam_declaration_instance11193();
    specparam_declaration11194 specparam_declaration_instance11194();
    specparam_declaration11195 specparam_declaration_instance11195();
    specparam_declaration11196 specparam_declaration_instance11196();
    specparam_declaration11197 specparam_declaration_instance11197();
    specparam_declaration11198 specparam_declaration_instance11198();
    specparam_declaration11199 specparam_declaration_instance11199();
    specparam_declaration11200 specparam_declaration_instance11200();
    specparam_declaration11201 specparam_declaration_instance11201();
    specparam_declaration11202 specparam_declaration_instance11202();
    specparam_declaration11203 specparam_declaration_instance11203();
    specparam_declaration11204 specparam_declaration_instance11204();
    specparam_declaration11205 specparam_declaration_instance11205();
    specparam_declaration11206 specparam_declaration_instance11206();
    specparam_declaration11207 specparam_declaration_instance11207();
    specparam_declaration11208 specparam_declaration_instance11208();
    specparam_declaration11209 specparam_declaration_instance11209();
    specparam_declaration11210 specparam_declaration_instance11210();
    specparam_declaration11211 specparam_declaration_instance11211();
    specparam_declaration11212 specparam_declaration_instance11212();
    specparam_declaration11213 specparam_declaration_instance11213();
    specparam_declaration11214 specparam_declaration_instance11214();
    specparam_declaration11215 specparam_declaration_instance11215();
    specparam_declaration11216 specparam_declaration_instance11216();
    specparam_declaration11217 specparam_declaration_instance11217();
    specparam_declaration11218 specparam_declaration_instance11218();
    specparam_declaration11219 specparam_declaration_instance11219();
    specparam_declaration11220 specparam_declaration_instance11220();
    specparam_declaration11221 specparam_declaration_instance11221();
    specparam_declaration11222 specparam_declaration_instance11222();
    specparam_declaration11223 specparam_declaration_instance11223();
    specparam_declaration11224 specparam_declaration_instance11224();
    specparam_declaration11225 specparam_declaration_instance11225();
    specparam_declaration11226 specparam_declaration_instance11226();
    specparam_declaration11227 specparam_declaration_instance11227();
    specparam_declaration11228 specparam_declaration_instance11228();
    specparam_declaration11229 specparam_declaration_instance11229();
    specparam_declaration11230 specparam_declaration_instance11230();
    specparam_declaration11231 specparam_declaration_instance11231();
    specparam_declaration11232 specparam_declaration_instance11232();
    specparam_declaration11233 specparam_declaration_instance11233();
    specparam_declaration11234 specparam_declaration_instance11234();
    specparam_declaration11235 specparam_declaration_instance11235();
    specparam_declaration11236 specparam_declaration_instance11236();
    specparam_declaration11237 specparam_declaration_instance11237();
    specparam_declaration11238 specparam_declaration_instance11238();
    specparam_declaration11239 specparam_declaration_instance11239();
    specparam_declaration11240 specparam_declaration_instance11240();
    specparam_declaration11241 specparam_declaration_instance11241();
    specparam_declaration11242 specparam_declaration_instance11242();
    specparam_declaration11243 specparam_declaration_instance11243();
    specparam_declaration11244 specparam_declaration_instance11244();
    specparam_declaration11245 specparam_declaration_instance11245();
    specparam_declaration11246 specparam_declaration_instance11246();
    specparam_declaration11247 specparam_declaration_instance11247();
    specparam_declaration11248 specparam_declaration_instance11248();
    specparam_declaration11249 specparam_declaration_instance11249();
    specparam_declaration11250 specparam_declaration_instance11250();
    specparam_declaration11251 specparam_declaration_instance11251();
    specparam_declaration11252 specparam_declaration_instance11252();
    specparam_declaration11253 specparam_declaration_instance11253();
    specparam_declaration11254 specparam_declaration_instance11254();
    specparam_declaration11255 specparam_declaration_instance11255();
    specparam_declaration11256 specparam_declaration_instance11256();
    specparam_declaration11257 specparam_declaration_instance11257();
    specparam_declaration11258 specparam_declaration_instance11258();
    specparam_declaration11259 specparam_declaration_instance11259();
    specparam_declaration11260 specparam_declaration_instance11260();
    specparam_declaration11261 specparam_declaration_instance11261();
    specparam_declaration11262 specparam_declaration_instance11262();
    specparam_declaration11263 specparam_declaration_instance11263();
    specparam_declaration11264 specparam_declaration_instance11264();
    specparam_declaration11265 specparam_declaration_instance11265();
    specparam_declaration11266 specparam_declaration_instance11266();
    specparam_declaration11267 specparam_declaration_instance11267();
    specparam_declaration11268 specparam_declaration_instance11268();
    specparam_declaration11269 specparam_declaration_instance11269();
    specparam_declaration11270 specparam_declaration_instance11270();
    specparam_declaration11271 specparam_declaration_instance11271();
    specparam_declaration11272 specparam_declaration_instance11272();
    specparam_declaration11273 specparam_declaration_instance11273();
    specparam_declaration11274 specparam_declaration_instance11274();
    specparam_declaration11275 specparam_declaration_instance11275();
    specparam_declaration11276 specparam_declaration_instance11276();
    specparam_declaration11277 specparam_declaration_instance11277();
    specparam_declaration11278 specparam_declaration_instance11278();
    specparam_declaration11279 specparam_declaration_instance11279();
    specparam_declaration11280 specparam_declaration_instance11280();
    specparam_declaration11281 specparam_declaration_instance11281();
    specparam_declaration11282 specparam_declaration_instance11282();
    specparam_declaration11283 specparam_declaration_instance11283();
    specparam_declaration11284 specparam_declaration_instance11284();
    specparam_declaration11285 specparam_declaration_instance11285();
    specparam_declaration11286 specparam_declaration_instance11286();
    specparam_declaration11287 specparam_declaration_instance11287();
    specparam_declaration11288 specparam_declaration_instance11288();
    specparam_declaration11289 specparam_declaration_instance11289();
    specparam_declaration11290 specparam_declaration_instance11290();
    specparam_declaration11291 specparam_declaration_instance11291();
    specparam_declaration11292 specparam_declaration_instance11292();
    specparam_declaration11293 specparam_declaration_instance11293();
    specparam_declaration11294 specparam_declaration_instance11294();
    specparam_declaration11295 specparam_declaration_instance11295();
    specparam_declaration11296 specparam_declaration_instance11296();
    specparam_declaration11297 specparam_declaration_instance11297();
    specparam_declaration11298 specparam_declaration_instance11298();
    specparam_declaration11299 specparam_declaration_instance11299();
    specparam_declaration11300 specparam_declaration_instance11300();
    specparam_declaration11301 specparam_declaration_instance11301();
    specparam_declaration11302 specparam_declaration_instance11302();
    specparam_declaration11303 specparam_declaration_instance11303();
    specparam_declaration11304 specparam_declaration_instance11304();
    specparam_declaration11305 specparam_declaration_instance11305();
    specparam_declaration11306 specparam_declaration_instance11306();
    specparam_declaration11307 specparam_declaration_instance11307();
    specparam_declaration11308 specparam_declaration_instance11308();
    specparam_declaration11309 specparam_declaration_instance11309();
    specparam_declaration11310 specparam_declaration_instance11310();
    specparam_declaration11311 specparam_declaration_instance11311();
    specparam_declaration11312 specparam_declaration_instance11312();
    specparam_declaration11313 specparam_declaration_instance11313();
    specparam_declaration11314 specparam_declaration_instance11314();
    specparam_declaration11315 specparam_declaration_instance11315();
    specparam_declaration11316 specparam_declaration_instance11316();
    specparam_declaration11317 specparam_declaration_instance11317();
    specparam_declaration11318 specparam_declaration_instance11318();
    specparam_declaration11319 specparam_declaration_instance11319();
    specparam_declaration11320 specparam_declaration_instance11320();
    specparam_declaration11321 specparam_declaration_instance11321();
    specparam_declaration11322 specparam_declaration_instance11322();
    specparam_declaration11323 specparam_declaration_instance11323();
    specparam_declaration11324 specparam_declaration_instance11324();
    specparam_declaration11325 specparam_declaration_instance11325();
    specparam_declaration11326 specparam_declaration_instance11326();
    specparam_declaration11327 specparam_declaration_instance11327();
    specparam_declaration11328 specparam_declaration_instance11328();
    specparam_declaration11329 specparam_declaration_instance11329();
    specparam_declaration11330 specparam_declaration_instance11330();
    specparam_declaration11331 specparam_declaration_instance11331();
    specparam_declaration11332 specparam_declaration_instance11332();
    specparam_declaration11333 specparam_declaration_instance11333();
    specparam_declaration11334 specparam_declaration_instance11334();
    specparam_declaration11335 specparam_declaration_instance11335();
    specparam_declaration11336 specparam_declaration_instance11336();
    specparam_declaration11337 specparam_declaration_instance11337();
    specparam_declaration11338 specparam_declaration_instance11338();
    specparam_declaration11339 specparam_declaration_instance11339();
    specparam_declaration11340 specparam_declaration_instance11340();
    specparam_declaration11341 specparam_declaration_instance11341();
    specparam_declaration11342 specparam_declaration_instance11342();
    specparam_declaration11343 specparam_declaration_instance11343();
    specparam_declaration11344 specparam_declaration_instance11344();
    specparam_declaration11345 specparam_declaration_instance11345();
    specparam_declaration11346 specparam_declaration_instance11346();
    specparam_declaration11347 specparam_declaration_instance11347();
    specparam_declaration11348 specparam_declaration_instance11348();
    specparam_declaration11349 specparam_declaration_instance11349();
    specparam_declaration11350 specparam_declaration_instance11350();
    specparam_declaration11351 specparam_declaration_instance11351();
    specparam_declaration11352 specparam_declaration_instance11352();
    specparam_declaration11353 specparam_declaration_instance11353();
    specparam_declaration11354 specparam_declaration_instance11354();
    specparam_declaration11355 specparam_declaration_instance11355();
    specparam_declaration11356 specparam_declaration_instance11356();
    specparam_declaration11357 specparam_declaration_instance11357();
    specparam_declaration11358 specparam_declaration_instance11358();
    specparam_declaration11359 specparam_declaration_instance11359();
    specparam_declaration11360 specparam_declaration_instance11360();
    specparam_declaration11361 specparam_declaration_instance11361();
    specparam_declaration11362 specparam_declaration_instance11362();
    specparam_declaration11363 specparam_declaration_instance11363();
    specparam_declaration11364 specparam_declaration_instance11364();
    specparam_declaration11365 specparam_declaration_instance11365();
    specparam_declaration11366 specparam_declaration_instance11366();
    specparam_declaration11367 specparam_declaration_instance11367();
    specparam_declaration11368 specparam_declaration_instance11368();
    specparam_declaration11369 specparam_declaration_instance11369();
    specparam_declaration11370 specparam_declaration_instance11370();
    specparam_declaration11371 specparam_declaration_instance11371();
    specparam_declaration11372 specparam_declaration_instance11372();
    specparam_declaration11373 specparam_declaration_instance11373();
    specparam_declaration11374 specparam_declaration_instance11374();
    specparam_declaration11375 specparam_declaration_instance11375();
    specparam_declaration11376 specparam_declaration_instance11376();
    specparam_declaration11377 specparam_declaration_instance11377();
    specparam_declaration11378 specparam_declaration_instance11378();
    specparam_declaration11379 specparam_declaration_instance11379();
    specparam_declaration11380 specparam_declaration_instance11380();
    specparam_declaration11381 specparam_declaration_instance11381();
    specparam_declaration11382 specparam_declaration_instance11382();
    specparam_declaration11383 specparam_declaration_instance11383();
    specparam_declaration11384 specparam_declaration_instance11384();
    specparam_declaration11385 specparam_declaration_instance11385();
    specparam_declaration11386 specparam_declaration_instance11386();
    specparam_declaration11387 specparam_declaration_instance11387();
    specparam_declaration11388 specparam_declaration_instance11388();
    specparam_declaration11389 specparam_declaration_instance11389();
    specparam_declaration11390 specparam_declaration_instance11390();
    specparam_declaration11391 specparam_declaration_instance11391();
    specparam_declaration11392 specparam_declaration_instance11392();
    specparam_declaration11393 specparam_declaration_instance11393();
    specparam_declaration11394 specparam_declaration_instance11394();
    specparam_declaration11395 specparam_declaration_instance11395();
    specparam_declaration11396 specparam_declaration_instance11396();
    specparam_declaration11397 specparam_declaration_instance11397();
    specparam_declaration11398 specparam_declaration_instance11398();
    specparam_declaration11399 specparam_declaration_instance11399();
    specparam_declaration11400 specparam_declaration_instance11400();
    specparam_declaration11401 specparam_declaration_instance11401();
    specparam_declaration11402 specparam_declaration_instance11402();
    specparam_declaration11403 specparam_declaration_instance11403();
    specparam_declaration11404 specparam_declaration_instance11404();
    specparam_declaration11405 specparam_declaration_instance11405();
    specparam_declaration11406 specparam_declaration_instance11406();
    specparam_declaration11407 specparam_declaration_instance11407();
    specparam_declaration11408 specparam_declaration_instance11408();
    specparam_declaration11409 specparam_declaration_instance11409();
    specparam_declaration11410 specparam_declaration_instance11410();
    specparam_declaration11411 specparam_declaration_instance11411();
    specparam_declaration11412 specparam_declaration_instance11412();
    specparam_declaration11413 specparam_declaration_instance11413();
    specparam_declaration11414 specparam_declaration_instance11414();
    specparam_declaration11415 specparam_declaration_instance11415();
    specparam_declaration11416 specparam_declaration_instance11416();
    specparam_declaration11417 specparam_declaration_instance11417();
    specparam_declaration11418 specparam_declaration_instance11418();
    specparam_declaration11419 specparam_declaration_instance11419();
    specparam_declaration11420 specparam_declaration_instance11420();
    specparam_declaration11421 specparam_declaration_instance11421();
    specparam_declaration11422 specparam_declaration_instance11422();
    specparam_declaration11423 specparam_declaration_instance11423();
    specparam_declaration11424 specparam_declaration_instance11424();
    specparam_declaration11425 specparam_declaration_instance11425();
    specparam_declaration11426 specparam_declaration_instance11426();
    specparam_declaration11427 specparam_declaration_instance11427();
    specparam_declaration11428 specparam_declaration_instance11428();
    specparam_declaration11429 specparam_declaration_instance11429();
    specparam_declaration11430 specparam_declaration_instance11430();
    specparam_declaration11431 specparam_declaration_instance11431();
    specparam_declaration11432 specparam_declaration_instance11432();
    specparam_declaration11433 specparam_declaration_instance11433();
    specparam_declaration11434 specparam_declaration_instance11434();
    specparam_declaration11435 specparam_declaration_instance11435();
    specparam_declaration11436 specparam_declaration_instance11436();
    specparam_declaration11437 specparam_declaration_instance11437();
    specparam_declaration11438 specparam_declaration_instance11438();
    specparam_declaration11439 specparam_declaration_instance11439();
    specparam_declaration11440 specparam_declaration_instance11440();
    specparam_declaration11441 specparam_declaration_instance11441();
    specparam_declaration11442 specparam_declaration_instance11442();
    specparam_declaration11443 specparam_declaration_instance11443();
    specparam_declaration11444 specparam_declaration_instance11444();
    specparam_declaration11445 specparam_declaration_instance11445();
    specparam_declaration11446 specparam_declaration_instance11446();
    specparam_declaration11447 specparam_declaration_instance11447();
    specparam_declaration11448 specparam_declaration_instance11448();
    specparam_declaration11449 specparam_declaration_instance11449();
    specparam_declaration11450 specparam_declaration_instance11450();
    specparam_declaration11451 specparam_declaration_instance11451();
    specparam_declaration11452 specparam_declaration_instance11452();
    specparam_declaration11453 specparam_declaration_instance11453();
    specparam_declaration11454 specparam_declaration_instance11454();
    specparam_declaration11455 specparam_declaration_instance11455();
    specparam_declaration11456 specparam_declaration_instance11456();
    specparam_declaration11457 specparam_declaration_instance11457();
    specparam_declaration11458 specparam_declaration_instance11458();
    specparam_declaration11459 specparam_declaration_instance11459();
    specparam_declaration11460 specparam_declaration_instance11460();
    specparam_declaration11461 specparam_declaration_instance11461();
    specparam_declaration11462 specparam_declaration_instance11462();
    specparam_declaration11463 specparam_declaration_instance11463();
    specparam_declaration11464 specparam_declaration_instance11464();
    specparam_declaration11465 specparam_declaration_instance11465();
    specparam_declaration11466 specparam_declaration_instance11466();
    specparam_declaration11467 specparam_declaration_instance11467();
    specparam_declaration11468 specparam_declaration_instance11468();
    specparam_declaration11469 specparam_declaration_instance11469();
    specparam_declaration11470 specparam_declaration_instance11470();
    specparam_declaration11471 specparam_declaration_instance11471();
    specparam_declaration11472 specparam_declaration_instance11472();
    specparam_declaration11473 specparam_declaration_instance11473();
    specparam_declaration11474 specparam_declaration_instance11474();
    specparam_declaration11475 specparam_declaration_instance11475();
    specparam_declaration11476 specparam_declaration_instance11476();
    specparam_declaration11477 specparam_declaration_instance11477();
    specparam_declaration11478 specparam_declaration_instance11478();
    specparam_declaration11479 specparam_declaration_instance11479();
    specparam_declaration11480 specparam_declaration_instance11480();
    specparam_declaration11481 specparam_declaration_instance11481();
    specparam_declaration11482 specparam_declaration_instance11482();
    specparam_declaration11483 specparam_declaration_instance11483();
    specparam_declaration11484 specparam_declaration_instance11484();
    specparam_declaration11485 specparam_declaration_instance11485();
    specparam_declaration11486 specparam_declaration_instance11486();
    specparam_declaration11487 specparam_declaration_instance11487();
    specparam_declaration11488 specparam_declaration_instance11488();
    specparam_declaration11489 specparam_declaration_instance11489();
    specparam_declaration11490 specparam_declaration_instance11490();
    specparam_declaration11491 specparam_declaration_instance11491();
    specparam_declaration11492 specparam_declaration_instance11492();
    specparam_declaration11493 specparam_declaration_instance11493();
    specparam_declaration11494 specparam_declaration_instance11494();
    specparam_declaration11495 specparam_declaration_instance11495();
    specparam_declaration11496 specparam_declaration_instance11496();
    specparam_declaration11497 specparam_declaration_instance11497();
    specparam_declaration11498 specparam_declaration_instance11498();
    specparam_declaration11499 specparam_declaration_instance11499();
    specparam_declaration11500 specparam_declaration_instance11500();
    specparam_declaration11501 specparam_declaration_instance11501();
    specparam_declaration11502 specparam_declaration_instance11502();
    specparam_declaration11503 specparam_declaration_instance11503();
    specparam_declaration11504 specparam_declaration_instance11504();
    specparam_declaration11505 specparam_declaration_instance11505();
    specparam_declaration11506 specparam_declaration_instance11506();
    specparam_declaration11507 specparam_declaration_instance11507();
    specparam_declaration11508 specparam_declaration_instance11508();
    specparam_declaration11509 specparam_declaration_instance11509();
    specparam_declaration11510 specparam_declaration_instance11510();
    specparam_declaration11511 specparam_declaration_instance11511();
    specparam_declaration11512 specparam_declaration_instance11512();
    specparam_declaration11513 specparam_declaration_instance11513();
    specparam_declaration11514 specparam_declaration_instance11514();
    specparam_declaration11515 specparam_declaration_instance11515();
    specparam_declaration11516 specparam_declaration_instance11516();
    specparam_declaration11517 specparam_declaration_instance11517();
    specparam_declaration11518 specparam_declaration_instance11518();
    specparam_declaration11519 specparam_declaration_instance11519();
    specparam_declaration11520 specparam_declaration_instance11520();
    specparam_declaration11521 specparam_declaration_instance11521();
    specparam_declaration11522 specparam_declaration_instance11522();
    specparam_declaration11523 specparam_declaration_instance11523();
    specparam_declaration11524 specparam_declaration_instance11524();
    specparam_declaration11525 specparam_declaration_instance11525();
    specparam_declaration11526 specparam_declaration_instance11526();
    specparam_declaration11527 specparam_declaration_instance11527();
    specparam_declaration11528 specparam_declaration_instance11528();
    specparam_declaration11529 specparam_declaration_instance11529();
    specparam_declaration11530 specparam_declaration_instance11530();
    specparam_declaration11531 specparam_declaration_instance11531();
    specparam_declaration11532 specparam_declaration_instance11532();
    specparam_declaration11533 specparam_declaration_instance11533();
    specparam_declaration11534 specparam_declaration_instance11534();
    specparam_declaration11535 specparam_declaration_instance11535();
    specparam_declaration11536 specparam_declaration_instance11536();
    specparam_declaration11537 specparam_declaration_instance11537();
    specparam_declaration11538 specparam_declaration_instance11538();
    specparam_declaration11539 specparam_declaration_instance11539();
    specparam_declaration11540 specparam_declaration_instance11540();
    specparam_declaration11541 specparam_declaration_instance11541();
    specparam_declaration11542 specparam_declaration_instance11542();
    specparam_declaration11543 specparam_declaration_instance11543();
    specparam_declaration11544 specparam_declaration_instance11544();
    specparam_declaration11545 specparam_declaration_instance11545();
    specparam_declaration11546 specparam_declaration_instance11546();
    specparam_declaration11547 specparam_declaration_instance11547();
    specparam_declaration11548 specparam_declaration_instance11548();
    specparam_declaration11549 specparam_declaration_instance11549();
    specparam_declaration11550 specparam_declaration_instance11550();
    specparam_declaration11551 specparam_declaration_instance11551();
    specparam_declaration11552 specparam_declaration_instance11552();
    specparam_declaration11553 specparam_declaration_instance11553();
    specparam_declaration11554 specparam_declaration_instance11554();
    specparam_declaration11555 specparam_declaration_instance11555();
    specparam_declaration11556 specparam_declaration_instance11556();
    specparam_declaration11557 specparam_declaration_instance11557();
    specparam_declaration11558 specparam_declaration_instance11558();
    specparam_declaration11559 specparam_declaration_instance11559();
    specparam_declaration11560 specparam_declaration_instance11560();
    specparam_declaration11561 specparam_declaration_instance11561();
    specparam_declaration11562 specparam_declaration_instance11562();
    specparam_declaration11563 specparam_declaration_instance11563();
    specparam_declaration11564 specparam_declaration_instance11564();
    specparam_declaration11565 specparam_declaration_instance11565();
    specparam_declaration11566 specparam_declaration_instance11566();
    specparam_declaration11567 specparam_declaration_instance11567();
    specparam_declaration11568 specparam_declaration_instance11568();
    specparam_declaration11569 specparam_declaration_instance11569();
    specparam_declaration11570 specparam_declaration_instance11570();
    specparam_declaration11571 specparam_declaration_instance11571();
    specparam_declaration11572 specparam_declaration_instance11572();
    specparam_declaration11573 specparam_declaration_instance11573();
    specparam_declaration11574 specparam_declaration_instance11574();
    specparam_declaration11575 specparam_declaration_instance11575();
    specparam_declaration11576 specparam_declaration_instance11576();
    specparam_declaration11577 specparam_declaration_instance11577();
    specparam_declaration11578 specparam_declaration_instance11578();
    specparam_declaration11579 specparam_declaration_instance11579();
    specparam_declaration11580 specparam_declaration_instance11580();
    specparam_declaration11581 specparam_declaration_instance11581();
    specparam_declaration11582 specparam_declaration_instance11582();
    specparam_declaration11583 specparam_declaration_instance11583();
    specparam_declaration11584 specparam_declaration_instance11584();
    specparam_declaration11585 specparam_declaration_instance11585();
    specparam_declaration11586 specparam_declaration_instance11586();
    specparam_declaration11587 specparam_declaration_instance11587();
    specparam_declaration11588 specparam_declaration_instance11588();
    specparam_declaration11589 specparam_declaration_instance11589();
    specparam_declaration11590 specparam_declaration_instance11590();
    specparam_declaration11591 specparam_declaration_instance11591();
    specparam_declaration11592 specparam_declaration_instance11592();
    specparam_declaration11593 specparam_declaration_instance11593();
    specparam_declaration11594 specparam_declaration_instance11594();
    specparam_declaration11595 specparam_declaration_instance11595();
    specparam_declaration11596 specparam_declaration_instance11596();
    specparam_declaration11597 specparam_declaration_instance11597();
    specparam_declaration11598 specparam_declaration_instance11598();
    specparam_declaration11599 specparam_declaration_instance11599();
    specparam_declaration11600 specparam_declaration_instance11600();
    specparam_declaration11601 specparam_declaration_instance11601();
    specparam_declaration11602 specparam_declaration_instance11602();
    specparam_declaration11603 specparam_declaration_instance11603();
    specparam_declaration11604 specparam_declaration_instance11604();
    specparam_declaration11605 specparam_declaration_instance11605();
    specparam_declaration11606 specparam_declaration_instance11606();
    specparam_declaration11607 specparam_declaration_instance11607();
    specparam_declaration11608 specparam_declaration_instance11608();
    specparam_declaration11609 specparam_declaration_instance11609();
    specparam_declaration11610 specparam_declaration_instance11610();
    specparam_declaration11611 specparam_declaration_instance11611();
    specparam_declaration11612 specparam_declaration_instance11612();
    specparam_declaration11613 specparam_declaration_instance11613();
    specparam_declaration11614 specparam_declaration_instance11614();
    specparam_declaration11615 specparam_declaration_instance11615();
    specparam_declaration11616 specparam_declaration_instance11616();
    specparam_declaration11617 specparam_declaration_instance11617();
    specparam_declaration11618 specparam_declaration_instance11618();
    specparam_declaration11619 specparam_declaration_instance11619();
    specparam_declaration11620 specparam_declaration_instance11620();
    specparam_declaration11621 specparam_declaration_instance11621();
    specparam_declaration11622 specparam_declaration_instance11622();
    specparam_declaration11623 specparam_declaration_instance11623();
    specparam_declaration11624 specparam_declaration_instance11624();
    specparam_declaration11625 specparam_declaration_instance11625();
    specparam_declaration11626 specparam_declaration_instance11626();
    specparam_declaration11627 specparam_declaration_instance11627();
    specparam_declaration11628 specparam_declaration_instance11628();
    specparam_declaration11629 specparam_declaration_instance11629();
    specparam_declaration11630 specparam_declaration_instance11630();
    specparam_declaration11631 specparam_declaration_instance11631();
    specparam_declaration11632 specparam_declaration_instance11632();
    specparam_declaration11633 specparam_declaration_instance11633();
    specparam_declaration11634 specparam_declaration_instance11634();
    specparam_declaration11635 specparam_declaration_instance11635();
    specparam_declaration11636 specparam_declaration_instance11636();
    specparam_declaration11637 specparam_declaration_instance11637();
    specparam_declaration11638 specparam_declaration_instance11638();
    specparam_declaration11639 specparam_declaration_instance11639();
    specparam_declaration11640 specparam_declaration_instance11640();
    specparam_declaration11641 specparam_declaration_instance11641();
    specparam_declaration11642 specparam_declaration_instance11642();
    specparam_declaration11643 specparam_declaration_instance11643();
    specparam_declaration11644 specparam_declaration_instance11644();
    specparam_declaration11645 specparam_declaration_instance11645();
    specparam_declaration11646 specparam_declaration_instance11646();
    specparam_declaration11647 specparam_declaration_instance11647();
    specparam_declaration11648 specparam_declaration_instance11648();
    specparam_declaration11649 specparam_declaration_instance11649();
    specparam_declaration11650 specparam_declaration_instance11650();
    specparam_declaration11651 specparam_declaration_instance11651();
    specparam_declaration11652 specparam_declaration_instance11652();
    specparam_declaration11653 specparam_declaration_instance11653();
    specparam_declaration11654 specparam_declaration_instance11654();
    specparam_declaration11655 specparam_declaration_instance11655();
    specparam_declaration11656 specparam_declaration_instance11656();
    specparam_declaration11657 specparam_declaration_instance11657();
    specparam_declaration11658 specparam_declaration_instance11658();
    specparam_declaration11659 specparam_declaration_instance11659();
    specparam_declaration11660 specparam_declaration_instance11660();
    specparam_declaration11661 specparam_declaration_instance11661();
    specparam_declaration11662 specparam_declaration_instance11662();
    specparam_declaration11663 specparam_declaration_instance11663();
    specparam_declaration11664 specparam_declaration_instance11664();
    specparam_declaration11665 specparam_declaration_instance11665();
    specparam_declaration11666 specparam_declaration_instance11666();
    specparam_declaration11667 specparam_declaration_instance11667();
    specparam_declaration11668 specparam_declaration_instance11668();
    specparam_declaration11669 specparam_declaration_instance11669();
    specparam_declaration11670 specparam_declaration_instance11670();
    specparam_declaration11671 specparam_declaration_instance11671();
    specparam_declaration11672 specparam_declaration_instance11672();
    specparam_declaration11673 specparam_declaration_instance11673();
    specparam_declaration11674 specparam_declaration_instance11674();
    specparam_declaration11675 specparam_declaration_instance11675();
    specparam_declaration11676 specparam_declaration_instance11676();
    specparam_declaration11677 specparam_declaration_instance11677();
    specparam_declaration11678 specparam_declaration_instance11678();
    specparam_declaration11679 specparam_declaration_instance11679();
    specparam_declaration11680 specparam_declaration_instance11680();
    specparam_declaration11681 specparam_declaration_instance11681();
    specparam_declaration11682 specparam_declaration_instance11682();
    specparam_declaration11683 specparam_declaration_instance11683();
    specparam_declaration11684 specparam_declaration_instance11684();
    specparam_declaration11685 specparam_declaration_instance11685();
    specparam_declaration11686 specparam_declaration_instance11686();
    specparam_declaration11687 specparam_declaration_instance11687();
    specparam_declaration11688 specparam_declaration_instance11688();
    specparam_declaration11689 specparam_declaration_instance11689();
    specparam_declaration11690 specparam_declaration_instance11690();
    specparam_declaration11691 specparam_declaration_instance11691();
    specparam_declaration11692 specparam_declaration_instance11692();
    specparam_declaration11693 specparam_declaration_instance11693();
    specparam_declaration11694 specparam_declaration_instance11694();
    specparam_declaration11695 specparam_declaration_instance11695();
    specparam_declaration11696 specparam_declaration_instance11696();
    specparam_declaration11697 specparam_declaration_instance11697();
    specparam_declaration11698 specparam_declaration_instance11698();
    specparam_declaration11699 specparam_declaration_instance11699();
    specparam_declaration11700 specparam_declaration_instance11700();
    specparam_declaration11701 specparam_declaration_instance11701();
    specparam_declaration11702 specparam_declaration_instance11702();
    specparam_declaration11703 specparam_declaration_instance11703();
    specparam_declaration11704 specparam_declaration_instance11704();
    specparam_declaration11705 specparam_declaration_instance11705();
    specparam_declaration11706 specparam_declaration_instance11706();
    specparam_declaration11707 specparam_declaration_instance11707();
    specparam_declaration11708 specparam_declaration_instance11708();
    specparam_declaration11709 specparam_declaration_instance11709();
    specparam_declaration11710 specparam_declaration_instance11710();
    specparam_declaration11711 specparam_declaration_instance11711();
    specparam_declaration11712 specparam_declaration_instance11712();
    specparam_declaration11713 specparam_declaration_instance11713();
    specparam_declaration11714 specparam_declaration_instance11714();
    specparam_declaration11715 specparam_declaration_instance11715();
    specparam_declaration11716 specparam_declaration_instance11716();
    specparam_declaration11717 specparam_declaration_instance11717();
    specparam_declaration11718 specparam_declaration_instance11718();
    specparam_declaration11719 specparam_declaration_instance11719();
    specparam_declaration11720 specparam_declaration_instance11720();
    specparam_declaration11721 specparam_declaration_instance11721();
    specparam_declaration11722 specparam_declaration_instance11722();
    specparam_declaration11723 specparam_declaration_instance11723();
    specparam_declaration11724 specparam_declaration_instance11724();
    specparam_declaration11725 specparam_declaration_instance11725();
    specparam_declaration11726 specparam_declaration_instance11726();
    specparam_declaration11727 specparam_declaration_instance11727();
    specparam_declaration11728 specparam_declaration_instance11728();
    specparam_declaration11729 specparam_declaration_instance11729();
    specparam_declaration11730 specparam_declaration_instance11730();
    specparam_declaration11731 specparam_declaration_instance11731();
    specparam_declaration11732 specparam_declaration_instance11732();
    specparam_declaration11733 specparam_declaration_instance11733();
    specparam_declaration11734 specparam_declaration_instance11734();
    specparam_declaration11735 specparam_declaration_instance11735();
    specparam_declaration11736 specparam_declaration_instance11736();
    specparam_declaration11737 specparam_declaration_instance11737();
    specparam_declaration11738 specparam_declaration_instance11738();
    specparam_declaration11739 specparam_declaration_instance11739();
    specparam_declaration11740 specparam_declaration_instance11740();
    specparam_declaration11741 specparam_declaration_instance11741();
    specparam_declaration11742 specparam_declaration_instance11742();
    specparam_declaration11743 specparam_declaration_instance11743();
    specparam_declaration11744 specparam_declaration_instance11744();
    specparam_declaration11745 specparam_declaration_instance11745();
    specparam_declaration11746 specparam_declaration_instance11746();
    specparam_declaration11747 specparam_declaration_instance11747();
    specparam_declaration11748 specparam_declaration_instance11748();
    specparam_declaration11749 specparam_declaration_instance11749();
    specparam_declaration11750 specparam_declaration_instance11750();
    specparam_declaration11751 specparam_declaration_instance11751();
    specparam_declaration11752 specparam_declaration_instance11752();
    specparam_declaration11753 specparam_declaration_instance11753();
    specparam_declaration11754 specparam_declaration_instance11754();
    specparam_declaration11755 specparam_declaration_instance11755();
    specparam_declaration11756 specparam_declaration_instance11756();
    specparam_declaration11757 specparam_declaration_instance11757();
    specparam_declaration11758 specparam_declaration_instance11758();
    specparam_declaration11759 specparam_declaration_instance11759();
    specparam_declaration11760 specparam_declaration_instance11760();
    specparam_declaration11761 specparam_declaration_instance11761();
    specparam_declaration11762 specparam_declaration_instance11762();
    specparam_declaration11763 specparam_declaration_instance11763();
    specparam_declaration11764 specparam_declaration_instance11764();
    specparam_declaration11765 specparam_declaration_instance11765();
    specparam_declaration11766 specparam_declaration_instance11766();
    specparam_declaration11767 specparam_declaration_instance11767();
    specparam_declaration11768 specparam_declaration_instance11768();
    specparam_declaration11769 specparam_declaration_instance11769();
    specparam_declaration11770 specparam_declaration_instance11770();
    specparam_declaration11771 specparam_declaration_instance11771();
    specparam_declaration11772 specparam_declaration_instance11772();
    specparam_declaration11773 specparam_declaration_instance11773();
    specparam_declaration11774 specparam_declaration_instance11774();
    specparam_declaration11775 specparam_declaration_instance11775();
    specparam_declaration11776 specparam_declaration_instance11776();
    specparam_declaration11777 specparam_declaration_instance11777();
    specparam_declaration11778 specparam_declaration_instance11778();
    specparam_declaration11779 specparam_declaration_instance11779();
    specparam_declaration11780 specparam_declaration_instance11780();
    specparam_declaration11781 specparam_declaration_instance11781();
    specparam_declaration11782 specparam_declaration_instance11782();
    specparam_declaration11783 specparam_declaration_instance11783();
    specparam_declaration11784 specparam_declaration_instance11784();
    specparam_declaration11785 specparam_declaration_instance11785();
    specparam_declaration11786 specparam_declaration_instance11786();
    specparam_declaration11787 specparam_declaration_instance11787();
    specparam_declaration11788 specparam_declaration_instance11788();
    specparam_declaration11789 specparam_declaration_instance11789();
    specparam_declaration11790 specparam_declaration_instance11790();
    specparam_declaration11791 specparam_declaration_instance11791();
    specparam_declaration11792 specparam_declaration_instance11792();
    specparam_declaration11793 specparam_declaration_instance11793();
    specparam_declaration11794 specparam_declaration_instance11794();
    specparam_declaration11795 specparam_declaration_instance11795();
    specparam_declaration11796 specparam_declaration_instance11796();
    specparam_declaration11797 specparam_declaration_instance11797();
    specparam_declaration11798 specparam_declaration_instance11798();
    specparam_declaration11799 specparam_declaration_instance11799();
    specparam_declaration11800 specparam_declaration_instance11800();
    specparam_declaration11801 specparam_declaration_instance11801();
    specparam_declaration11802 specparam_declaration_instance11802();
    specparam_declaration11803 specparam_declaration_instance11803();
    specparam_declaration11804 specparam_declaration_instance11804();
    specparam_declaration11805 specparam_declaration_instance11805();
    specparam_declaration11806 specparam_declaration_instance11806();
    specparam_declaration11807 specparam_declaration_instance11807();
    specparam_declaration11808 specparam_declaration_instance11808();
    specparam_declaration11809 specparam_declaration_instance11809();
    specparam_declaration11810 specparam_declaration_instance11810();
    specparam_declaration11811 specparam_declaration_instance11811();
    specparam_declaration11812 specparam_declaration_instance11812();
    specparam_declaration11813 specparam_declaration_instance11813();
    specparam_declaration11814 specparam_declaration_instance11814();
    specparam_declaration11815 specparam_declaration_instance11815();
    specparam_declaration11816 specparam_declaration_instance11816();
    specparam_declaration11817 specparam_declaration_instance11817();
    specparam_declaration11818 specparam_declaration_instance11818();
    specparam_declaration11819 specparam_declaration_instance11819();
    specparam_declaration11820 specparam_declaration_instance11820();
    specparam_declaration11821 specparam_declaration_instance11821();
    specparam_declaration11822 specparam_declaration_instance11822();
    specparam_declaration11823 specparam_declaration_instance11823();
    specparam_declaration11824 specparam_declaration_instance11824();
    specparam_declaration11825 specparam_declaration_instance11825();
    specparam_declaration11826 specparam_declaration_instance11826();
    specparam_declaration11827 specparam_declaration_instance11827();
    specparam_declaration11828 specparam_declaration_instance11828();
    specparam_declaration11829 specparam_declaration_instance11829();
    specparam_declaration11830 specparam_declaration_instance11830();
    specparam_declaration11831 specparam_declaration_instance11831();
    specparam_declaration11832 specparam_declaration_instance11832();
    specparam_declaration11833 specparam_declaration_instance11833();
    specparam_declaration11834 specparam_declaration_instance11834();
    specparam_declaration11835 specparam_declaration_instance11835();
    specparam_declaration11836 specparam_declaration_instance11836();
    specparam_declaration11837 specparam_declaration_instance11837();
    specparam_declaration11838 specparam_declaration_instance11838();
    specparam_declaration11839 specparam_declaration_instance11839();
    specparam_declaration11840 specparam_declaration_instance11840();
    specparam_declaration11841 specparam_declaration_instance11841();
    specparam_declaration11842 specparam_declaration_instance11842();
    specparam_declaration11843 specparam_declaration_instance11843();
    specparam_declaration11844 specparam_declaration_instance11844();
    specparam_declaration11845 specparam_declaration_instance11845();
    specparam_declaration11846 specparam_declaration_instance11846();
    specparam_declaration11847 specparam_declaration_instance11847();
    specparam_declaration11848 specparam_declaration_instance11848();
    specparam_declaration11849 specparam_declaration_instance11849();
    specparam_declaration11850 specparam_declaration_instance11850();
    specparam_declaration11851 specparam_declaration_instance11851();
    specparam_declaration11852 specparam_declaration_instance11852();
    specparam_declaration11853 specparam_declaration_instance11853();
    specparam_declaration11854 specparam_declaration_instance11854();
    specparam_declaration11855 specparam_declaration_instance11855();
    specparam_declaration11856 specparam_declaration_instance11856();
    specparam_declaration11857 specparam_declaration_instance11857();
    specparam_declaration11858 specparam_declaration_instance11858();
    specparam_declaration11859 specparam_declaration_instance11859();
    specparam_declaration11860 specparam_declaration_instance11860();
    specparam_declaration11861 specparam_declaration_instance11861();
    specparam_declaration11862 specparam_declaration_instance11862();
    specparam_declaration11863 specparam_declaration_instance11863();
    specparam_declaration11864 specparam_declaration_instance11864();
    specparam_declaration11865 specparam_declaration_instance11865();
    specparam_declaration11866 specparam_declaration_instance11866();
    specparam_declaration11867 specparam_declaration_instance11867();
    specparam_declaration11868 specparam_declaration_instance11868();
    specparam_declaration11869 specparam_declaration_instance11869();
    specparam_declaration11870 specparam_declaration_instance11870();
    specparam_declaration11871 specparam_declaration_instance11871();
    specparam_declaration11872 specparam_declaration_instance11872();
    specparam_declaration11873 specparam_declaration_instance11873();
    specparam_declaration11874 specparam_declaration_instance11874();
    specparam_declaration11875 specparam_declaration_instance11875();
    specparam_declaration11876 specparam_declaration_instance11876();
    specparam_declaration11877 specparam_declaration_instance11877();
    specparam_declaration11878 specparam_declaration_instance11878();
    specparam_declaration11879 specparam_declaration_instance11879();
    specparam_declaration11880 specparam_declaration_instance11880();
    specparam_declaration11881 specparam_declaration_instance11881();
    specparam_declaration11882 specparam_declaration_instance11882();
    specparam_declaration11883 specparam_declaration_instance11883();
    specparam_declaration11884 specparam_declaration_instance11884();
    specparam_declaration11885 specparam_declaration_instance11885();
    specparam_declaration11886 specparam_declaration_instance11886();
    specparam_declaration11887 specparam_declaration_instance11887();
    specparam_declaration11888 specparam_declaration_instance11888();
    specparam_declaration11889 specparam_declaration_instance11889();
    specparam_declaration11890 specparam_declaration_instance11890();
    specparam_declaration11891 specparam_declaration_instance11891();
    specparam_declaration11892 specparam_declaration_instance11892();
    specparam_declaration11893 specparam_declaration_instance11893();
    specparam_declaration11894 specparam_declaration_instance11894();
    specparam_declaration11895 specparam_declaration_instance11895();
    specparam_declaration11896 specparam_declaration_instance11896();
    specparam_declaration11897 specparam_declaration_instance11897();
    specparam_declaration11898 specparam_declaration_instance11898();
    specparam_declaration11899 specparam_declaration_instance11899();
    specparam_declaration11900 specparam_declaration_instance11900();
    specparam_declaration11901 specparam_declaration_instance11901();
    specparam_declaration11902 specparam_declaration_instance11902();
    specparam_declaration11903 specparam_declaration_instance11903();
    specparam_declaration11904 specparam_declaration_instance11904();
    specparam_declaration11905 specparam_declaration_instance11905();
    specparam_declaration11906 specparam_declaration_instance11906();
    specparam_declaration11907 specparam_declaration_instance11907();
    specparam_declaration11908 specparam_declaration_instance11908();
    specparam_declaration11909 specparam_declaration_instance11909();
    specparam_declaration11910 specparam_declaration_instance11910();
    specparam_declaration11911 specparam_declaration_instance11911();
    specparam_declaration11912 specparam_declaration_instance11912();
    specparam_declaration11913 specparam_declaration_instance11913();
    specparam_declaration11914 specparam_declaration_instance11914();
    specparam_declaration11915 specparam_declaration_instance11915();
    specparam_declaration11916 specparam_declaration_instance11916();
    specparam_declaration11917 specparam_declaration_instance11917();
    specparam_declaration11918 specparam_declaration_instance11918();
    specparam_declaration11919 specparam_declaration_instance11919();
    specparam_declaration11920 specparam_declaration_instance11920();
    specparam_declaration11921 specparam_declaration_instance11921();
    specparam_declaration11922 specparam_declaration_instance11922();
    specparam_declaration11923 specparam_declaration_instance11923();
    specparam_declaration11924 specparam_declaration_instance11924();
    specparam_declaration11925 specparam_declaration_instance11925();
    specparam_declaration11926 specparam_declaration_instance11926();
    specparam_declaration11927 specparam_declaration_instance11927();
    specparam_declaration11928 specparam_declaration_instance11928();
    specparam_declaration11929 specparam_declaration_instance11929();
    specparam_declaration11930 specparam_declaration_instance11930();
    specparam_declaration11931 specparam_declaration_instance11931();
    specparam_declaration11932 specparam_declaration_instance11932();
    specparam_declaration11933 specparam_declaration_instance11933();
    specparam_declaration11934 specparam_declaration_instance11934();
    specparam_declaration11935 specparam_declaration_instance11935();
    specparam_declaration11936 specparam_declaration_instance11936();
    specparam_declaration11937 specparam_declaration_instance11937();
    specparam_declaration11938 specparam_declaration_instance11938();
    specparam_declaration11939 specparam_declaration_instance11939();
    specparam_declaration11940 specparam_declaration_instance11940();
    specparam_declaration11941 specparam_declaration_instance11941();
    specparam_declaration11942 specparam_declaration_instance11942();
    specparam_declaration11943 specparam_declaration_instance11943();
    specparam_declaration11944 specparam_declaration_instance11944();
    specparam_declaration11945 specparam_declaration_instance11945();
    specparam_declaration11946 specparam_declaration_instance11946();
    specparam_declaration11947 specparam_declaration_instance11947();
    specparam_declaration11948 specparam_declaration_instance11948();
    specparam_declaration11949 specparam_declaration_instance11949();
    specparam_declaration11950 specparam_declaration_instance11950();
    specparam_declaration11951 specparam_declaration_instance11951();
    specparam_declaration11952 specparam_declaration_instance11952();
    specparam_declaration11953 specparam_declaration_instance11953();
    specparam_declaration11954 specparam_declaration_instance11954();
    specparam_declaration11955 specparam_declaration_instance11955();
    specparam_declaration11956 specparam_declaration_instance11956();
    specparam_declaration11957 specparam_declaration_instance11957();
    specparam_declaration11958 specparam_declaration_instance11958();
    specparam_declaration11959 specparam_declaration_instance11959();
    specparam_declaration11960 specparam_declaration_instance11960();
    specparam_declaration11961 specparam_declaration_instance11961();
    specparam_declaration11962 specparam_declaration_instance11962();
    specparam_declaration11963 specparam_declaration_instance11963();
    specparam_declaration11964 specparam_declaration_instance11964();
    specparam_declaration11965 specparam_declaration_instance11965();
    specparam_declaration11966 specparam_declaration_instance11966();
    specparam_declaration11967 specparam_declaration_instance11967();
    specparam_declaration11968 specparam_declaration_instance11968();
    specparam_declaration11969 specparam_declaration_instance11969();
    specparam_declaration11970 specparam_declaration_instance11970();
    specparam_declaration11971 specparam_declaration_instance11971();
    specparam_declaration11972 specparam_declaration_instance11972();
    specparam_declaration11973 specparam_declaration_instance11973();
    specparam_declaration11974 specparam_declaration_instance11974();
    specparam_declaration11975 specparam_declaration_instance11975();
    specparam_declaration11976 specparam_declaration_instance11976();
    specparam_declaration11977 specparam_declaration_instance11977();
    specparam_declaration11978 specparam_declaration_instance11978();
    specparam_declaration11979 specparam_declaration_instance11979();
    specparam_declaration11980 specparam_declaration_instance11980();
    specparam_declaration11981 specparam_declaration_instance11981();
    specparam_declaration11982 specparam_declaration_instance11982();
    specparam_declaration11983 specparam_declaration_instance11983();
    specparam_declaration11984 specparam_declaration_instance11984();
    specparam_declaration11985 specparam_declaration_instance11985();
    specparam_declaration11986 specparam_declaration_instance11986();
    specparam_declaration11987 specparam_declaration_instance11987();
    specparam_declaration11988 specparam_declaration_instance11988();
    specparam_declaration11989 specparam_declaration_instance11989();
    specparam_declaration11990 specparam_declaration_instance11990();
    specparam_declaration11991 specparam_declaration_instance11991();
    specparam_declaration11992 specparam_declaration_instance11992();
    specparam_declaration11993 specparam_declaration_instance11993();
    specparam_declaration11994 specparam_declaration_instance11994();
    specparam_declaration11995 specparam_declaration_instance11995();
    specparam_declaration11996 specparam_declaration_instance11996();
    specparam_declaration11997 specparam_declaration_instance11997();
    specparam_declaration11998 specparam_declaration_instance11998();
    specparam_declaration11999 specparam_declaration_instance11999();
    specparam_declaration12000 specparam_declaration_instance12000();
    specparam_declaration12001 specparam_declaration_instance12001();
    specparam_declaration12002 specparam_declaration_instance12002();
    specparam_declaration12003 specparam_declaration_instance12003();
    specparam_declaration12004 specparam_declaration_instance12004();
    specparam_declaration12005 specparam_declaration_instance12005();
    specparam_declaration12006 specparam_declaration_instance12006();
    specparam_declaration12007 specparam_declaration_instance12007();
    specparam_declaration12008 specparam_declaration_instance12008();
    specparam_declaration12009 specparam_declaration_instance12009();
    specparam_declaration12010 specparam_declaration_instance12010();
    specparam_declaration12011 specparam_declaration_instance12011();
    specparam_declaration12012 specparam_declaration_instance12012();
    specparam_declaration12013 specparam_declaration_instance12013();
    specparam_declaration12014 specparam_declaration_instance12014();
    specparam_declaration12015 specparam_declaration_instance12015();
    specparam_declaration12016 specparam_declaration_instance12016();
    specparam_declaration12017 specparam_declaration_instance12017();
    specparam_declaration12018 specparam_declaration_instance12018();
    specparam_declaration12019 specparam_declaration_instance12019();
    specparam_declaration12020 specparam_declaration_instance12020();
    specparam_declaration12021 specparam_declaration_instance12021();
    specparam_declaration12022 specparam_declaration_instance12022();
    specparam_declaration12023 specparam_declaration_instance12023();
    specparam_declaration12024 specparam_declaration_instance12024();
    specparam_declaration12025 specparam_declaration_instance12025();
    specparam_declaration12026 specparam_declaration_instance12026();
    specparam_declaration12027 specparam_declaration_instance12027();
    specparam_declaration12028 specparam_declaration_instance12028();
    specparam_declaration12029 specparam_declaration_instance12029();
    specparam_declaration12030 specparam_declaration_instance12030();
    specparam_declaration12031 specparam_declaration_instance12031();
    specparam_declaration12032 specparam_declaration_instance12032();
    specparam_declaration12033 specparam_declaration_instance12033();
    specparam_declaration12034 specparam_declaration_instance12034();
    specparam_declaration12035 specparam_declaration_instance12035();
    specparam_declaration12036 specparam_declaration_instance12036();
    specparam_declaration12037 specparam_declaration_instance12037();
    specparam_declaration12038 specparam_declaration_instance12038();
    specparam_declaration12039 specparam_declaration_instance12039();
    specparam_declaration12040 specparam_declaration_instance12040();
    specparam_declaration12041 specparam_declaration_instance12041();
    specparam_declaration12042 specparam_declaration_instance12042();
    specparam_declaration12043 specparam_declaration_instance12043();
    specparam_declaration12044 specparam_declaration_instance12044();
    specparam_declaration12045 specparam_declaration_instance12045();
    specparam_declaration12046 specparam_declaration_instance12046();
    specparam_declaration12047 specparam_declaration_instance12047();
    specparam_declaration12048 specparam_declaration_instance12048();
    specparam_declaration12049 specparam_declaration_instance12049();
    specparam_declaration12050 specparam_declaration_instance12050();
    specparam_declaration12051 specparam_declaration_instance12051();
    specparam_declaration12052 specparam_declaration_instance12052();
    specparam_declaration12053 specparam_declaration_instance12053();
    specparam_declaration12054 specparam_declaration_instance12054();
    specparam_declaration12055 specparam_declaration_instance12055();
    specparam_declaration12056 specparam_declaration_instance12056();
    specparam_declaration12057 specparam_declaration_instance12057();
    specparam_declaration12058 specparam_declaration_instance12058();
    specparam_declaration12059 specparam_declaration_instance12059();
    specparam_declaration12060 specparam_declaration_instance12060();
    specparam_declaration12061 specparam_declaration_instance12061();
    specparam_declaration12062 specparam_declaration_instance12062();
    specparam_declaration12063 specparam_declaration_instance12063();
    specparam_declaration12064 specparam_declaration_instance12064();
    specparam_declaration12065 specparam_declaration_instance12065();
    specparam_declaration12066 specparam_declaration_instance12066();
    specparam_declaration12067 specparam_declaration_instance12067();
    specparam_declaration12068 specparam_declaration_instance12068();
    specparam_declaration12069 specparam_declaration_instance12069();
    specparam_declaration12070 specparam_declaration_instance12070();
    specparam_declaration12071 specparam_declaration_instance12071();
    specparam_declaration12072 specparam_declaration_instance12072();
    specparam_declaration12073 specparam_declaration_instance12073();
    specparam_declaration12074 specparam_declaration_instance12074();
    specparam_declaration12075 specparam_declaration_instance12075();
    specparam_declaration12076 specparam_declaration_instance12076();
    specparam_declaration12077 specparam_declaration_instance12077();
    specparam_declaration12078 specparam_declaration_instance12078();
    specparam_declaration12079 specparam_declaration_instance12079();
    specparam_declaration12080 specparam_declaration_instance12080();
    specparam_declaration12081 specparam_declaration_instance12081();
    specparam_declaration12082 specparam_declaration_instance12082();
    specparam_declaration12083 specparam_declaration_instance12083();
    specparam_declaration12084 specparam_declaration_instance12084();
    specparam_declaration12085 specparam_declaration_instance12085();
    specparam_declaration12086 specparam_declaration_instance12086();
    specparam_declaration12087 specparam_declaration_instance12087();
    specparam_declaration12088 specparam_declaration_instance12088();
    specparam_declaration12089 specparam_declaration_instance12089();
    specparam_declaration12090 specparam_declaration_instance12090();
    specparam_declaration12091 specparam_declaration_instance12091();
    specparam_declaration12092 specparam_declaration_instance12092();
    specparam_declaration12093 specparam_declaration_instance12093();
    specparam_declaration12094 specparam_declaration_instance12094();
    specparam_declaration12095 specparam_declaration_instance12095();
    specparam_declaration12096 specparam_declaration_instance12096();
    specparam_declaration12097 specparam_declaration_instance12097();
    specparam_declaration12098 specparam_declaration_instance12098();
    specparam_declaration12099 specparam_declaration_instance12099();
    specparam_declaration12100 specparam_declaration_instance12100();
    specparam_declaration12101 specparam_declaration_instance12101();
    specparam_declaration12102 specparam_declaration_instance12102();
    specparam_declaration12103 specparam_declaration_instance12103();
    specparam_declaration12104 specparam_declaration_instance12104();
    specparam_declaration12105 specparam_declaration_instance12105();
    specparam_declaration12106 specparam_declaration_instance12106();
    specparam_declaration12107 specparam_declaration_instance12107();
    specparam_declaration12108 specparam_declaration_instance12108();
    specparam_declaration12109 specparam_declaration_instance12109();
    specparam_declaration12110 specparam_declaration_instance12110();
    specparam_declaration12111 specparam_declaration_instance12111();
    specparam_declaration12112 specparam_declaration_instance12112();
    specparam_declaration12113 specparam_declaration_instance12113();
    specparam_declaration12114 specparam_declaration_instance12114();
    specparam_declaration12115 specparam_declaration_instance12115();
    specparam_declaration12116 specparam_declaration_instance12116();
    specparam_declaration12117 specparam_declaration_instance12117();
    specparam_declaration12118 specparam_declaration_instance12118();
    specparam_declaration12119 specparam_declaration_instance12119();
    specparam_declaration12120 specparam_declaration_instance12120();
    specparam_declaration12121 specparam_declaration_instance12121();
    specparam_declaration12122 specparam_declaration_instance12122();
    specparam_declaration12123 specparam_declaration_instance12123();
    specparam_declaration12124 specparam_declaration_instance12124();
    specparam_declaration12125 specparam_declaration_instance12125();
    specparam_declaration12126 specparam_declaration_instance12126();
    specparam_declaration12127 specparam_declaration_instance12127();
    specparam_declaration12128 specparam_declaration_instance12128();
    specparam_declaration12129 specparam_declaration_instance12129();
    specparam_declaration12130 specparam_declaration_instance12130();
    specparam_declaration12131 specparam_declaration_instance12131();
    specparam_declaration12132 specparam_declaration_instance12132();
    specparam_declaration12133 specparam_declaration_instance12133();
    specparam_declaration12134 specparam_declaration_instance12134();
    specparam_declaration12135 specparam_declaration_instance12135();
    specparam_declaration12136 specparam_declaration_instance12136();
    specparam_declaration12137 specparam_declaration_instance12137();
    specparam_declaration12138 specparam_declaration_instance12138();
    specparam_declaration12139 specparam_declaration_instance12139();
    specparam_declaration12140 specparam_declaration_instance12140();
    specparam_declaration12141 specparam_declaration_instance12141();
    specparam_declaration12142 specparam_declaration_instance12142();
    specparam_declaration12143 specparam_declaration_instance12143();
    specparam_declaration12144 specparam_declaration_instance12144();
    specparam_declaration12145 specparam_declaration_instance12145();
    specparam_declaration12146 specparam_declaration_instance12146();
    specparam_declaration12147 specparam_declaration_instance12147();
    specparam_declaration12148 specparam_declaration_instance12148();
    specparam_declaration12149 specparam_declaration_instance12149();
    specparam_declaration12150 specparam_declaration_instance12150();
    specparam_declaration12151 specparam_declaration_instance12151();
    specparam_declaration12152 specparam_declaration_instance12152();
    specparam_declaration12153 specparam_declaration_instance12153();
    specparam_declaration12154 specparam_declaration_instance12154();
    specparam_declaration12155 specparam_declaration_instance12155();
    specparam_declaration12156 specparam_declaration_instance12156();
    specparam_declaration12157 specparam_declaration_instance12157();
    specparam_declaration12158 specparam_declaration_instance12158();
    specparam_declaration12159 specparam_declaration_instance12159();
    specparam_declaration12160 specparam_declaration_instance12160();
    specparam_declaration12161 specparam_declaration_instance12161();
    specparam_declaration12162 specparam_declaration_instance12162();
    specparam_declaration12163 specparam_declaration_instance12163();
    specparam_declaration12164 specparam_declaration_instance12164();
    specparam_declaration12165 specparam_declaration_instance12165();
    specparam_declaration12166 specparam_declaration_instance12166();
    specparam_declaration12167 specparam_declaration_instance12167();
    specparam_declaration12168 specparam_declaration_instance12168();
    specparam_declaration12169 specparam_declaration_instance12169();
    specparam_declaration12170 specparam_declaration_instance12170();
    specparam_declaration12171 specparam_declaration_instance12171();
    specparam_declaration12172 specparam_declaration_instance12172();
    specparam_declaration12173 specparam_declaration_instance12173();
    specparam_declaration12174 specparam_declaration_instance12174();
    specparam_declaration12175 specparam_declaration_instance12175();
    specparam_declaration12176 specparam_declaration_instance12176();
    specparam_declaration12177 specparam_declaration_instance12177();
    specparam_declaration12178 specparam_declaration_instance12178();
    specparam_declaration12179 specparam_declaration_instance12179();
    specparam_declaration12180 specparam_declaration_instance12180();
    specparam_declaration12181 specparam_declaration_instance12181();
    specparam_declaration12182 specparam_declaration_instance12182();
    specparam_declaration12183 specparam_declaration_instance12183();
    specparam_declaration12184 specparam_declaration_instance12184();
    specparam_declaration12185 specparam_declaration_instance12185();
    specparam_declaration12186 specparam_declaration_instance12186();
    specparam_declaration12187 specparam_declaration_instance12187();
    specparam_declaration12188 specparam_declaration_instance12188();
    specparam_declaration12189 specparam_declaration_instance12189();
    specparam_declaration12190 specparam_declaration_instance12190();
    specparam_declaration12191 specparam_declaration_instance12191();
    specparam_declaration12192 specparam_declaration_instance12192();
    specparam_declaration12193 specparam_declaration_instance12193();
    specparam_declaration12194 specparam_declaration_instance12194();
    specparam_declaration12195 specparam_declaration_instance12195();
    specparam_declaration12196 specparam_declaration_instance12196();
    specparam_declaration12197 specparam_declaration_instance12197();
    specparam_declaration12198 specparam_declaration_instance12198();
    specparam_declaration12199 specparam_declaration_instance12199();
    specparam_declaration12200 specparam_declaration_instance12200();
    specparam_declaration12201 specparam_declaration_instance12201();
    specparam_declaration12202 specparam_declaration_instance12202();
    specparam_declaration12203 specparam_declaration_instance12203();
    specparam_declaration12204 specparam_declaration_instance12204();
    specparam_declaration12205 specparam_declaration_instance12205();
    specparam_declaration12206 specparam_declaration_instance12206();
    specparam_declaration12207 specparam_declaration_instance12207();
    specparam_declaration12208 specparam_declaration_instance12208();
    specparam_declaration12209 specparam_declaration_instance12209();
    specparam_declaration12210 specparam_declaration_instance12210();
    specparam_declaration12211 specparam_declaration_instance12211();
    specparam_declaration12212 specparam_declaration_instance12212();
    specparam_declaration12213 specparam_declaration_instance12213();
    specparam_declaration12214 specparam_declaration_instance12214();
    specparam_declaration12215 specparam_declaration_instance12215();
    specparam_declaration12216 specparam_declaration_instance12216();
    specparam_declaration12217 specparam_declaration_instance12217();
    specparam_declaration12218 specparam_declaration_instance12218();
    specparam_declaration12219 specparam_declaration_instance12219();
    specparam_declaration12220 specparam_declaration_instance12220();
    specparam_declaration12221 specparam_declaration_instance12221();
    specparam_declaration12222 specparam_declaration_instance12222();
    specparam_declaration12223 specparam_declaration_instance12223();
    specparam_declaration12224 specparam_declaration_instance12224();
    specparam_declaration12225 specparam_declaration_instance12225();
    specparam_declaration12226 specparam_declaration_instance12226();
    specparam_declaration12227 specparam_declaration_instance12227();
    specparam_declaration12228 specparam_declaration_instance12228();
    specparam_declaration12229 specparam_declaration_instance12229();
    specparam_declaration12230 specparam_declaration_instance12230();
    specparam_declaration12231 specparam_declaration_instance12231();
    specparam_declaration12232 specparam_declaration_instance12232();
    specparam_declaration12233 specparam_declaration_instance12233();
    specparam_declaration12234 specparam_declaration_instance12234();
    specparam_declaration12235 specparam_declaration_instance12235();
    specparam_declaration12236 specparam_declaration_instance12236();
    specparam_declaration12237 specparam_declaration_instance12237();
    specparam_declaration12238 specparam_declaration_instance12238();
    specparam_declaration12239 specparam_declaration_instance12239();
    specparam_declaration12240 specparam_declaration_instance12240();
    specparam_declaration12241 specparam_declaration_instance12241();
    specparam_declaration12242 specparam_declaration_instance12242();
    specparam_declaration12243 specparam_declaration_instance12243();
    specparam_declaration12244 specparam_declaration_instance12244();
    specparam_declaration12245 specparam_declaration_instance12245();
    specparam_declaration12246 specparam_declaration_instance12246();
    specparam_declaration12247 specparam_declaration_instance12247();
    specparam_declaration12248 specparam_declaration_instance12248();
    specparam_declaration12249 specparam_declaration_instance12249();
    specparam_declaration12250 specparam_declaration_instance12250();
    specparam_declaration12251 specparam_declaration_instance12251();
    specparam_declaration12252 specparam_declaration_instance12252();
    specparam_declaration12253 specparam_declaration_instance12253();
    specparam_declaration12254 specparam_declaration_instance12254();
    specparam_declaration12255 specparam_declaration_instance12255();
    specparam_declaration12256 specparam_declaration_instance12256();
    specparam_declaration12257 specparam_declaration_instance12257();
    specparam_declaration12258 specparam_declaration_instance12258();
    specparam_declaration12259 specparam_declaration_instance12259();
    specparam_declaration12260 specparam_declaration_instance12260();
    specparam_declaration12261 specparam_declaration_instance12261();
    specparam_declaration12262 specparam_declaration_instance12262();
    specparam_declaration12263 specparam_declaration_instance12263();
    specparam_declaration12264 specparam_declaration_instance12264();
    specparam_declaration12265 specparam_declaration_instance12265();
    specparam_declaration12266 specparam_declaration_instance12266();
    specparam_declaration12267 specparam_declaration_instance12267();
    specparam_declaration12268 specparam_declaration_instance12268();
    specparam_declaration12269 specparam_declaration_instance12269();
    specparam_declaration12270 specparam_declaration_instance12270();
    specparam_declaration12271 specparam_declaration_instance12271();
    specparam_declaration12272 specparam_declaration_instance12272();
    specparam_declaration12273 specparam_declaration_instance12273();
    specparam_declaration12274 specparam_declaration_instance12274();
    specparam_declaration12275 specparam_declaration_instance12275();
    specparam_declaration12276 specparam_declaration_instance12276();
    specparam_declaration12277 specparam_declaration_instance12277();
    specparam_declaration12278 specparam_declaration_instance12278();
    specparam_declaration12279 specparam_declaration_instance12279();
    specparam_declaration12280 specparam_declaration_instance12280();
    specparam_declaration12281 specparam_declaration_instance12281();
    specparam_declaration12282 specparam_declaration_instance12282();
    specparam_declaration12283 specparam_declaration_instance12283();
    specparam_declaration12284 specparam_declaration_instance12284();
    specparam_declaration12285 specparam_declaration_instance12285();
    specparam_declaration12286 specparam_declaration_instance12286();
    specparam_declaration12287 specparam_declaration_instance12287();
    specparam_declaration12288 specparam_declaration_instance12288();
    specparam_declaration12289 specparam_declaration_instance12289();
    specparam_declaration12290 specparam_declaration_instance12290();
    specparam_declaration12291 specparam_declaration_instance12291();
    specparam_declaration12292 specparam_declaration_instance12292();
    specparam_declaration12293 specparam_declaration_instance12293();
    specparam_declaration12294 specparam_declaration_instance12294();
    specparam_declaration12295 specparam_declaration_instance12295();
    specparam_declaration12296 specparam_declaration_instance12296();
    specparam_declaration12297 specparam_declaration_instance12297();
    specparam_declaration12298 specparam_declaration_instance12298();
    specparam_declaration12299 specparam_declaration_instance12299();
    specparam_declaration12300 specparam_declaration_instance12300();
    specparam_declaration12301 specparam_declaration_instance12301();
    specparam_declaration12302 specparam_declaration_instance12302();
    specparam_declaration12303 specparam_declaration_instance12303();
    specparam_declaration12304 specparam_declaration_instance12304();
    specparam_declaration12305 specparam_declaration_instance12305();
    specparam_declaration12306 specparam_declaration_instance12306();
    specparam_declaration12307 specparam_declaration_instance12307();
    specparam_declaration12308 specparam_declaration_instance12308();
    specparam_declaration12309 specparam_declaration_instance12309();
    specparam_declaration12310 specparam_declaration_instance12310();
    specparam_declaration12311 specparam_declaration_instance12311();
    specparam_declaration12312 specparam_declaration_instance12312();
    specparam_declaration12313 specparam_declaration_instance12313();
    specparam_declaration12314 specparam_declaration_instance12314();
    specparam_declaration12315 specparam_declaration_instance12315();
    specparam_declaration12316 specparam_declaration_instance12316();
    specparam_declaration12317 specparam_declaration_instance12317();
    specparam_declaration12318 specparam_declaration_instance12318();
    specparam_declaration12319 specparam_declaration_instance12319();
    specparam_declaration12320 specparam_declaration_instance12320();
    specparam_declaration12321 specparam_declaration_instance12321();
    specparam_declaration12322 specparam_declaration_instance12322();
    specparam_declaration12323 specparam_declaration_instance12323();
    specparam_declaration12324 specparam_declaration_instance12324();
    specparam_declaration12325 specparam_declaration_instance12325();
    specparam_declaration12326 specparam_declaration_instance12326();
    specparam_declaration12327 specparam_declaration_instance12327();
    specparam_declaration12328 specparam_declaration_instance12328();
    specparam_declaration12329 specparam_declaration_instance12329();
    specparam_declaration12330 specparam_declaration_instance12330();
    specparam_declaration12331 specparam_declaration_instance12331();
    specparam_declaration12332 specparam_declaration_instance12332();
    specparam_declaration12333 specparam_declaration_instance12333();
    specparam_declaration12334 specparam_declaration_instance12334();
    specparam_declaration12335 specparam_declaration_instance12335();
    specparam_declaration12336 specparam_declaration_instance12336();
    specparam_declaration12337 specparam_declaration_instance12337();
    specparam_declaration12338 specparam_declaration_instance12338();
    specparam_declaration12339 specparam_declaration_instance12339();
    specparam_declaration12340 specparam_declaration_instance12340();
    specparam_declaration12341 specparam_declaration_instance12341();
    specparam_declaration12342 specparam_declaration_instance12342();
    specparam_declaration12343 specparam_declaration_instance12343();
    specparam_declaration12344 specparam_declaration_instance12344();
    specparam_declaration12345 specparam_declaration_instance12345();
    specparam_declaration12346 specparam_declaration_instance12346();
    specparam_declaration12347 specparam_declaration_instance12347();
    specparam_declaration12348 specparam_declaration_instance12348();
    specparam_declaration12349 specparam_declaration_instance12349();
    specparam_declaration12350 specparam_declaration_instance12350();
    specparam_declaration12351 specparam_declaration_instance12351();
    specparam_declaration12352 specparam_declaration_instance12352();
    specparam_declaration12353 specparam_declaration_instance12353();
    specparam_declaration12354 specparam_declaration_instance12354();
    specparam_declaration12355 specparam_declaration_instance12355();
    specparam_declaration12356 specparam_declaration_instance12356();
    specparam_declaration12357 specparam_declaration_instance12357();
    specparam_declaration12358 specparam_declaration_instance12358();
    specparam_declaration12359 specparam_declaration_instance12359();
    specparam_declaration12360 specparam_declaration_instance12360();
    specparam_declaration12361 specparam_declaration_instance12361();
    specparam_declaration12362 specparam_declaration_instance12362();
    specparam_declaration12363 specparam_declaration_instance12363();
    specparam_declaration12364 specparam_declaration_instance12364();
    specparam_declaration12365 specparam_declaration_instance12365();
    specparam_declaration12366 specparam_declaration_instance12366();
    specparam_declaration12367 specparam_declaration_instance12367();
    specparam_declaration12368 specparam_declaration_instance12368();
    specparam_declaration12369 specparam_declaration_instance12369();
    specparam_declaration12370 specparam_declaration_instance12370();
    specparam_declaration12371 specparam_declaration_instance12371();
    specparam_declaration12372 specparam_declaration_instance12372();
    specparam_declaration12373 specparam_declaration_instance12373();
    specparam_declaration12374 specparam_declaration_instance12374();
    specparam_declaration12375 specparam_declaration_instance12375();
    specparam_declaration12376 specparam_declaration_instance12376();
    specparam_declaration12377 specparam_declaration_instance12377();
    specparam_declaration12378 specparam_declaration_instance12378();
    specparam_declaration12379 specparam_declaration_instance12379();
    specparam_declaration12380 specparam_declaration_instance12380();
    specparam_declaration12381 specparam_declaration_instance12381();
    specparam_declaration12382 specparam_declaration_instance12382();
    specparam_declaration12383 specparam_declaration_instance12383();
    specparam_declaration12384 specparam_declaration_instance12384();
    specparam_declaration12385 specparam_declaration_instance12385();
    specparam_declaration12386 specparam_declaration_instance12386();
    specparam_declaration12387 specparam_declaration_instance12387();
    specparam_declaration12388 specparam_declaration_instance12388();
    specparam_declaration12389 specparam_declaration_instance12389();
    specparam_declaration12390 specparam_declaration_instance12390();
    specparam_declaration12391 specparam_declaration_instance12391();
    specparam_declaration12392 specparam_declaration_instance12392();
    specparam_declaration12393 specparam_declaration_instance12393();
    specparam_declaration12394 specparam_declaration_instance12394();
    specparam_declaration12395 specparam_declaration_instance12395();
    specparam_declaration12396 specparam_declaration_instance12396();
    specparam_declaration12397 specparam_declaration_instance12397();
    specparam_declaration12398 specparam_declaration_instance12398();
    specparam_declaration12399 specparam_declaration_instance12399();
    specparam_declaration12400 specparam_declaration_instance12400();
    specparam_declaration12401 specparam_declaration_instance12401();
    specparam_declaration12402 specparam_declaration_instance12402();
    specparam_declaration12403 specparam_declaration_instance12403();
    specparam_declaration12404 specparam_declaration_instance12404();
    specparam_declaration12405 specparam_declaration_instance12405();
    specparam_declaration12406 specparam_declaration_instance12406();
    specparam_declaration12407 specparam_declaration_instance12407();
    specparam_declaration12408 specparam_declaration_instance12408();
    specparam_declaration12409 specparam_declaration_instance12409();
    specparam_declaration12410 specparam_declaration_instance12410();
    specparam_declaration12411 specparam_declaration_instance12411();
    specparam_declaration12412 specparam_declaration_instance12412();
    specparam_declaration12413 specparam_declaration_instance12413();
    specparam_declaration12414 specparam_declaration_instance12414();
    specparam_declaration12415 specparam_declaration_instance12415();
    specparam_declaration12416 specparam_declaration_instance12416();
    specparam_declaration12417 specparam_declaration_instance12417();
    specparam_declaration12418 specparam_declaration_instance12418();
    specparam_declaration12419 specparam_declaration_instance12419();
    specparam_declaration12420 specparam_declaration_instance12420();
    specparam_declaration12421 specparam_declaration_instance12421();
    specparam_declaration12422 specparam_declaration_instance12422();
    specparam_declaration12423 specparam_declaration_instance12423();
    specparam_declaration12424 specparam_declaration_instance12424();
    specparam_declaration12425 specparam_declaration_instance12425();
    specparam_declaration12426 specparam_declaration_instance12426();
    specparam_declaration12427 specparam_declaration_instance12427();
    specparam_declaration12428 specparam_declaration_instance12428();
    specparam_declaration12429 specparam_declaration_instance12429();
    specparam_declaration12430 specparam_declaration_instance12430();
    specparam_declaration12431 specparam_declaration_instance12431();
    specparam_declaration12432 specparam_declaration_instance12432();
    specparam_declaration12433 specparam_declaration_instance12433();
    specparam_declaration12434 specparam_declaration_instance12434();
    specparam_declaration12435 specparam_declaration_instance12435();
    specparam_declaration12436 specparam_declaration_instance12436();
    specparam_declaration12437 specparam_declaration_instance12437();
    specparam_declaration12438 specparam_declaration_instance12438();
    specparam_declaration12439 specparam_declaration_instance12439();
    specparam_declaration12440 specparam_declaration_instance12440();
    specparam_declaration12441 specparam_declaration_instance12441();
    specparam_declaration12442 specparam_declaration_instance12442();
    specparam_declaration12443 specparam_declaration_instance12443();
    specparam_declaration12444 specparam_declaration_instance12444();
    specparam_declaration12445 specparam_declaration_instance12445();
    specparam_declaration12446 specparam_declaration_instance12446();
    specparam_declaration12447 specparam_declaration_instance12447();
    specparam_declaration12448 specparam_declaration_instance12448();
    specparam_declaration12449 specparam_declaration_instance12449();
    specparam_declaration12450 specparam_declaration_instance12450();
    specparam_declaration12451 specparam_declaration_instance12451();
    specparam_declaration12452 specparam_declaration_instance12452();
    specparam_declaration12453 specparam_declaration_instance12453();
    specparam_declaration12454 specparam_declaration_instance12454();
    specparam_declaration12455 specparam_declaration_instance12455();
    specparam_declaration12456 specparam_declaration_instance12456();
    specparam_declaration12457 specparam_declaration_instance12457();
    specparam_declaration12458 specparam_declaration_instance12458();
    specparam_declaration12459 specparam_declaration_instance12459();
    specparam_declaration12460 specparam_declaration_instance12460();
    specparam_declaration12461 specparam_declaration_instance12461();
    specparam_declaration12462 specparam_declaration_instance12462();
    specparam_declaration12463 specparam_declaration_instance12463();
    specparam_declaration12464 specparam_declaration_instance12464();
    specparam_declaration12465 specparam_declaration_instance12465();
    specparam_declaration12466 specparam_declaration_instance12466();
    specparam_declaration12467 specparam_declaration_instance12467();
    specparam_declaration12468 specparam_declaration_instance12468();
    specparam_declaration12469 specparam_declaration_instance12469();
    specparam_declaration12470 specparam_declaration_instance12470();
    specparam_declaration12471 specparam_declaration_instance12471();
    specparam_declaration12472 specparam_declaration_instance12472();
    specparam_declaration12473 specparam_declaration_instance12473();
    specparam_declaration12474 specparam_declaration_instance12474();
    specparam_declaration12475 specparam_declaration_instance12475();
    specparam_declaration12476 specparam_declaration_instance12476();
    specparam_declaration12477 specparam_declaration_instance12477();
    specparam_declaration12478 specparam_declaration_instance12478();
    specparam_declaration12479 specparam_declaration_instance12479();
    specparam_declaration12480 specparam_declaration_instance12480();
    specparam_declaration12481 specparam_declaration_instance12481();
    specparam_declaration12482 specparam_declaration_instance12482();
    specparam_declaration12483 specparam_declaration_instance12483();
    specparam_declaration12484 specparam_declaration_instance12484();
    specparam_declaration12485 specparam_declaration_instance12485();
    specparam_declaration12486 specparam_declaration_instance12486();
    specparam_declaration12487 specparam_declaration_instance12487();
    specparam_declaration12488 specparam_declaration_instance12488();
    specparam_declaration12489 specparam_declaration_instance12489();
    specparam_declaration12490 specparam_declaration_instance12490();
    specparam_declaration12491 specparam_declaration_instance12491();
    specparam_declaration12492 specparam_declaration_instance12492();
    specparam_declaration12493 specparam_declaration_instance12493();
    specparam_declaration12494 specparam_declaration_instance12494();
    specparam_declaration12495 specparam_declaration_instance12495();
    specparam_declaration12496 specparam_declaration_instance12496();
    specparam_declaration12497 specparam_declaration_instance12497();
    specparam_declaration12498 specparam_declaration_instance12498();
    specparam_declaration12499 specparam_declaration_instance12499();
    specparam_declaration12500 specparam_declaration_instance12500();
    specparam_declaration12501 specparam_declaration_instance12501();
    specparam_declaration12502 specparam_declaration_instance12502();
    specparam_declaration12503 specparam_declaration_instance12503();
    specparam_declaration12504 specparam_declaration_instance12504();
    specparam_declaration12505 specparam_declaration_instance12505();
    specparam_declaration12506 specparam_declaration_instance12506();
    specparam_declaration12507 specparam_declaration_instance12507();
    specparam_declaration12508 specparam_declaration_instance12508();
    specparam_declaration12509 specparam_declaration_instance12509();
    specparam_declaration12510 specparam_declaration_instance12510();
    specparam_declaration12511 specparam_declaration_instance12511();
    specparam_declaration12512 specparam_declaration_instance12512();
    specparam_declaration12513 specparam_declaration_instance12513();
    specparam_declaration12514 specparam_declaration_instance12514();
    specparam_declaration12515 specparam_declaration_instance12515();
    specparam_declaration12516 specparam_declaration_instance12516();
    specparam_declaration12517 specparam_declaration_instance12517();
    specparam_declaration12518 specparam_declaration_instance12518();
    specparam_declaration12519 specparam_declaration_instance12519();
    specparam_declaration12520 specparam_declaration_instance12520();
    specparam_declaration12521 specparam_declaration_instance12521();
    specparam_declaration12522 specparam_declaration_instance12522();
    specparam_declaration12523 specparam_declaration_instance12523();
    specparam_declaration12524 specparam_declaration_instance12524();
    specparam_declaration12525 specparam_declaration_instance12525();
    specparam_declaration12526 specparam_declaration_instance12526();
    specparam_declaration12527 specparam_declaration_instance12527();
    specparam_declaration12528 specparam_declaration_instance12528();
    specparam_declaration12529 specparam_declaration_instance12529();
    specparam_declaration12530 specparam_declaration_instance12530();
    specparam_declaration12531 specparam_declaration_instance12531();
    specparam_declaration12532 specparam_declaration_instance12532();
    specparam_declaration12533 specparam_declaration_instance12533();
    specparam_declaration12534 specparam_declaration_instance12534();
    specparam_declaration12535 specparam_declaration_instance12535();
    specparam_declaration12536 specparam_declaration_instance12536();
    specparam_declaration12537 specparam_declaration_instance12537();
    specparam_declaration12538 specparam_declaration_instance12538();
    specparam_declaration12539 specparam_declaration_instance12539();
    specparam_declaration12540 specparam_declaration_instance12540();
    specparam_declaration12541 specparam_declaration_instance12541();
    specparam_declaration12542 specparam_declaration_instance12542();
    specparam_declaration12543 specparam_declaration_instance12543();
    specparam_declaration12544 specparam_declaration_instance12544();
    specparam_declaration12545 specparam_declaration_instance12545();
    specparam_declaration12546 specparam_declaration_instance12546();
    specparam_declaration12547 specparam_declaration_instance12547();
    specparam_declaration12548 specparam_declaration_instance12548();
    specparam_declaration12549 specparam_declaration_instance12549();
    specparam_declaration12550 specparam_declaration_instance12550();
    specparam_declaration12551 specparam_declaration_instance12551();
    specparam_declaration12552 specparam_declaration_instance12552();
    specparam_declaration12553 specparam_declaration_instance12553();
    specparam_declaration12554 specparam_declaration_instance12554();
    specparam_declaration12555 specparam_declaration_instance12555();
    specparam_declaration12556 specparam_declaration_instance12556();
    specparam_declaration12557 specparam_declaration_instance12557();
    specparam_declaration12558 specparam_declaration_instance12558();
    specparam_declaration12559 specparam_declaration_instance12559();
    specparam_declaration12560 specparam_declaration_instance12560();
    specparam_declaration12561 specparam_declaration_instance12561();
    specparam_declaration12562 specparam_declaration_instance12562();
    specparam_declaration12563 specparam_declaration_instance12563();
    specparam_declaration12564 specparam_declaration_instance12564();
    specparam_declaration12565 specparam_declaration_instance12565();
    specparam_declaration12566 specparam_declaration_instance12566();
    specparam_declaration12567 specparam_declaration_instance12567();
    specparam_declaration12568 specparam_declaration_instance12568();
    specparam_declaration12569 specparam_declaration_instance12569();
    specparam_declaration12570 specparam_declaration_instance12570();
    specparam_declaration12571 specparam_declaration_instance12571();
    specparam_declaration12572 specparam_declaration_instance12572();
    specparam_declaration12573 specparam_declaration_instance12573();
    specparam_declaration12574 specparam_declaration_instance12574();
    specparam_declaration12575 specparam_declaration_instance12575();
    specparam_declaration12576 specparam_declaration_instance12576();
    specparam_declaration12577 specparam_declaration_instance12577();
    specparam_declaration12578 specparam_declaration_instance12578();
    specparam_declaration12579 specparam_declaration_instance12579();
    specparam_declaration12580 specparam_declaration_instance12580();
    specparam_declaration12581 specparam_declaration_instance12581();
    specparam_declaration12582 specparam_declaration_instance12582();
    specparam_declaration12583 specparam_declaration_instance12583();
    specparam_declaration12584 specparam_declaration_instance12584();
    specparam_declaration12585 specparam_declaration_instance12585();
    specparam_declaration12586 specparam_declaration_instance12586();
    specparam_declaration12587 specparam_declaration_instance12587();
    specparam_declaration12588 specparam_declaration_instance12588();
    specparam_declaration12589 specparam_declaration_instance12589();
    specparam_declaration12590 specparam_declaration_instance12590();
    specparam_declaration12591 specparam_declaration_instance12591();
    specparam_declaration12592 specparam_declaration_instance12592();
    specparam_declaration12593 specparam_declaration_instance12593();
    specparam_declaration12594 specparam_declaration_instance12594();
    specparam_declaration12595 specparam_declaration_instance12595();
    specparam_declaration12596 specparam_declaration_instance12596();
    specparam_declaration12597 specparam_declaration_instance12597();
    specparam_declaration12598 specparam_declaration_instance12598();
    specparam_declaration12599 specparam_declaration_instance12599();
    specparam_declaration12600 specparam_declaration_instance12600();
    specparam_declaration12601 specparam_declaration_instance12601();
    specparam_declaration12602 specparam_declaration_instance12602();
    specparam_declaration12603 specparam_declaration_instance12603();
    specparam_declaration12604 specparam_declaration_instance12604();
    specparam_declaration12605 specparam_declaration_instance12605();
    specparam_declaration12606 specparam_declaration_instance12606();
    specparam_declaration12607 specparam_declaration_instance12607();
    specparam_declaration12608 specparam_declaration_instance12608();
    specparam_declaration12609 specparam_declaration_instance12609();
    specparam_declaration12610 specparam_declaration_instance12610();
    specparam_declaration12611 specparam_declaration_instance12611();
    specparam_declaration12612 specparam_declaration_instance12612();
    specparam_declaration12613 specparam_declaration_instance12613();
    specparam_declaration12614 specparam_declaration_instance12614();
    specparam_declaration12615 specparam_declaration_instance12615();
    specparam_declaration12616 specparam_declaration_instance12616();
    specparam_declaration12617 specparam_declaration_instance12617();
    specparam_declaration12618 specparam_declaration_instance12618();
    specparam_declaration12619 specparam_declaration_instance12619();
    specparam_declaration12620 specparam_declaration_instance12620();
    specparam_declaration12621 specparam_declaration_instance12621();
    specparam_declaration12622 specparam_declaration_instance12622();
    specparam_declaration12623 specparam_declaration_instance12623();
    specparam_declaration12624 specparam_declaration_instance12624();
    specparam_declaration12625 specparam_declaration_instance12625();
    specparam_declaration12626 specparam_declaration_instance12626();
    specparam_declaration12627 specparam_declaration_instance12627();
    specparam_declaration12628 specparam_declaration_instance12628();
    specparam_declaration12629 specparam_declaration_instance12629();
    specparam_declaration12630 specparam_declaration_instance12630();
    specparam_declaration12631 specparam_declaration_instance12631();
    specparam_declaration12632 specparam_declaration_instance12632();
    specparam_declaration12633 specparam_declaration_instance12633();
    specparam_declaration12634 specparam_declaration_instance12634();
    specparam_declaration12635 specparam_declaration_instance12635();
    specparam_declaration12636 specparam_declaration_instance12636();
    specparam_declaration12637 specparam_declaration_instance12637();
    specparam_declaration12638 specparam_declaration_instance12638();
    specparam_declaration12639 specparam_declaration_instance12639();
    specparam_declaration12640 specparam_declaration_instance12640();
    specparam_declaration12641 specparam_declaration_instance12641();
    specparam_declaration12642 specparam_declaration_instance12642();
    specparam_declaration12643 specparam_declaration_instance12643();
    specparam_declaration12644 specparam_declaration_instance12644();
    specparam_declaration12645 specparam_declaration_instance12645();
    specparam_declaration12646 specparam_declaration_instance12646();
    specparam_declaration12647 specparam_declaration_instance12647();
    specparam_declaration12648 specparam_declaration_instance12648();
    specparam_declaration12649 specparam_declaration_instance12649();
    specparam_declaration12650 specparam_declaration_instance12650();
    specparam_declaration12651 specparam_declaration_instance12651();
    specparam_declaration12652 specparam_declaration_instance12652();
    specparam_declaration12653 specparam_declaration_instance12653();
    specparam_declaration12654 specparam_declaration_instance12654();
    specparam_declaration12655 specparam_declaration_instance12655();
    specparam_declaration12656 specparam_declaration_instance12656();
    specparam_declaration12657 specparam_declaration_instance12657();
    specparam_declaration12658 specparam_declaration_instance12658();
    specparam_declaration12659 specparam_declaration_instance12659();
    specparam_declaration12660 specparam_declaration_instance12660();
    specparam_declaration12661 specparam_declaration_instance12661();
    specparam_declaration12662 specparam_declaration_instance12662();
    specparam_declaration12663 specparam_declaration_instance12663();
    specparam_declaration12664 specparam_declaration_instance12664();
    specparam_declaration12665 specparam_declaration_instance12665();
    specparam_declaration12666 specparam_declaration_instance12666();
    specparam_declaration12667 specparam_declaration_instance12667();
    specparam_declaration12668 specparam_declaration_instance12668();
    specparam_declaration12669 specparam_declaration_instance12669();
    specparam_declaration12670 specparam_declaration_instance12670();
    specparam_declaration12671 specparam_declaration_instance12671();
    specparam_declaration12672 specparam_declaration_instance12672();
    specparam_declaration12673 specparam_declaration_instance12673();
    specparam_declaration12674 specparam_declaration_instance12674();
    specparam_declaration12675 specparam_declaration_instance12675();
    specparam_declaration12676 specparam_declaration_instance12676();
    specparam_declaration12677 specparam_declaration_instance12677();
    specparam_declaration12678 specparam_declaration_instance12678();
    specparam_declaration12679 specparam_declaration_instance12679();
    specparam_declaration12680 specparam_declaration_instance12680();
    specparam_declaration12681 specparam_declaration_instance12681();
    specparam_declaration12682 specparam_declaration_instance12682();
    specparam_declaration12683 specparam_declaration_instance12683();
    specparam_declaration12684 specparam_declaration_instance12684();
    specparam_declaration12685 specparam_declaration_instance12685();
    specparam_declaration12686 specparam_declaration_instance12686();
    specparam_declaration12687 specparam_declaration_instance12687();
    specparam_declaration12688 specparam_declaration_instance12688();
    specparam_declaration12689 specparam_declaration_instance12689();
    specparam_declaration12690 specparam_declaration_instance12690();
    specparam_declaration12691 specparam_declaration_instance12691();
    specparam_declaration12692 specparam_declaration_instance12692();
    specparam_declaration12693 specparam_declaration_instance12693();
    specparam_declaration12694 specparam_declaration_instance12694();
    specparam_declaration12695 specparam_declaration_instance12695();
    specparam_declaration12696 specparam_declaration_instance12696();
    specparam_declaration12697 specparam_declaration_instance12697();
    specparam_declaration12698 specparam_declaration_instance12698();
    specparam_declaration12699 specparam_declaration_instance12699();
    specparam_declaration12700 specparam_declaration_instance12700();
    specparam_declaration12701 specparam_declaration_instance12701();
    specparam_declaration12702 specparam_declaration_instance12702();
    specparam_declaration12703 specparam_declaration_instance12703();
    specparam_declaration12704 specparam_declaration_instance12704();
    specparam_declaration12705 specparam_declaration_instance12705();
    specparam_declaration12706 specparam_declaration_instance12706();
    specparam_declaration12707 specparam_declaration_instance12707();
    specparam_declaration12708 specparam_declaration_instance12708();
    specparam_declaration12709 specparam_declaration_instance12709();
    specparam_declaration12710 specparam_declaration_instance12710();
    specparam_declaration12711 specparam_declaration_instance12711();
    specparam_declaration12712 specparam_declaration_instance12712();
    specparam_declaration12713 specparam_declaration_instance12713();
    specparam_declaration12714 specparam_declaration_instance12714();
    specparam_declaration12715 specparam_declaration_instance12715();
    specparam_declaration12716 specparam_declaration_instance12716();
    specparam_declaration12717 specparam_declaration_instance12717();
    specparam_declaration12718 specparam_declaration_instance12718();
    specparam_declaration12719 specparam_declaration_instance12719();
    specparam_declaration12720 specparam_declaration_instance12720();
    specparam_declaration12721 specparam_declaration_instance12721();
    specparam_declaration12722 specparam_declaration_instance12722();
    specparam_declaration12723 specparam_declaration_instance12723();
    specparam_declaration12724 specparam_declaration_instance12724();
    specparam_declaration12725 specparam_declaration_instance12725();
    specparam_declaration12726 specparam_declaration_instance12726();
    specparam_declaration12727 specparam_declaration_instance12727();
    specparam_declaration12728 specparam_declaration_instance12728();
    specparam_declaration12729 specparam_declaration_instance12729();
    specparam_declaration12730 specparam_declaration_instance12730();
    specparam_declaration12731 specparam_declaration_instance12731();
    specparam_declaration12732 specparam_declaration_instance12732();
    specparam_declaration12733 specparam_declaration_instance12733();
    specparam_declaration12734 specparam_declaration_instance12734();
    specparam_declaration12735 specparam_declaration_instance12735();
    specparam_declaration12736 specparam_declaration_instance12736();
    specparam_declaration12737 specparam_declaration_instance12737();
    specparam_declaration12738 specparam_declaration_instance12738();
    specparam_declaration12739 specparam_declaration_instance12739();
    specparam_declaration12740 specparam_declaration_instance12740();
    specparam_declaration12741 specparam_declaration_instance12741();
    specparam_declaration12742 specparam_declaration_instance12742();
    specparam_declaration12743 specparam_declaration_instance12743();
    specparam_declaration12744 specparam_declaration_instance12744();
    specparam_declaration12745 specparam_declaration_instance12745();
    specparam_declaration12746 specparam_declaration_instance12746();
    specparam_declaration12747 specparam_declaration_instance12747();
    specparam_declaration12748 specparam_declaration_instance12748();
    specparam_declaration12749 specparam_declaration_instance12749();
    specparam_declaration12750 specparam_declaration_instance12750();
    specparam_declaration12751 specparam_declaration_instance12751();
    specparam_declaration12752 specparam_declaration_instance12752();
    specparam_declaration12753 specparam_declaration_instance12753();
    specparam_declaration12754 specparam_declaration_instance12754();
    specparam_declaration12755 specparam_declaration_instance12755();
    specparam_declaration12756 specparam_declaration_instance12756();
    specparam_declaration12757 specparam_declaration_instance12757();
    specparam_declaration12758 specparam_declaration_instance12758();
    specparam_declaration12759 specparam_declaration_instance12759();
    specparam_declaration12760 specparam_declaration_instance12760();
    specparam_declaration12761 specparam_declaration_instance12761();
    specparam_declaration12762 specparam_declaration_instance12762();
    specparam_declaration12763 specparam_declaration_instance12763();
    specparam_declaration12764 specparam_declaration_instance12764();
    specparam_declaration12765 specparam_declaration_instance12765();
    specparam_declaration12766 specparam_declaration_instance12766();
    specparam_declaration12767 specparam_declaration_instance12767();
    specparam_declaration12768 specparam_declaration_instance12768();
    specparam_declaration12769 specparam_declaration_instance12769();
    specparam_declaration12770 specparam_declaration_instance12770();
    specparam_declaration12771 specparam_declaration_instance12771();
    specparam_declaration12772 specparam_declaration_instance12772();
    specparam_declaration12773 specparam_declaration_instance12773();
    specparam_declaration12774 specparam_declaration_instance12774();
    specparam_declaration12775 specparam_declaration_instance12775();
    specparam_declaration12776 specparam_declaration_instance12776();
    specparam_declaration12777 specparam_declaration_instance12777();
    specparam_declaration12778 specparam_declaration_instance12778();
    specparam_declaration12779 specparam_declaration_instance12779();
    specparam_declaration12780 specparam_declaration_instance12780();
    specparam_declaration12781 specparam_declaration_instance12781();
    specparam_declaration12782 specparam_declaration_instance12782();
    specparam_declaration12783 specparam_declaration_instance12783();
    specparam_declaration12784 specparam_declaration_instance12784();
    specparam_declaration12785 specparam_declaration_instance12785();
    specparam_declaration12786 specparam_declaration_instance12786();
    specparam_declaration12787 specparam_declaration_instance12787();
    specparam_declaration12788 specparam_declaration_instance12788();
    specparam_declaration12789 specparam_declaration_instance12789();
    specparam_declaration12790 specparam_declaration_instance12790();
    specparam_declaration12791 specparam_declaration_instance12791();
    specparam_declaration12792 specparam_declaration_instance12792();
    specparam_declaration12793 specparam_declaration_instance12793();
    specparam_declaration12794 specparam_declaration_instance12794();
    specparam_declaration12795 specparam_declaration_instance12795();
    specparam_declaration12796 specparam_declaration_instance12796();
    specparam_declaration12797 specparam_declaration_instance12797();
    specparam_declaration12798 specparam_declaration_instance12798();
    specparam_declaration12799 specparam_declaration_instance12799();
    specparam_declaration12800 specparam_declaration_instance12800();
    specparam_declaration12801 specparam_declaration_instance12801();
    specparam_declaration12802 specparam_declaration_instance12802();
    specparam_declaration12803 specparam_declaration_instance12803();
    specparam_declaration12804 specparam_declaration_instance12804();
    specparam_declaration12805 specparam_declaration_instance12805();
    specparam_declaration12806 specparam_declaration_instance12806();
    specparam_declaration12807 specparam_declaration_instance12807();
    specparam_declaration12808 specparam_declaration_instance12808();
    specparam_declaration12809 specparam_declaration_instance12809();
    specparam_declaration12810 specparam_declaration_instance12810();
    specparam_declaration12811 specparam_declaration_instance12811();
    specparam_declaration12812 specparam_declaration_instance12812();
    specparam_declaration12813 specparam_declaration_instance12813();
    specparam_declaration12814 specparam_declaration_instance12814();
    specparam_declaration12815 specparam_declaration_instance12815();
    specparam_declaration12816 specparam_declaration_instance12816();
    specparam_declaration12817 specparam_declaration_instance12817();
    specparam_declaration12818 specparam_declaration_instance12818();
    specparam_declaration12819 specparam_declaration_instance12819();
    specparam_declaration12820 specparam_declaration_instance12820();
    specparam_declaration12821 specparam_declaration_instance12821();
    specparam_declaration12822 specparam_declaration_instance12822();
    specparam_declaration12823 specparam_declaration_instance12823();
    specparam_declaration12824 specparam_declaration_instance12824();
    specparam_declaration12825 specparam_declaration_instance12825();
    specparam_declaration12826 specparam_declaration_instance12826();
    specparam_declaration12827 specparam_declaration_instance12827();
    specparam_declaration12828 specparam_declaration_instance12828();
    specparam_declaration12829 specparam_declaration_instance12829();
    specparam_declaration12830 specparam_declaration_instance12830();
    specparam_declaration12831 specparam_declaration_instance12831();
    specparam_declaration12832 specparam_declaration_instance12832();
    specparam_declaration12833 specparam_declaration_instance12833();
    specparam_declaration12834 specparam_declaration_instance12834();
    specparam_declaration12835 specparam_declaration_instance12835();
    specparam_declaration12836 specparam_declaration_instance12836();
    specparam_declaration12837 specparam_declaration_instance12837();
    specparam_declaration12838 specparam_declaration_instance12838();
    specparam_declaration12839 specparam_declaration_instance12839();
    specparam_declaration12840 specparam_declaration_instance12840();
    specparam_declaration12841 specparam_declaration_instance12841();
    specparam_declaration12842 specparam_declaration_instance12842();
    specparam_declaration12843 specparam_declaration_instance12843();
    specparam_declaration12844 specparam_declaration_instance12844();
    specparam_declaration12845 specparam_declaration_instance12845();
    specparam_declaration12846 specparam_declaration_instance12846();
    specparam_declaration12847 specparam_declaration_instance12847();
    specparam_declaration12848 specparam_declaration_instance12848();
    specparam_declaration12849 specparam_declaration_instance12849();
    specparam_declaration12850 specparam_declaration_instance12850();
    specparam_declaration12851 specparam_declaration_instance12851();
    specparam_declaration12852 specparam_declaration_instance12852();
    specparam_declaration12853 specparam_declaration_instance12853();
    specparam_declaration12854 specparam_declaration_instance12854();
    specparam_declaration12855 specparam_declaration_instance12855();
    specparam_declaration12856 specparam_declaration_instance12856();
    specparam_declaration12857 specparam_declaration_instance12857();
    specparam_declaration12858 specparam_declaration_instance12858();
    specparam_declaration12859 specparam_declaration_instance12859();
    specparam_declaration12860 specparam_declaration_instance12860();
    specparam_declaration12861 specparam_declaration_instance12861();
    specparam_declaration12862 specparam_declaration_instance12862();
    specparam_declaration12863 specparam_declaration_instance12863();
    specparam_declaration12864 specparam_declaration_instance12864();
    specparam_declaration12865 specparam_declaration_instance12865();
    specparam_declaration12866 specparam_declaration_instance12866();
    specparam_declaration12867 specparam_declaration_instance12867();
    specparam_declaration12868 specparam_declaration_instance12868();
    specparam_declaration12869 specparam_declaration_instance12869();
    specparam_declaration12870 specparam_declaration_instance12870();
    specparam_declaration12871 specparam_declaration_instance12871();
    specparam_declaration12872 specparam_declaration_instance12872();
    specparam_declaration12873 specparam_declaration_instance12873();
    specparam_declaration12874 specparam_declaration_instance12874();
    specparam_declaration12875 specparam_declaration_instance12875();
    specparam_declaration12876 specparam_declaration_instance12876();
    specparam_declaration12877 specparam_declaration_instance12877();
    specparam_declaration12878 specparam_declaration_instance12878();
    specparam_declaration12879 specparam_declaration_instance12879();
    specparam_declaration12880 specparam_declaration_instance12880();
    specparam_declaration12881 specparam_declaration_instance12881();
    specparam_declaration12882 specparam_declaration_instance12882();
    specparam_declaration12883 specparam_declaration_instance12883();
    specparam_declaration12884 specparam_declaration_instance12884();
    specparam_declaration12885 specparam_declaration_instance12885();
    specparam_declaration12886 specparam_declaration_instance12886();
    specparam_declaration12887 specparam_declaration_instance12887();
    specparam_declaration12888 specparam_declaration_instance12888();
    specparam_declaration12889 specparam_declaration_instance12889();
    specparam_declaration12890 specparam_declaration_instance12890();
    specparam_declaration12891 specparam_declaration_instance12891();
    specparam_declaration12892 specparam_declaration_instance12892();
    specparam_declaration12893 specparam_declaration_instance12893();
    specparam_declaration12894 specparam_declaration_instance12894();
    specparam_declaration12895 specparam_declaration_instance12895();
    specparam_declaration12896 specparam_declaration_instance12896();
    specparam_declaration12897 specparam_declaration_instance12897();
    specparam_declaration12898 specparam_declaration_instance12898();
    specparam_declaration12899 specparam_declaration_instance12899();
    specparam_declaration12900 specparam_declaration_instance12900();
    specparam_declaration12901 specparam_declaration_instance12901();
    specparam_declaration12902 specparam_declaration_instance12902();
    specparam_declaration12903 specparam_declaration_instance12903();
    specparam_declaration12904 specparam_declaration_instance12904();
    specparam_declaration12905 specparam_declaration_instance12905();
    specparam_declaration12906 specparam_declaration_instance12906();
    specparam_declaration12907 specparam_declaration_instance12907();
    specparam_declaration12908 specparam_declaration_instance12908();
    specparam_declaration12909 specparam_declaration_instance12909();
    specparam_declaration12910 specparam_declaration_instance12910();
    specparam_declaration12911 specparam_declaration_instance12911();
    specparam_declaration12912 specparam_declaration_instance12912();
    specparam_declaration12913 specparam_declaration_instance12913();
    specparam_declaration12914 specparam_declaration_instance12914();
    specparam_declaration12915 specparam_declaration_instance12915();
    specparam_declaration12916 specparam_declaration_instance12916();
    specparam_declaration12917 specparam_declaration_instance12917();
    specparam_declaration12918 specparam_declaration_instance12918();
    specparam_declaration12919 specparam_declaration_instance12919();
    specparam_declaration12920 specparam_declaration_instance12920();
    specparam_declaration12921 specparam_declaration_instance12921();
    specparam_declaration12922 specparam_declaration_instance12922();
    specparam_declaration12923 specparam_declaration_instance12923();
    specparam_declaration12924 specparam_declaration_instance12924();
    specparam_declaration12925 specparam_declaration_instance12925();
    specparam_declaration12926 specparam_declaration_instance12926();
    specparam_declaration12927 specparam_declaration_instance12927();
    specparam_declaration12928 specparam_declaration_instance12928();
    specparam_declaration12929 specparam_declaration_instance12929();
    specparam_declaration12930 specparam_declaration_instance12930();
    specparam_declaration12931 specparam_declaration_instance12931();
    specparam_declaration12932 specparam_declaration_instance12932();
    specparam_declaration12933 specparam_declaration_instance12933();
    specparam_declaration12934 specparam_declaration_instance12934();
    specparam_declaration12935 specparam_declaration_instance12935();
    specparam_declaration12936 specparam_declaration_instance12936();
    specparam_declaration12937 specparam_declaration_instance12937();
    specparam_declaration12938 specparam_declaration_instance12938();
    specparam_declaration12939 specparam_declaration_instance12939();
    specparam_declaration12940 specparam_declaration_instance12940();
    specparam_declaration12941 specparam_declaration_instance12941();
    specparam_declaration12942 specparam_declaration_instance12942();
    specparam_declaration12943 specparam_declaration_instance12943();
    specparam_declaration12944 specparam_declaration_instance12944();
    specparam_declaration12945 specparam_declaration_instance12945();
    specparam_declaration12946 specparam_declaration_instance12946();
    specparam_declaration12947 specparam_declaration_instance12947();
    specparam_declaration12948 specparam_declaration_instance12948();
    specparam_declaration12949 specparam_declaration_instance12949();
    specparam_declaration12950 specparam_declaration_instance12950();
    specparam_declaration12951 specparam_declaration_instance12951();
    specparam_declaration12952 specparam_declaration_instance12952();
    specparam_declaration12953 specparam_declaration_instance12953();
    specparam_declaration12954 specparam_declaration_instance12954();
    specparam_declaration12955 specparam_declaration_instance12955();
    specparam_declaration12956 specparam_declaration_instance12956();
    specparam_declaration12957 specparam_declaration_instance12957();
    specparam_declaration12958 specparam_declaration_instance12958();
    specparam_declaration12959 specparam_declaration_instance12959();
    specparam_declaration12960 specparam_declaration_instance12960();
    specparam_declaration12961 specparam_declaration_instance12961();
    specparam_declaration12962 specparam_declaration_instance12962();
    specparam_declaration12963 specparam_declaration_instance12963();
    specparam_declaration12964 specparam_declaration_instance12964();
    specparam_declaration12965 specparam_declaration_instance12965();
    specparam_declaration12966 specparam_declaration_instance12966();
    specparam_declaration12967 specparam_declaration_instance12967();
    specparam_declaration12968 specparam_declaration_instance12968();
    specparam_declaration12969 specparam_declaration_instance12969();
    specparam_declaration12970 specparam_declaration_instance12970();
    specparam_declaration12971 specparam_declaration_instance12971();
    specparam_declaration12972 specparam_declaration_instance12972();
    specparam_declaration12973 specparam_declaration_instance12973();
    specparam_declaration12974 specparam_declaration_instance12974();
    specparam_declaration12975 specparam_declaration_instance12975();
    specparam_declaration12976 specparam_declaration_instance12976();
    specparam_declaration12977 specparam_declaration_instance12977();
    specparam_declaration12978 specparam_declaration_instance12978();
    specparam_declaration12979 specparam_declaration_instance12979();
    specparam_declaration12980 specparam_declaration_instance12980();
    specparam_declaration12981 specparam_declaration_instance12981();
    specparam_declaration12982 specparam_declaration_instance12982();
    specparam_declaration12983 specparam_declaration_instance12983();
    specparam_declaration12984 specparam_declaration_instance12984();
    specparam_declaration12985 specparam_declaration_instance12985();
    specparam_declaration12986 specparam_declaration_instance12986();
    specparam_declaration12987 specparam_declaration_instance12987();
    specparam_declaration12988 specparam_declaration_instance12988();
    specparam_declaration12989 specparam_declaration_instance12989();
    specparam_declaration12990 specparam_declaration_instance12990();
    specparam_declaration12991 specparam_declaration_instance12991();
    specparam_declaration12992 specparam_declaration_instance12992();
    specparam_declaration12993 specparam_declaration_instance12993();
    specparam_declaration12994 specparam_declaration_instance12994();
    specparam_declaration12995 specparam_declaration_instance12995();
    specparam_declaration12996 specparam_declaration_instance12996();
    specparam_declaration12997 specparam_declaration_instance12997();
    specparam_declaration12998 specparam_declaration_instance12998();
    specparam_declaration12999 specparam_declaration_instance12999();
    specparam_declaration13000 specparam_declaration_instance13000();
    specparam_declaration13001 specparam_declaration_instance13001();
    specparam_declaration13002 specparam_declaration_instance13002();
    specparam_declaration13003 specparam_declaration_instance13003();
    specparam_declaration13004 specparam_declaration_instance13004();
    specparam_declaration13005 specparam_declaration_instance13005();
    specparam_declaration13006 specparam_declaration_instance13006();
    specparam_declaration13007 specparam_declaration_instance13007();
    specparam_declaration13008 specparam_declaration_instance13008();
    specparam_declaration13009 specparam_declaration_instance13009();
    specparam_declaration13010 specparam_declaration_instance13010();
    specparam_declaration13011 specparam_declaration_instance13011();
    specparam_declaration13012 specparam_declaration_instance13012();
    specparam_declaration13013 specparam_declaration_instance13013();
    specparam_declaration13014 specparam_declaration_instance13014();
    specparam_declaration13015 specparam_declaration_instance13015();
    specparam_declaration13016 specparam_declaration_instance13016();
    specparam_declaration13017 specparam_declaration_instance13017();
    specparam_declaration13018 specparam_declaration_instance13018();
    specparam_declaration13019 specparam_declaration_instance13019();
    specparam_declaration13020 specparam_declaration_instance13020();
    specparam_declaration13021 specparam_declaration_instance13021();
    specparam_declaration13022 specparam_declaration_instance13022();
    specparam_declaration13023 specparam_declaration_instance13023();
    specparam_declaration13024 specparam_declaration_instance13024();
    specparam_declaration13025 specparam_declaration_instance13025();
    specparam_declaration13026 specparam_declaration_instance13026();
    specparam_declaration13027 specparam_declaration_instance13027();
    specparam_declaration13028 specparam_declaration_instance13028();
    specparam_declaration13029 specparam_declaration_instance13029();
    specparam_declaration13030 specparam_declaration_instance13030();
    specparam_declaration13031 specparam_declaration_instance13031();
    specparam_declaration13032 specparam_declaration_instance13032();
    specparam_declaration13033 specparam_declaration_instance13033();
    specparam_declaration13034 specparam_declaration_instance13034();
    specparam_declaration13035 specparam_declaration_instance13035();
    specparam_declaration13036 specparam_declaration_instance13036();
    specparam_declaration13037 specparam_declaration_instance13037();
    specparam_declaration13038 specparam_declaration_instance13038();
    specparam_declaration13039 specparam_declaration_instance13039();
    specparam_declaration13040 specparam_declaration_instance13040();
    specparam_declaration13041 specparam_declaration_instance13041();
    specparam_declaration13042 specparam_declaration_instance13042();
    specparam_declaration13043 specparam_declaration_instance13043();
    specparam_declaration13044 specparam_declaration_instance13044();
    specparam_declaration13045 specparam_declaration_instance13045();
    specparam_declaration13046 specparam_declaration_instance13046();
    specparam_declaration13047 specparam_declaration_instance13047();
    specparam_declaration13048 specparam_declaration_instance13048();
    specparam_declaration13049 specparam_declaration_instance13049();
    specparam_declaration13050 specparam_declaration_instance13050();
    specparam_declaration13051 specparam_declaration_instance13051();
    specparam_declaration13052 specparam_declaration_instance13052();
    specparam_declaration13053 specparam_declaration_instance13053();
    specparam_declaration13054 specparam_declaration_instance13054();
    specparam_declaration13055 specparam_declaration_instance13055();
    specparam_declaration13056 specparam_declaration_instance13056();
    specparam_declaration13057 specparam_declaration_instance13057();
    specparam_declaration13058 specparam_declaration_instance13058();
    specparam_declaration13059 specparam_declaration_instance13059();
    specparam_declaration13060 specparam_declaration_instance13060();
    specparam_declaration13061 specparam_declaration_instance13061();
    specparam_declaration13062 specparam_declaration_instance13062();
    specparam_declaration13063 specparam_declaration_instance13063();
    specparam_declaration13064 specparam_declaration_instance13064();
    specparam_declaration13065 specparam_declaration_instance13065();
    specparam_declaration13066 specparam_declaration_instance13066();
    specparam_declaration13067 specparam_declaration_instance13067();
    specparam_declaration13068 specparam_declaration_instance13068();
    specparam_declaration13069 specparam_declaration_instance13069();
    specparam_declaration13070 specparam_declaration_instance13070();
    specparam_declaration13071 specparam_declaration_instance13071();
    specparam_declaration13072 specparam_declaration_instance13072();
    specparam_declaration13073 specparam_declaration_instance13073();
    specparam_declaration13074 specparam_declaration_instance13074();
    specparam_declaration13075 specparam_declaration_instance13075();
    specparam_declaration13076 specparam_declaration_instance13076();
    specparam_declaration13077 specparam_declaration_instance13077();
    specparam_declaration13078 specparam_declaration_instance13078();
    specparam_declaration13079 specparam_declaration_instance13079();
    specparam_declaration13080 specparam_declaration_instance13080();
    specparam_declaration13081 specparam_declaration_instance13081();
    specparam_declaration13082 specparam_declaration_instance13082();
    specparam_declaration13083 specparam_declaration_instance13083();
    specparam_declaration13084 specparam_declaration_instance13084();
    specparam_declaration13085 specparam_declaration_instance13085();
    specparam_declaration13086 specparam_declaration_instance13086();
    specparam_declaration13087 specparam_declaration_instance13087();
    specparam_declaration13088 specparam_declaration_instance13088();
    specparam_declaration13089 specparam_declaration_instance13089();
    specparam_declaration13090 specparam_declaration_instance13090();
    specparam_declaration13091 specparam_declaration_instance13091();
    specparam_declaration13092 specparam_declaration_instance13092();
    specparam_declaration13093 specparam_declaration_instance13093();
    specparam_declaration13094 specparam_declaration_instance13094();
    specparam_declaration13095 specparam_declaration_instance13095();
    specparam_declaration13096 specparam_declaration_instance13096();
    specparam_declaration13097 specparam_declaration_instance13097();
    specparam_declaration13098 specparam_declaration_instance13098();
    specparam_declaration13099 specparam_declaration_instance13099();
    specparam_declaration13100 specparam_declaration_instance13100();
    specparam_declaration13101 specparam_declaration_instance13101();
    specparam_declaration13102 specparam_declaration_instance13102();
    specparam_declaration13103 specparam_declaration_instance13103();
    specparam_declaration13104 specparam_declaration_instance13104();
    specparam_declaration13105 specparam_declaration_instance13105();
    specparam_declaration13106 specparam_declaration_instance13106();
    specparam_declaration13107 specparam_declaration_instance13107();
    specparam_declaration13108 specparam_declaration_instance13108();
    specparam_declaration13109 specparam_declaration_instance13109();
    specparam_declaration13110 specparam_declaration_instance13110();
    specparam_declaration13111 specparam_declaration_instance13111();
    specparam_declaration13112 specparam_declaration_instance13112();
    specparam_declaration13113 specparam_declaration_instance13113();
    specparam_declaration13114 specparam_declaration_instance13114();
    specparam_declaration13115 specparam_declaration_instance13115();
    specparam_declaration13116 specparam_declaration_instance13116();
    specparam_declaration13117 specparam_declaration_instance13117();
    specparam_declaration13118 specparam_declaration_instance13118();
    specparam_declaration13119 specparam_declaration_instance13119();
    specparam_declaration13120 specparam_declaration_instance13120();
    specparam_declaration13121 specparam_declaration_instance13121();
    specparam_declaration13122 specparam_declaration_instance13122();
    specparam_declaration13123 specparam_declaration_instance13123();
    specparam_declaration13124 specparam_declaration_instance13124();
    specparam_declaration13125 specparam_declaration_instance13125();
    specparam_declaration13126 specparam_declaration_instance13126();
    specparam_declaration13127 specparam_declaration_instance13127();
    specparam_declaration13128 specparam_declaration_instance13128();
    specparam_declaration13129 specparam_declaration_instance13129();
    specparam_declaration13130 specparam_declaration_instance13130();
    specparam_declaration13131 specparam_declaration_instance13131();
    specparam_declaration13132 specparam_declaration_instance13132();
    specparam_declaration13133 specparam_declaration_instance13133();
    specparam_declaration13134 specparam_declaration_instance13134();
    specparam_declaration13135 specparam_declaration_instance13135();
    specparam_declaration13136 specparam_declaration_instance13136();
    specparam_declaration13137 specparam_declaration_instance13137();
    specparam_declaration13138 specparam_declaration_instance13138();
    specparam_declaration13139 specparam_declaration_instance13139();
    specparam_declaration13140 specparam_declaration_instance13140();
    specparam_declaration13141 specparam_declaration_instance13141();
    specparam_declaration13142 specparam_declaration_instance13142();
    specparam_declaration13143 specparam_declaration_instance13143();
    specparam_declaration13144 specparam_declaration_instance13144();
    specparam_declaration13145 specparam_declaration_instance13145();
    specparam_declaration13146 specparam_declaration_instance13146();
    specparam_declaration13147 specparam_declaration_instance13147();
    specparam_declaration13148 specparam_declaration_instance13148();
    specparam_declaration13149 specparam_declaration_instance13149();
    specparam_declaration13150 specparam_declaration_instance13150();
    specparam_declaration13151 specparam_declaration_instance13151();
    specparam_declaration13152 specparam_declaration_instance13152();
    specparam_declaration13153 specparam_declaration_instance13153();
    specparam_declaration13154 specparam_declaration_instance13154();
    specparam_declaration13155 specparam_declaration_instance13155();
    specparam_declaration13156 specparam_declaration_instance13156();
    specparam_declaration13157 specparam_declaration_instance13157();
    specparam_declaration13158 specparam_declaration_instance13158();
    specparam_declaration13159 specparam_declaration_instance13159();
    specparam_declaration13160 specparam_declaration_instance13160();
    specparam_declaration13161 specparam_declaration_instance13161();
    specparam_declaration13162 specparam_declaration_instance13162();
    specparam_declaration13163 specparam_declaration_instance13163();
    specparam_declaration13164 specparam_declaration_instance13164();
    specparam_declaration13165 specparam_declaration_instance13165();
    specparam_declaration13166 specparam_declaration_instance13166();
    specparam_declaration13167 specparam_declaration_instance13167();
    specparam_declaration13168 specparam_declaration_instance13168();
    specparam_declaration13169 specparam_declaration_instance13169();
    specparam_declaration13170 specparam_declaration_instance13170();
    specparam_declaration13171 specparam_declaration_instance13171();
    specparam_declaration13172 specparam_declaration_instance13172();
    specparam_declaration13173 specparam_declaration_instance13173();
    specparam_declaration13174 specparam_declaration_instance13174();
    specparam_declaration13175 specparam_declaration_instance13175();
    specparam_declaration13176 specparam_declaration_instance13176();
    specparam_declaration13177 specparam_declaration_instance13177();
    specparam_declaration13178 specparam_declaration_instance13178();
    specparam_declaration13179 specparam_declaration_instance13179();
    specparam_declaration13180 specparam_declaration_instance13180();
    specparam_declaration13181 specparam_declaration_instance13181();
    specparam_declaration13182 specparam_declaration_instance13182();
    specparam_declaration13183 specparam_declaration_instance13183();
    specparam_declaration13184 specparam_declaration_instance13184();
    specparam_declaration13185 specparam_declaration_instance13185();
    specparam_declaration13186 specparam_declaration_instance13186();
    specparam_declaration13187 specparam_declaration_instance13187();
    specparam_declaration13188 specparam_declaration_instance13188();
    specparam_declaration13189 specparam_declaration_instance13189();
    specparam_declaration13190 specparam_declaration_instance13190();
    specparam_declaration13191 specparam_declaration_instance13191();
    specparam_declaration13192 specparam_declaration_instance13192();
    specparam_declaration13193 specparam_declaration_instance13193();
    specparam_declaration13194 specparam_declaration_instance13194();
    specparam_declaration13195 specparam_declaration_instance13195();
    specparam_declaration13196 specparam_declaration_instance13196();
    specparam_declaration13197 specparam_declaration_instance13197();
    specparam_declaration13198 specparam_declaration_instance13198();
    specparam_declaration13199 specparam_declaration_instance13199();
    specparam_declaration13200 specparam_declaration_instance13200();
    specparam_declaration13201 specparam_declaration_instance13201();
    specparam_declaration13202 specparam_declaration_instance13202();
    specparam_declaration13203 specparam_declaration_instance13203();
    specparam_declaration13204 specparam_declaration_instance13204();
    specparam_declaration13205 specparam_declaration_instance13205();
    specparam_declaration13206 specparam_declaration_instance13206();
    specparam_declaration13207 specparam_declaration_instance13207();
    specparam_declaration13208 specparam_declaration_instance13208();
    specparam_declaration13209 specparam_declaration_instance13209();
    specparam_declaration13210 specparam_declaration_instance13210();
    specparam_declaration13211 specparam_declaration_instance13211();
    specparam_declaration13212 specparam_declaration_instance13212();
    specparam_declaration13213 specparam_declaration_instance13213();
    specparam_declaration13214 specparam_declaration_instance13214();
    specparam_declaration13215 specparam_declaration_instance13215();
    specparam_declaration13216 specparam_declaration_instance13216();
    specparam_declaration13217 specparam_declaration_instance13217();
    specparam_declaration13218 specparam_declaration_instance13218();
    specparam_declaration13219 specparam_declaration_instance13219();
    specparam_declaration13220 specparam_declaration_instance13220();
    specparam_declaration13221 specparam_declaration_instance13221();
    specparam_declaration13222 specparam_declaration_instance13222();
    specparam_declaration13223 specparam_declaration_instance13223();
    specparam_declaration13224 specparam_declaration_instance13224();
    specparam_declaration13225 specparam_declaration_instance13225();
    specparam_declaration13226 specparam_declaration_instance13226();
    specparam_declaration13227 specparam_declaration_instance13227();
    specparam_declaration13228 specparam_declaration_instance13228();
    specparam_declaration13229 specparam_declaration_instance13229();
    specparam_declaration13230 specparam_declaration_instance13230();
    specparam_declaration13231 specparam_declaration_instance13231();
    specparam_declaration13232 specparam_declaration_instance13232();
    specparam_declaration13233 specparam_declaration_instance13233();
    specparam_declaration13234 specparam_declaration_instance13234();
    specparam_declaration13235 specparam_declaration_instance13235();
    specparam_declaration13236 specparam_declaration_instance13236();
    specparam_declaration13237 specparam_declaration_instance13237();
    specparam_declaration13238 specparam_declaration_instance13238();
    specparam_declaration13239 specparam_declaration_instance13239();
    specparam_declaration13240 specparam_declaration_instance13240();
    specparam_declaration13241 specparam_declaration_instance13241();
    specparam_declaration13242 specparam_declaration_instance13242();
    specparam_declaration13243 specparam_declaration_instance13243();
    specparam_declaration13244 specparam_declaration_instance13244();
    specparam_declaration13245 specparam_declaration_instance13245();
    specparam_declaration13246 specparam_declaration_instance13246();
    specparam_declaration13247 specparam_declaration_instance13247();
    specparam_declaration13248 specparam_declaration_instance13248();
    specparam_declaration13249 specparam_declaration_instance13249();
    specparam_declaration13250 specparam_declaration_instance13250();
    specparam_declaration13251 specparam_declaration_instance13251();
    specparam_declaration13252 specparam_declaration_instance13252();
    specparam_declaration13253 specparam_declaration_instance13253();
    specparam_declaration13254 specparam_declaration_instance13254();
    specparam_declaration13255 specparam_declaration_instance13255();
    specparam_declaration13256 specparam_declaration_instance13256();
    specparam_declaration13257 specparam_declaration_instance13257();
    specparam_declaration13258 specparam_declaration_instance13258();
    specparam_declaration13259 specparam_declaration_instance13259();
    specparam_declaration13260 specparam_declaration_instance13260();
    specparam_declaration13261 specparam_declaration_instance13261();
    specparam_declaration13262 specparam_declaration_instance13262();
    specparam_declaration13263 specparam_declaration_instance13263();
    specparam_declaration13264 specparam_declaration_instance13264();
    specparam_declaration13265 specparam_declaration_instance13265();
    specparam_declaration13266 specparam_declaration_instance13266();
    specparam_declaration13267 specparam_declaration_instance13267();
    specparam_declaration13268 specparam_declaration_instance13268();
    specparam_declaration13269 specparam_declaration_instance13269();
    specparam_declaration13270 specparam_declaration_instance13270();
    specparam_declaration13271 specparam_declaration_instance13271();
    specparam_declaration13272 specparam_declaration_instance13272();
    specparam_declaration13273 specparam_declaration_instance13273();
    specparam_declaration13274 specparam_declaration_instance13274();
    specparam_declaration13275 specparam_declaration_instance13275();
    specparam_declaration13276 specparam_declaration_instance13276();
    specparam_declaration13277 specparam_declaration_instance13277();
    specparam_declaration13278 specparam_declaration_instance13278();
    specparam_declaration13279 specparam_declaration_instance13279();
    specparam_declaration13280 specparam_declaration_instance13280();
    specparam_declaration13281 specparam_declaration_instance13281();
    specparam_declaration13282 specparam_declaration_instance13282();
    specparam_declaration13283 specparam_declaration_instance13283();
    specparam_declaration13284 specparam_declaration_instance13284();
    specparam_declaration13285 specparam_declaration_instance13285();
    specparam_declaration13286 specparam_declaration_instance13286();
    specparam_declaration13287 specparam_declaration_instance13287();
    specparam_declaration13288 specparam_declaration_instance13288();
    specparam_declaration13289 specparam_declaration_instance13289();
    specparam_declaration13290 specparam_declaration_instance13290();
    specparam_declaration13291 specparam_declaration_instance13291();
    specparam_declaration13292 specparam_declaration_instance13292();
    specparam_declaration13293 specparam_declaration_instance13293();
    specparam_declaration13294 specparam_declaration_instance13294();
    specparam_declaration13295 specparam_declaration_instance13295();
    specparam_declaration13296 specparam_declaration_instance13296();
    specparam_declaration13297 specparam_declaration_instance13297();
    specparam_declaration13298 specparam_declaration_instance13298();
    specparam_declaration13299 specparam_declaration_instance13299();
    specparam_declaration13300 specparam_declaration_instance13300();
    specparam_declaration13301 specparam_declaration_instance13301();
    specparam_declaration13302 specparam_declaration_instance13302();
    specparam_declaration13303 specparam_declaration_instance13303();
    specparam_declaration13304 specparam_declaration_instance13304();
    specparam_declaration13305 specparam_declaration_instance13305();
    specparam_declaration13306 specparam_declaration_instance13306();
    specparam_declaration13307 specparam_declaration_instance13307();
    specparam_declaration13308 specparam_declaration_instance13308();
    specparam_declaration13309 specparam_declaration_instance13309();
    specparam_declaration13310 specparam_declaration_instance13310();
    specparam_declaration13311 specparam_declaration_instance13311();
    specparam_declaration13312 specparam_declaration_instance13312();
    specparam_declaration13313 specparam_declaration_instance13313();
    specparam_declaration13314 specparam_declaration_instance13314();
    specparam_declaration13315 specparam_declaration_instance13315();
    specparam_declaration13316 specparam_declaration_instance13316();
    specparam_declaration13317 specparam_declaration_instance13317();
    specparam_declaration13318 specparam_declaration_instance13318();
    specparam_declaration13319 specparam_declaration_instance13319();
    specparam_declaration13320 specparam_declaration_instance13320();
    specparam_declaration13321 specparam_declaration_instance13321();
    specparam_declaration13322 specparam_declaration_instance13322();
    specparam_declaration13323 specparam_declaration_instance13323();
    specparam_declaration13324 specparam_declaration_instance13324();
    specparam_declaration13325 specparam_declaration_instance13325();
    specparam_declaration13326 specparam_declaration_instance13326();
    specparam_declaration13327 specparam_declaration_instance13327();
    specparam_declaration13328 specparam_declaration_instance13328();
    specparam_declaration13329 specparam_declaration_instance13329();
    specparam_declaration13330 specparam_declaration_instance13330();
    specparam_declaration13331 specparam_declaration_instance13331();
    specparam_declaration13332 specparam_declaration_instance13332();
    specparam_declaration13333 specparam_declaration_instance13333();
    specparam_declaration13334 specparam_declaration_instance13334();
    specparam_declaration13335 specparam_declaration_instance13335();
    specparam_declaration13336 specparam_declaration_instance13336();
    specparam_declaration13337 specparam_declaration_instance13337();
    specparam_declaration13338 specparam_declaration_instance13338();
    specparam_declaration13339 specparam_declaration_instance13339();
    specparam_declaration13340 specparam_declaration_instance13340();
    specparam_declaration13341 specparam_declaration_instance13341();
    specparam_declaration13342 specparam_declaration_instance13342();
    specparam_declaration13343 specparam_declaration_instance13343();
    specparam_declaration13344 specparam_declaration_instance13344();
    specparam_declaration13345 specparam_declaration_instance13345();
    specparam_declaration13346 specparam_declaration_instance13346();
    specparam_declaration13347 specparam_declaration_instance13347();
    specparam_declaration13348 specparam_declaration_instance13348();
    specparam_declaration13349 specparam_declaration_instance13349();
    specparam_declaration13350 specparam_declaration_instance13350();
    specparam_declaration13351 specparam_declaration_instance13351();
    specparam_declaration13352 specparam_declaration_instance13352();
    specparam_declaration13353 specparam_declaration_instance13353();
    specparam_declaration13354 specparam_declaration_instance13354();
    specparam_declaration13355 specparam_declaration_instance13355();
    specparam_declaration13356 specparam_declaration_instance13356();
    specparam_declaration13357 specparam_declaration_instance13357();
    specparam_declaration13358 specparam_declaration_instance13358();
    specparam_declaration13359 specparam_declaration_instance13359();
    specparam_declaration13360 specparam_declaration_instance13360();
    specparam_declaration13361 specparam_declaration_instance13361();
    specparam_declaration13362 specparam_declaration_instance13362();
    specparam_declaration13363 specparam_declaration_instance13363();
    specparam_declaration13364 specparam_declaration_instance13364();
    specparam_declaration13365 specparam_declaration_instance13365();
    specparam_declaration13366 specparam_declaration_instance13366();
    specparam_declaration13367 specparam_declaration_instance13367();
    specparam_declaration13368 specparam_declaration_instance13368();
    specparam_declaration13369 specparam_declaration_instance13369();
    specparam_declaration13370 specparam_declaration_instance13370();
    specparam_declaration13371 specparam_declaration_instance13371();
    specparam_declaration13372 specparam_declaration_instance13372();
    specparam_declaration13373 specparam_declaration_instance13373();
    specparam_declaration13374 specparam_declaration_instance13374();
    specparam_declaration13375 specparam_declaration_instance13375();
    specparam_declaration13376 specparam_declaration_instance13376();
    specparam_declaration13377 specparam_declaration_instance13377();
    specparam_declaration13378 specparam_declaration_instance13378();
    specparam_declaration13379 specparam_declaration_instance13379();
    specparam_declaration13380 specparam_declaration_instance13380();
    specparam_declaration13381 specparam_declaration_instance13381();
    specparam_declaration13382 specparam_declaration_instance13382();
    specparam_declaration13383 specparam_declaration_instance13383();
    specparam_declaration13384 specparam_declaration_instance13384();
    specparam_declaration13385 specparam_declaration_instance13385();
    specparam_declaration13386 specparam_declaration_instance13386();
    specparam_declaration13387 specparam_declaration_instance13387();
    specparam_declaration13388 specparam_declaration_instance13388();
    specparam_declaration13389 specparam_declaration_instance13389();
    specparam_declaration13390 specparam_declaration_instance13390();
    specparam_declaration13391 specparam_declaration_instance13391();
    specparam_declaration13392 specparam_declaration_instance13392();
    specparam_declaration13393 specparam_declaration_instance13393();
    specparam_declaration13394 specparam_declaration_instance13394();
    specparam_declaration13395 specparam_declaration_instance13395();
    specparam_declaration13396 specparam_declaration_instance13396();
    specparam_declaration13397 specparam_declaration_instance13397();
    specparam_declaration13398 specparam_declaration_instance13398();
    specparam_declaration13399 specparam_declaration_instance13399();
    specparam_declaration13400 specparam_declaration_instance13400();
    specparam_declaration13401 specparam_declaration_instance13401();
    specparam_declaration13402 specparam_declaration_instance13402();
    specparam_declaration13403 specparam_declaration_instance13403();
    specparam_declaration13404 specparam_declaration_instance13404();
    specparam_declaration13405 specparam_declaration_instance13405();
    specparam_declaration13406 specparam_declaration_instance13406();
    specparam_declaration13407 specparam_declaration_instance13407();
    specparam_declaration13408 specparam_declaration_instance13408();
    specparam_declaration13409 specparam_declaration_instance13409();
    specparam_declaration13410 specparam_declaration_instance13410();
    specparam_declaration13411 specparam_declaration_instance13411();
    specparam_declaration13412 specparam_declaration_instance13412();
    specparam_declaration13413 specparam_declaration_instance13413();
    specparam_declaration13414 specparam_declaration_instance13414();
    specparam_declaration13415 specparam_declaration_instance13415();
    specparam_declaration13416 specparam_declaration_instance13416();
    specparam_declaration13417 specparam_declaration_instance13417();
    specparam_declaration13418 specparam_declaration_instance13418();
    specparam_declaration13419 specparam_declaration_instance13419();
    specparam_declaration13420 specparam_declaration_instance13420();
    specparam_declaration13421 specparam_declaration_instance13421();
    specparam_declaration13422 specparam_declaration_instance13422();
    specparam_declaration13423 specparam_declaration_instance13423();
    specparam_declaration13424 specparam_declaration_instance13424();
    specparam_declaration13425 specparam_declaration_instance13425();
    specparam_declaration13426 specparam_declaration_instance13426();
    specparam_declaration13427 specparam_declaration_instance13427();
    specparam_declaration13428 specparam_declaration_instance13428();
    specparam_declaration13429 specparam_declaration_instance13429();
    specparam_declaration13430 specparam_declaration_instance13430();
    specparam_declaration13431 specparam_declaration_instance13431();
    specparam_declaration13432 specparam_declaration_instance13432();
    specparam_declaration13433 specparam_declaration_instance13433();
    specparam_declaration13434 specparam_declaration_instance13434();
    specparam_declaration13435 specparam_declaration_instance13435();
    specparam_declaration13436 specparam_declaration_instance13436();
    specparam_declaration13437 specparam_declaration_instance13437();
    specparam_declaration13438 specparam_declaration_instance13438();
    specparam_declaration13439 specparam_declaration_instance13439();
    specparam_declaration13440 specparam_declaration_instance13440();
    specparam_declaration13441 specparam_declaration_instance13441();
    specparam_declaration13442 specparam_declaration_instance13442();
    specparam_declaration13443 specparam_declaration_instance13443();
    specparam_declaration13444 specparam_declaration_instance13444();
    specparam_declaration13445 specparam_declaration_instance13445();
    specparam_declaration13446 specparam_declaration_instance13446();
    specparam_declaration13447 specparam_declaration_instance13447();
    specparam_declaration13448 specparam_declaration_instance13448();
    specparam_declaration13449 specparam_declaration_instance13449();
    specparam_declaration13450 specparam_declaration_instance13450();
    specparam_declaration13451 specparam_declaration_instance13451();
    specparam_declaration13452 specparam_declaration_instance13452();
    specparam_declaration13453 specparam_declaration_instance13453();
    specparam_declaration13454 specparam_declaration_instance13454();
    specparam_declaration13455 specparam_declaration_instance13455();
    specparam_declaration13456 specparam_declaration_instance13456();
    specparam_declaration13457 specparam_declaration_instance13457();
    specparam_declaration13458 specparam_declaration_instance13458();
    specparam_declaration13459 specparam_declaration_instance13459();
    specparam_declaration13460 specparam_declaration_instance13460();
    specparam_declaration13461 specparam_declaration_instance13461();
    specparam_declaration13462 specparam_declaration_instance13462();
    specparam_declaration13463 specparam_declaration_instance13463();
    specparam_declaration13464 specparam_declaration_instance13464();
    specparam_declaration13465 specparam_declaration_instance13465();
    specparam_declaration13466 specparam_declaration_instance13466();
    specparam_declaration13467 specparam_declaration_instance13467();
    specparam_declaration13468 specparam_declaration_instance13468();
    specparam_declaration13469 specparam_declaration_instance13469();
    specparam_declaration13470 specparam_declaration_instance13470();
    specparam_declaration13471 specparam_declaration_instance13471();
    specparam_declaration13472 specparam_declaration_instance13472();
    specparam_declaration13473 specparam_declaration_instance13473();
    specparam_declaration13474 specparam_declaration_instance13474();
    specparam_declaration13475 specparam_declaration_instance13475();
    specparam_declaration13476 specparam_declaration_instance13476();
    specparam_declaration13477 specparam_declaration_instance13477();
    specparam_declaration13478 specparam_declaration_instance13478();
    specparam_declaration13479 specparam_declaration_instance13479();
    specparam_declaration13480 specparam_declaration_instance13480();
    specparam_declaration13481 specparam_declaration_instance13481();
    specparam_declaration13482 specparam_declaration_instance13482();
    specparam_declaration13483 specparam_declaration_instance13483();
    specparam_declaration13484 specparam_declaration_instance13484();
    specparam_declaration13485 specparam_declaration_instance13485();
    specparam_declaration13486 specparam_declaration_instance13486();
    specparam_declaration13487 specparam_declaration_instance13487();
    specparam_declaration13488 specparam_declaration_instance13488();
    specparam_declaration13489 specparam_declaration_instance13489();
    specparam_declaration13490 specparam_declaration_instance13490();
    specparam_declaration13491 specparam_declaration_instance13491();
    specparam_declaration13492 specparam_declaration_instance13492();
    specparam_declaration13493 specparam_declaration_instance13493();
    specparam_declaration13494 specparam_declaration_instance13494();
    specparam_declaration13495 specparam_declaration_instance13495();
    specparam_declaration13496 specparam_declaration_instance13496();
    specparam_declaration13497 specparam_declaration_instance13497();
    specparam_declaration13498 specparam_declaration_instance13498();
    specparam_declaration13499 specparam_declaration_instance13499();
    specparam_declaration13500 specparam_declaration_instance13500();
    specparam_declaration13501 specparam_declaration_instance13501();
    specparam_declaration13502 specparam_declaration_instance13502();
    specparam_declaration13503 specparam_declaration_instance13503();
    specparam_declaration13504 specparam_declaration_instance13504();
    specparam_declaration13505 specparam_declaration_instance13505();
    specparam_declaration13506 specparam_declaration_instance13506();
    specparam_declaration13507 specparam_declaration_instance13507();
    specparam_declaration13508 specparam_declaration_instance13508();
    specparam_declaration13509 specparam_declaration_instance13509();
    specparam_declaration13510 specparam_declaration_instance13510();
    specparam_declaration13511 specparam_declaration_instance13511();
    specparam_declaration13512 specparam_declaration_instance13512();
    specparam_declaration13513 specparam_declaration_instance13513();
    specparam_declaration13514 specparam_declaration_instance13514();
    specparam_declaration13515 specparam_declaration_instance13515();
    specparam_declaration13516 specparam_declaration_instance13516();
    specparam_declaration13517 specparam_declaration_instance13517();
    specparam_declaration13518 specparam_declaration_instance13518();
    specparam_declaration13519 specparam_declaration_instance13519();
    specparam_declaration13520 specparam_declaration_instance13520();
    specparam_declaration13521 specparam_declaration_instance13521();
    specparam_declaration13522 specparam_declaration_instance13522();
    specparam_declaration13523 specparam_declaration_instance13523();
    specparam_declaration13524 specparam_declaration_instance13524();
    specparam_declaration13525 specparam_declaration_instance13525();
    specparam_declaration13526 specparam_declaration_instance13526();
    specparam_declaration13527 specparam_declaration_instance13527();
    specparam_declaration13528 specparam_declaration_instance13528();
    specparam_declaration13529 specparam_declaration_instance13529();
    specparam_declaration13530 specparam_declaration_instance13530();
    specparam_declaration13531 specparam_declaration_instance13531();
    specparam_declaration13532 specparam_declaration_instance13532();
    specparam_declaration13533 specparam_declaration_instance13533();
    specparam_declaration13534 specparam_declaration_instance13534();
    specparam_declaration13535 specparam_declaration_instance13535();
    specparam_declaration13536 specparam_declaration_instance13536();
    specparam_declaration13537 specparam_declaration_instance13537();
    specparam_declaration13538 specparam_declaration_instance13538();
    specparam_declaration13539 specparam_declaration_instance13539();
    specparam_declaration13540 specparam_declaration_instance13540();
    specparam_declaration13541 specparam_declaration_instance13541();
    specparam_declaration13542 specparam_declaration_instance13542();
    specparam_declaration13543 specparam_declaration_instance13543();
    specparam_declaration13544 specparam_declaration_instance13544();
    specparam_declaration13545 specparam_declaration_instance13545();
    specparam_declaration13546 specparam_declaration_instance13546();
    specparam_declaration13547 specparam_declaration_instance13547();
    specparam_declaration13548 specparam_declaration_instance13548();
    specparam_declaration13549 specparam_declaration_instance13549();
    specparam_declaration13550 specparam_declaration_instance13550();
    specparam_declaration13551 specparam_declaration_instance13551();
    specparam_declaration13552 specparam_declaration_instance13552();
    specparam_declaration13553 specparam_declaration_instance13553();
    specparam_declaration13554 specparam_declaration_instance13554();
    specparam_declaration13555 specparam_declaration_instance13555();
    specparam_declaration13556 specparam_declaration_instance13556();
    specparam_declaration13557 specparam_declaration_instance13557();
    specparam_declaration13558 specparam_declaration_instance13558();
    specparam_declaration13559 specparam_declaration_instance13559();
    specparam_declaration13560 specparam_declaration_instance13560();
    specparam_declaration13561 specparam_declaration_instance13561();
    specparam_declaration13562 specparam_declaration_instance13562();
    specparam_declaration13563 specparam_declaration_instance13563();
    specparam_declaration13564 specparam_declaration_instance13564();
    specparam_declaration13565 specparam_declaration_instance13565();
    specparam_declaration13566 specparam_declaration_instance13566();
    specparam_declaration13567 specparam_declaration_instance13567();
    specparam_declaration13568 specparam_declaration_instance13568();
    specparam_declaration13569 specparam_declaration_instance13569();
    specparam_declaration13570 specparam_declaration_instance13570();
    specparam_declaration13571 specparam_declaration_instance13571();
    specparam_declaration13572 specparam_declaration_instance13572();
    specparam_declaration13573 specparam_declaration_instance13573();
    specparam_declaration13574 specparam_declaration_instance13574();
    specparam_declaration13575 specparam_declaration_instance13575();
    specparam_declaration13576 specparam_declaration_instance13576();
    specparam_declaration13577 specparam_declaration_instance13577();
    specparam_declaration13578 specparam_declaration_instance13578();
    specparam_declaration13579 specparam_declaration_instance13579();
    specparam_declaration13580 specparam_declaration_instance13580();
    specparam_declaration13581 specparam_declaration_instance13581();
    specparam_declaration13582 specparam_declaration_instance13582();
    specparam_declaration13583 specparam_declaration_instance13583();
    specparam_declaration13584 specparam_declaration_instance13584();
    specparam_declaration13585 specparam_declaration_instance13585();
    specparam_declaration13586 specparam_declaration_instance13586();
    specparam_declaration13587 specparam_declaration_instance13587();
    specparam_declaration13588 specparam_declaration_instance13588();
    specparam_declaration13589 specparam_declaration_instance13589();
    specparam_declaration13590 specparam_declaration_instance13590();
    specparam_declaration13591 specparam_declaration_instance13591();
    specparam_declaration13592 specparam_declaration_instance13592();
    specparam_declaration13593 specparam_declaration_instance13593();
    specparam_declaration13594 specparam_declaration_instance13594();
    specparam_declaration13595 specparam_declaration_instance13595();
    specparam_declaration13596 specparam_declaration_instance13596();
    specparam_declaration13597 specparam_declaration_instance13597();
    specparam_declaration13598 specparam_declaration_instance13598();
    specparam_declaration13599 specparam_declaration_instance13599();
    specparam_declaration13600 specparam_declaration_instance13600();
    specparam_declaration13601 specparam_declaration_instance13601();
    specparam_declaration13602 specparam_declaration_instance13602();
    specparam_declaration13603 specparam_declaration_instance13603();
    specparam_declaration13604 specparam_declaration_instance13604();
    specparam_declaration13605 specparam_declaration_instance13605();
    specparam_declaration13606 specparam_declaration_instance13606();
    specparam_declaration13607 specparam_declaration_instance13607();
    specparam_declaration13608 specparam_declaration_instance13608();
    specparam_declaration13609 specparam_declaration_instance13609();
    specparam_declaration13610 specparam_declaration_instance13610();
    specparam_declaration13611 specparam_declaration_instance13611();
    specparam_declaration13612 specparam_declaration_instance13612();
    specparam_declaration13613 specparam_declaration_instance13613();
    specparam_declaration13614 specparam_declaration_instance13614();
    specparam_declaration13615 specparam_declaration_instance13615();
    specparam_declaration13616 specparam_declaration_instance13616();
    specparam_declaration13617 specparam_declaration_instance13617();
    specparam_declaration13618 specparam_declaration_instance13618();
    specparam_declaration13619 specparam_declaration_instance13619();
    specparam_declaration13620 specparam_declaration_instance13620();
    specparam_declaration13621 specparam_declaration_instance13621();
    specparam_declaration13622 specparam_declaration_instance13622();
    specparam_declaration13623 specparam_declaration_instance13623();
    specparam_declaration13624 specparam_declaration_instance13624();
    specparam_declaration13625 specparam_declaration_instance13625();
    specparam_declaration13626 specparam_declaration_instance13626();
    specparam_declaration13627 specparam_declaration_instance13627();
    specparam_declaration13628 specparam_declaration_instance13628();
    specparam_declaration13629 specparam_declaration_instance13629();
    specparam_declaration13630 specparam_declaration_instance13630();
    specparam_declaration13631 specparam_declaration_instance13631();
    specparam_declaration13632 specparam_declaration_instance13632();
    specparam_declaration13633 specparam_declaration_instance13633();
    specparam_declaration13634 specparam_declaration_instance13634();
    specparam_declaration13635 specparam_declaration_instance13635();
    specparam_declaration13636 specparam_declaration_instance13636();
    specparam_declaration13637 specparam_declaration_instance13637();
    specparam_declaration13638 specparam_declaration_instance13638();
    specparam_declaration13639 specparam_declaration_instance13639();
    specparam_declaration13640 specparam_declaration_instance13640();
    specparam_declaration13641 specparam_declaration_instance13641();
    specparam_declaration13642 specparam_declaration_instance13642();
    specparam_declaration13643 specparam_declaration_instance13643();
    specparam_declaration13644 specparam_declaration_instance13644();
    specparam_declaration13645 specparam_declaration_instance13645();
    specparam_declaration13646 specparam_declaration_instance13646();
    specparam_declaration13647 specparam_declaration_instance13647();
    specparam_declaration13648 specparam_declaration_instance13648();
    specparam_declaration13649 specparam_declaration_instance13649();
    specparam_declaration13650 specparam_declaration_instance13650();
    specparam_declaration13651 specparam_declaration_instance13651();
    specparam_declaration13652 specparam_declaration_instance13652();
    specparam_declaration13653 specparam_declaration_instance13653();
    specparam_declaration13654 specparam_declaration_instance13654();
    specparam_declaration13655 specparam_declaration_instance13655();
    specparam_declaration13656 specparam_declaration_instance13656();
    specparam_declaration13657 specparam_declaration_instance13657();
    specparam_declaration13658 specparam_declaration_instance13658();
    specparam_declaration13659 specparam_declaration_instance13659();
    specparam_declaration13660 specparam_declaration_instance13660();
    specparam_declaration13661 specparam_declaration_instance13661();
    specparam_declaration13662 specparam_declaration_instance13662();
    specparam_declaration13663 specparam_declaration_instance13663();
    specparam_declaration13664 specparam_declaration_instance13664();
    specparam_declaration13665 specparam_declaration_instance13665();
    specparam_declaration13666 specparam_declaration_instance13666();
    specparam_declaration13667 specparam_declaration_instance13667();
    specparam_declaration13668 specparam_declaration_instance13668();
    specparam_declaration13669 specparam_declaration_instance13669();
    specparam_declaration13670 specparam_declaration_instance13670();
    specparam_declaration13671 specparam_declaration_instance13671();
    specparam_declaration13672 specparam_declaration_instance13672();
    specparam_declaration13673 specparam_declaration_instance13673();
    specparam_declaration13674 specparam_declaration_instance13674();
    specparam_declaration13675 specparam_declaration_instance13675();
    specparam_declaration13676 specparam_declaration_instance13676();
    specparam_declaration13677 specparam_declaration_instance13677();
    specparam_declaration13678 specparam_declaration_instance13678();
    specparam_declaration13679 specparam_declaration_instance13679();
    specparam_declaration13680 specparam_declaration_instance13680();
    specparam_declaration13681 specparam_declaration_instance13681();
    specparam_declaration13682 specparam_declaration_instance13682();
    specparam_declaration13683 specparam_declaration_instance13683();
    specparam_declaration13684 specparam_declaration_instance13684();
    specparam_declaration13685 specparam_declaration_instance13685();
    specparam_declaration13686 specparam_declaration_instance13686();
    specparam_declaration13687 specparam_declaration_instance13687();
    specparam_declaration13688 specparam_declaration_instance13688();
    specparam_declaration13689 specparam_declaration_instance13689();
    specparam_declaration13690 specparam_declaration_instance13690();
    specparam_declaration13691 specparam_declaration_instance13691();
    specparam_declaration13692 specparam_declaration_instance13692();
    specparam_declaration13693 specparam_declaration_instance13693();
    specparam_declaration13694 specparam_declaration_instance13694();
    specparam_declaration13695 specparam_declaration_instance13695();
    specparam_declaration13696 specparam_declaration_instance13696();
    specparam_declaration13697 specparam_declaration_instance13697();
    specparam_declaration13698 specparam_declaration_instance13698();
    specparam_declaration13699 specparam_declaration_instance13699();
    specparam_declaration13700 specparam_declaration_instance13700();
    specparam_declaration13701 specparam_declaration_instance13701();
    specparam_declaration13702 specparam_declaration_instance13702();
    specparam_declaration13703 specparam_declaration_instance13703();
    specparam_declaration13704 specparam_declaration_instance13704();
    specparam_declaration13705 specparam_declaration_instance13705();
    specparam_declaration13706 specparam_declaration_instance13706();
    specparam_declaration13707 specparam_declaration_instance13707();
    specparam_declaration13708 specparam_declaration_instance13708();
    specparam_declaration13709 specparam_declaration_instance13709();
    specparam_declaration13710 specparam_declaration_instance13710();
    specparam_declaration13711 specparam_declaration_instance13711();
    specparam_declaration13712 specparam_declaration_instance13712();
    specparam_declaration13713 specparam_declaration_instance13713();
    specparam_declaration13714 specparam_declaration_instance13714();
    specparam_declaration13715 specparam_declaration_instance13715();
    specparam_declaration13716 specparam_declaration_instance13716();
    specparam_declaration13717 specparam_declaration_instance13717();
    specparam_declaration13718 specparam_declaration_instance13718();
    specparam_declaration13719 specparam_declaration_instance13719();
    specparam_declaration13720 specparam_declaration_instance13720();
    specparam_declaration13721 specparam_declaration_instance13721();
    specparam_declaration13722 specparam_declaration_instance13722();
    specparam_declaration13723 specparam_declaration_instance13723();
    specparam_declaration13724 specparam_declaration_instance13724();
    specparam_declaration13725 specparam_declaration_instance13725();
    specparam_declaration13726 specparam_declaration_instance13726();
    specparam_declaration13727 specparam_declaration_instance13727();
    specparam_declaration13728 specparam_declaration_instance13728();
    specparam_declaration13729 specparam_declaration_instance13729();
    specparam_declaration13730 specparam_declaration_instance13730();
    specparam_declaration13731 specparam_declaration_instance13731();
    specparam_declaration13732 specparam_declaration_instance13732();
    specparam_declaration13733 specparam_declaration_instance13733();
    specparam_declaration13734 specparam_declaration_instance13734();
    specparam_declaration13735 specparam_declaration_instance13735();
    specparam_declaration13736 specparam_declaration_instance13736();
    specparam_declaration13737 specparam_declaration_instance13737();
    specparam_declaration13738 specparam_declaration_instance13738();
    specparam_declaration13739 specparam_declaration_instance13739();
    specparam_declaration13740 specparam_declaration_instance13740();
    specparam_declaration13741 specparam_declaration_instance13741();
    specparam_declaration13742 specparam_declaration_instance13742();
    specparam_declaration13743 specparam_declaration_instance13743();
    specparam_declaration13744 specparam_declaration_instance13744();
    specparam_declaration13745 specparam_declaration_instance13745();
    specparam_declaration13746 specparam_declaration_instance13746();
    specparam_declaration13747 specparam_declaration_instance13747();
    specparam_declaration13748 specparam_declaration_instance13748();
    specparam_declaration13749 specparam_declaration_instance13749();
    specparam_declaration13750 specparam_declaration_instance13750();
    specparam_declaration13751 specparam_declaration_instance13751();
    specparam_declaration13752 specparam_declaration_instance13752();
    specparam_declaration13753 specparam_declaration_instance13753();
    specparam_declaration13754 specparam_declaration_instance13754();
    specparam_declaration13755 specparam_declaration_instance13755();
    specparam_declaration13756 specparam_declaration_instance13756();
    specparam_declaration13757 specparam_declaration_instance13757();
    specparam_declaration13758 specparam_declaration_instance13758();
    specparam_declaration13759 specparam_declaration_instance13759();
    specparam_declaration13760 specparam_declaration_instance13760();
    specparam_declaration13761 specparam_declaration_instance13761();
    specparam_declaration13762 specparam_declaration_instance13762();
    specparam_declaration13763 specparam_declaration_instance13763();
    specparam_declaration13764 specparam_declaration_instance13764();
    specparam_declaration13765 specparam_declaration_instance13765();
    specparam_declaration13766 specparam_declaration_instance13766();
    specparam_declaration13767 specparam_declaration_instance13767();
    specparam_declaration13768 specparam_declaration_instance13768();
    specparam_declaration13769 specparam_declaration_instance13769();
    specparam_declaration13770 specparam_declaration_instance13770();
    specparam_declaration13771 specparam_declaration_instance13771();
    specparam_declaration13772 specparam_declaration_instance13772();
    specparam_declaration13773 specparam_declaration_instance13773();
    specparam_declaration13774 specparam_declaration_instance13774();
    specparam_declaration13775 specparam_declaration_instance13775();
    specparam_declaration13776 specparam_declaration_instance13776();
    specparam_declaration13777 specparam_declaration_instance13777();
    specparam_declaration13778 specparam_declaration_instance13778();
    specparam_declaration13779 specparam_declaration_instance13779();
    specparam_declaration13780 specparam_declaration_instance13780();
    specparam_declaration13781 specparam_declaration_instance13781();
    specparam_declaration13782 specparam_declaration_instance13782();
    specparam_declaration13783 specparam_declaration_instance13783();
    specparam_declaration13784 specparam_declaration_instance13784();
    specparam_declaration13785 specparam_declaration_instance13785();
    specparam_declaration13786 specparam_declaration_instance13786();
    specparam_declaration13787 specparam_declaration_instance13787();
    specparam_declaration13788 specparam_declaration_instance13788();
    specparam_declaration13789 specparam_declaration_instance13789();
    specparam_declaration13790 specparam_declaration_instance13790();
    specparam_declaration13791 specparam_declaration_instance13791();
    specparam_declaration13792 specparam_declaration_instance13792();
    specparam_declaration13793 specparam_declaration_instance13793();
    specparam_declaration13794 specparam_declaration_instance13794();
    specparam_declaration13795 specparam_declaration_instance13795();
    specparam_declaration13796 specparam_declaration_instance13796();
    specparam_declaration13797 specparam_declaration_instance13797();
    specparam_declaration13798 specparam_declaration_instance13798();
    specparam_declaration13799 specparam_declaration_instance13799();
    specparam_declaration13800 specparam_declaration_instance13800();
    specparam_declaration13801 specparam_declaration_instance13801();
    specparam_declaration13802 specparam_declaration_instance13802();
    specparam_declaration13803 specparam_declaration_instance13803();
    specparam_declaration13804 specparam_declaration_instance13804();
    specparam_declaration13805 specparam_declaration_instance13805();
    specparam_declaration13806 specparam_declaration_instance13806();
    specparam_declaration13807 specparam_declaration_instance13807();
    specparam_declaration13808 specparam_declaration_instance13808();
    specparam_declaration13809 specparam_declaration_instance13809();
    specparam_declaration13810 specparam_declaration_instance13810();
    specparam_declaration13811 specparam_declaration_instance13811();
    specparam_declaration13812 specparam_declaration_instance13812();
    specparam_declaration13813 specparam_declaration_instance13813();
    specparam_declaration13814 specparam_declaration_instance13814();
    specparam_declaration13815 specparam_declaration_instance13815();
    specparam_declaration13816 specparam_declaration_instance13816();
    specparam_declaration13817 specparam_declaration_instance13817();
    specparam_declaration13818 specparam_declaration_instance13818();
    specparam_declaration13819 specparam_declaration_instance13819();
    specparam_declaration13820 specparam_declaration_instance13820();
    specparam_declaration13821 specparam_declaration_instance13821();
    specparam_declaration13822 specparam_declaration_instance13822();
    specparam_declaration13823 specparam_declaration_instance13823();
    specparam_declaration13824 specparam_declaration_instance13824();
    specparam_declaration13825 specparam_declaration_instance13825();
    specparam_declaration13826 specparam_declaration_instance13826();
    specparam_declaration13827 specparam_declaration_instance13827();
    specparam_declaration13828 specparam_declaration_instance13828();
    specparam_declaration13829 specparam_declaration_instance13829();
    specparam_declaration13830 specparam_declaration_instance13830();
    specparam_declaration13831 specparam_declaration_instance13831();
    specparam_declaration13832 specparam_declaration_instance13832();
    specparam_declaration13833 specparam_declaration_instance13833();
    specparam_declaration13834 specparam_declaration_instance13834();
    specparam_declaration13835 specparam_declaration_instance13835();
    specparam_declaration13836 specparam_declaration_instance13836();
    specparam_declaration13837 specparam_declaration_instance13837();
    specparam_declaration13838 specparam_declaration_instance13838();
    specparam_declaration13839 specparam_declaration_instance13839();
    specparam_declaration13840 specparam_declaration_instance13840();
    specparam_declaration13841 specparam_declaration_instance13841();
    specparam_declaration13842 specparam_declaration_instance13842();
    specparam_declaration13843 specparam_declaration_instance13843();
    specparam_declaration13844 specparam_declaration_instance13844();
    specparam_declaration13845 specparam_declaration_instance13845();
    specparam_declaration13846 specparam_declaration_instance13846();
    specparam_declaration13847 specparam_declaration_instance13847();
    specparam_declaration13848 specparam_declaration_instance13848();
    specparam_declaration13849 specparam_declaration_instance13849();
    specparam_declaration13850 specparam_declaration_instance13850();
    specparam_declaration13851 specparam_declaration_instance13851();
    specparam_declaration13852 specparam_declaration_instance13852();
    specparam_declaration13853 specparam_declaration_instance13853();
    specparam_declaration13854 specparam_declaration_instance13854();
    specparam_declaration13855 specparam_declaration_instance13855();
    specparam_declaration13856 specparam_declaration_instance13856();
    specparam_declaration13857 specparam_declaration_instance13857();
    specparam_declaration13858 specparam_declaration_instance13858();
    specparam_declaration13859 specparam_declaration_instance13859();
    specparam_declaration13860 specparam_declaration_instance13860();
    specparam_declaration13861 specparam_declaration_instance13861();
    specparam_declaration13862 specparam_declaration_instance13862();
    specparam_declaration13863 specparam_declaration_instance13863();
    specparam_declaration13864 specparam_declaration_instance13864();
    specparam_declaration13865 specparam_declaration_instance13865();
    specparam_declaration13866 specparam_declaration_instance13866();
    specparam_declaration13867 specparam_declaration_instance13867();
    specparam_declaration13868 specparam_declaration_instance13868();
    specparam_declaration13869 specparam_declaration_instance13869();
    specparam_declaration13870 specparam_declaration_instance13870();
    specparam_declaration13871 specparam_declaration_instance13871();
    specparam_declaration13872 specparam_declaration_instance13872();
    specparam_declaration13873 specparam_declaration_instance13873();
    specparam_declaration13874 specparam_declaration_instance13874();
    specparam_declaration13875 specparam_declaration_instance13875();
    specparam_declaration13876 specparam_declaration_instance13876();
    specparam_declaration13877 specparam_declaration_instance13877();
    specparam_declaration13878 specparam_declaration_instance13878();
    specparam_declaration13879 specparam_declaration_instance13879();
    specparam_declaration13880 specparam_declaration_instance13880();
    specparam_declaration13881 specparam_declaration_instance13881();
    specparam_declaration13882 specparam_declaration_instance13882();
    specparam_declaration13883 specparam_declaration_instance13883();
    specparam_declaration13884 specparam_declaration_instance13884();
    specparam_declaration13885 specparam_declaration_instance13885();
    specparam_declaration13886 specparam_declaration_instance13886();
    specparam_declaration13887 specparam_declaration_instance13887();
    specparam_declaration13888 specparam_declaration_instance13888();
    specparam_declaration13889 specparam_declaration_instance13889();
    specparam_declaration13890 specparam_declaration_instance13890();
    specparam_declaration13891 specparam_declaration_instance13891();
    specparam_declaration13892 specparam_declaration_instance13892();
    specparam_declaration13893 specparam_declaration_instance13893();
    specparam_declaration13894 specparam_declaration_instance13894();
    specparam_declaration13895 specparam_declaration_instance13895();
    specparam_declaration13896 specparam_declaration_instance13896();
    specparam_declaration13897 specparam_declaration_instance13897();
    specparam_declaration13898 specparam_declaration_instance13898();
    specparam_declaration13899 specparam_declaration_instance13899();
    specparam_declaration13900 specparam_declaration_instance13900();
    specparam_declaration13901 specparam_declaration_instance13901();
    specparam_declaration13902 specparam_declaration_instance13902();
    specparam_declaration13903 specparam_declaration_instance13903();
    specparam_declaration13904 specparam_declaration_instance13904();
    specparam_declaration13905 specparam_declaration_instance13905();
    specparam_declaration13906 specparam_declaration_instance13906();
    specparam_declaration13907 specparam_declaration_instance13907();
    specparam_declaration13908 specparam_declaration_instance13908();
    specparam_declaration13909 specparam_declaration_instance13909();
    specparam_declaration13910 specparam_declaration_instance13910();
    specparam_declaration13911 specparam_declaration_instance13911();
    specparam_declaration13912 specparam_declaration_instance13912();
    specparam_declaration13913 specparam_declaration_instance13913();
    specparam_declaration13914 specparam_declaration_instance13914();
    specparam_declaration13915 specparam_declaration_instance13915();
    specparam_declaration13916 specparam_declaration_instance13916();
    specparam_declaration13917 specparam_declaration_instance13917();
    specparam_declaration13918 specparam_declaration_instance13918();
    specparam_declaration13919 specparam_declaration_instance13919();
    specparam_declaration13920 specparam_declaration_instance13920();
    specparam_declaration13921 specparam_declaration_instance13921();
    specparam_declaration13922 specparam_declaration_instance13922();
    specparam_declaration13923 specparam_declaration_instance13923();
    specparam_declaration13924 specparam_declaration_instance13924();
    specparam_declaration13925 specparam_declaration_instance13925();
    specparam_declaration13926 specparam_declaration_instance13926();
    specparam_declaration13927 specparam_declaration_instance13927();
    specparam_declaration13928 specparam_declaration_instance13928();
    specparam_declaration13929 specparam_declaration_instance13929();
    specparam_declaration13930 specparam_declaration_instance13930();
    specparam_declaration13931 specparam_declaration_instance13931();
    specparam_declaration13932 specparam_declaration_instance13932();
    specparam_declaration13933 specparam_declaration_instance13933();
    specparam_declaration13934 specparam_declaration_instance13934();
    specparam_declaration13935 specparam_declaration_instance13935();
    specparam_declaration13936 specparam_declaration_instance13936();
    specparam_declaration13937 specparam_declaration_instance13937();
    specparam_declaration13938 specparam_declaration_instance13938();
    specparam_declaration13939 specparam_declaration_instance13939();
    specparam_declaration13940 specparam_declaration_instance13940();
    specparam_declaration13941 specparam_declaration_instance13941();
    specparam_declaration13942 specparam_declaration_instance13942();
    specparam_declaration13943 specparam_declaration_instance13943();
    specparam_declaration13944 specparam_declaration_instance13944();
    specparam_declaration13945 specparam_declaration_instance13945();
    specparam_declaration13946 specparam_declaration_instance13946();
    specparam_declaration13947 specparam_declaration_instance13947();
    specparam_declaration13948 specparam_declaration_instance13948();
    specparam_declaration13949 specparam_declaration_instance13949();
    specparam_declaration13950 specparam_declaration_instance13950();
    specparam_declaration13951 specparam_declaration_instance13951();
    specparam_declaration13952 specparam_declaration_instance13952();
    specparam_declaration13953 specparam_declaration_instance13953();
    specparam_declaration13954 specparam_declaration_instance13954();
    specparam_declaration13955 specparam_declaration_instance13955();
    specparam_declaration13956 specparam_declaration_instance13956();
    specparam_declaration13957 specparam_declaration_instance13957();
    specparam_declaration13958 specparam_declaration_instance13958();
    specparam_declaration13959 specparam_declaration_instance13959();
    specparam_declaration13960 specparam_declaration_instance13960();
    specparam_declaration13961 specparam_declaration_instance13961();
    specparam_declaration13962 specparam_declaration_instance13962();
    specparam_declaration13963 specparam_declaration_instance13963();
    specparam_declaration13964 specparam_declaration_instance13964();
    specparam_declaration13965 specparam_declaration_instance13965();
    specparam_declaration13966 specparam_declaration_instance13966();
    specparam_declaration13967 specparam_declaration_instance13967();
    specparam_declaration13968 specparam_declaration_instance13968();
    specparam_declaration13969 specparam_declaration_instance13969();
    specparam_declaration13970 specparam_declaration_instance13970();
    specparam_declaration13971 specparam_declaration_instance13971();
    specparam_declaration13972 specparam_declaration_instance13972();
    specparam_declaration13973 specparam_declaration_instance13973();
    specparam_declaration13974 specparam_declaration_instance13974();
    specparam_declaration13975 specparam_declaration_instance13975();
    specparam_declaration13976 specparam_declaration_instance13976();
    specparam_declaration13977 specparam_declaration_instance13977();
    specparam_declaration13978 specparam_declaration_instance13978();
    specparam_declaration13979 specparam_declaration_instance13979();
    specparam_declaration13980 specparam_declaration_instance13980();
    specparam_declaration13981 specparam_declaration_instance13981();
    specparam_declaration13982 specparam_declaration_instance13982();
    specparam_declaration13983 specparam_declaration_instance13983();
    specparam_declaration13984 specparam_declaration_instance13984();
    specparam_declaration13985 specparam_declaration_instance13985();
    specparam_declaration13986 specparam_declaration_instance13986();
    specparam_declaration13987 specparam_declaration_instance13987();
    specparam_declaration13988 specparam_declaration_instance13988();
    specparam_declaration13989 specparam_declaration_instance13989();
    specparam_declaration13990 specparam_declaration_instance13990();
    specparam_declaration13991 specparam_declaration_instance13991();
    specparam_declaration13992 specparam_declaration_instance13992();
    specparam_declaration13993 specparam_declaration_instance13993();
    specparam_declaration13994 specparam_declaration_instance13994();
    specparam_declaration13995 specparam_declaration_instance13995();
    specparam_declaration13996 specparam_declaration_instance13996();
    specparam_declaration13997 specparam_declaration_instance13997();
    specparam_declaration13998 specparam_declaration_instance13998();
    specparam_declaration13999 specparam_declaration_instance13999();
    specparam_declaration14000 specparam_declaration_instance14000();
    specparam_declaration14001 specparam_declaration_instance14001();
    specparam_declaration14002 specparam_declaration_instance14002();
    specparam_declaration14003 specparam_declaration_instance14003();
    specparam_declaration14004 specparam_declaration_instance14004();
    specparam_declaration14005 specparam_declaration_instance14005();
    specparam_declaration14006 specparam_declaration_instance14006();
    specparam_declaration14007 specparam_declaration_instance14007();
    specparam_declaration14008 specparam_declaration_instance14008();
    specparam_declaration14009 specparam_declaration_instance14009();
    specparam_declaration14010 specparam_declaration_instance14010();
    specparam_declaration14011 specparam_declaration_instance14011();
    specparam_declaration14012 specparam_declaration_instance14012();
    specparam_declaration14013 specparam_declaration_instance14013();
    specparam_declaration14014 specparam_declaration_instance14014();
    specparam_declaration14015 specparam_declaration_instance14015();
    specparam_declaration14016 specparam_declaration_instance14016();
    specparam_declaration14017 specparam_declaration_instance14017();
    specparam_declaration14018 specparam_declaration_instance14018();
    specparam_declaration14019 specparam_declaration_instance14019();
    specparam_declaration14020 specparam_declaration_instance14020();
    specparam_declaration14021 specparam_declaration_instance14021();
    specparam_declaration14022 specparam_declaration_instance14022();
    specparam_declaration14023 specparam_declaration_instance14023();
    specparam_declaration14024 specparam_declaration_instance14024();
    specparam_declaration14025 specparam_declaration_instance14025();
    specparam_declaration14026 specparam_declaration_instance14026();
    specparam_declaration14027 specparam_declaration_instance14027();
    specparam_declaration14028 specparam_declaration_instance14028();
    specparam_declaration14029 specparam_declaration_instance14029();
    specparam_declaration14030 specparam_declaration_instance14030();
    specparam_declaration14031 specparam_declaration_instance14031();
    specparam_declaration14032 specparam_declaration_instance14032();
    specparam_declaration14033 specparam_declaration_instance14033();
    specparam_declaration14034 specparam_declaration_instance14034();
    specparam_declaration14035 specparam_declaration_instance14035();
    specparam_declaration14036 specparam_declaration_instance14036();
    specparam_declaration14037 specparam_declaration_instance14037();
    specparam_declaration14038 specparam_declaration_instance14038();
    specparam_declaration14039 specparam_declaration_instance14039();
    specparam_declaration14040 specparam_declaration_instance14040();
    specparam_declaration14041 specparam_declaration_instance14041();
    specparam_declaration14042 specparam_declaration_instance14042();
    specparam_declaration14043 specparam_declaration_instance14043();
    specparam_declaration14044 specparam_declaration_instance14044();
    specparam_declaration14045 specparam_declaration_instance14045();
    specparam_declaration14046 specparam_declaration_instance14046();
    specparam_declaration14047 specparam_declaration_instance14047();
    specparam_declaration14048 specparam_declaration_instance14048();
    specparam_declaration14049 specparam_declaration_instance14049();
    specparam_declaration14050 specparam_declaration_instance14050();
    specparam_declaration14051 specparam_declaration_instance14051();
    specparam_declaration14052 specparam_declaration_instance14052();
    specparam_declaration14053 specparam_declaration_instance14053();
    specparam_declaration14054 specparam_declaration_instance14054();
    specparam_declaration14055 specparam_declaration_instance14055();
    specparam_declaration14056 specparam_declaration_instance14056();
    specparam_declaration14057 specparam_declaration_instance14057();
    specparam_declaration14058 specparam_declaration_instance14058();
    specparam_declaration14059 specparam_declaration_instance14059();
    specparam_declaration14060 specparam_declaration_instance14060();
    specparam_declaration14061 specparam_declaration_instance14061();
    specparam_declaration14062 specparam_declaration_instance14062();
    specparam_declaration14063 specparam_declaration_instance14063();
    specparam_declaration14064 specparam_declaration_instance14064();
    specparam_declaration14065 specparam_declaration_instance14065();
    specparam_declaration14066 specparam_declaration_instance14066();
    specparam_declaration14067 specparam_declaration_instance14067();
    specparam_declaration14068 specparam_declaration_instance14068();
    specparam_declaration14069 specparam_declaration_instance14069();
    specparam_declaration14070 specparam_declaration_instance14070();
    specparam_declaration14071 specparam_declaration_instance14071();
    specparam_declaration14072 specparam_declaration_instance14072();
    specparam_declaration14073 specparam_declaration_instance14073();
    specparam_declaration14074 specparam_declaration_instance14074();
    specparam_declaration14075 specparam_declaration_instance14075();
    specparam_declaration14076 specparam_declaration_instance14076();
    specparam_declaration14077 specparam_declaration_instance14077();
    specparam_declaration14078 specparam_declaration_instance14078();
    specparam_declaration14079 specparam_declaration_instance14079();
    specparam_declaration14080 specparam_declaration_instance14080();
    specparam_declaration14081 specparam_declaration_instance14081();
    specparam_declaration14082 specparam_declaration_instance14082();
    specparam_declaration14083 specparam_declaration_instance14083();
    specparam_declaration14084 specparam_declaration_instance14084();
    specparam_declaration14085 specparam_declaration_instance14085();
    specparam_declaration14086 specparam_declaration_instance14086();
    specparam_declaration14087 specparam_declaration_instance14087();
    specparam_declaration14088 specparam_declaration_instance14088();
    specparam_declaration14089 specparam_declaration_instance14089();
    specparam_declaration14090 specparam_declaration_instance14090();
    specparam_declaration14091 specparam_declaration_instance14091();
    specparam_declaration14092 specparam_declaration_instance14092();
    specparam_declaration14093 specparam_declaration_instance14093();
    specparam_declaration14094 specparam_declaration_instance14094();
    specparam_declaration14095 specparam_declaration_instance14095();
    specparam_declaration14096 specparam_declaration_instance14096();
    specparam_declaration14097 specparam_declaration_instance14097();
    specparam_declaration14098 specparam_declaration_instance14098();
    specparam_declaration14099 specparam_declaration_instance14099();
    specparam_declaration14100 specparam_declaration_instance14100();
    specparam_declaration14101 specparam_declaration_instance14101();
    specparam_declaration14102 specparam_declaration_instance14102();
    specparam_declaration14103 specparam_declaration_instance14103();
    specparam_declaration14104 specparam_declaration_instance14104();
    specparam_declaration14105 specparam_declaration_instance14105();
    specparam_declaration14106 specparam_declaration_instance14106();
    specparam_declaration14107 specparam_declaration_instance14107();
    specparam_declaration14108 specparam_declaration_instance14108();
    specparam_declaration14109 specparam_declaration_instance14109();
    specparam_declaration14110 specparam_declaration_instance14110();
    specparam_declaration14111 specparam_declaration_instance14111();
    specparam_declaration14112 specparam_declaration_instance14112();
    specparam_declaration14113 specparam_declaration_instance14113();
    specparam_declaration14114 specparam_declaration_instance14114();
    specparam_declaration14115 specparam_declaration_instance14115();
    specparam_declaration14116 specparam_declaration_instance14116();
    specparam_declaration14117 specparam_declaration_instance14117();
    specparam_declaration14118 specparam_declaration_instance14118();
    specparam_declaration14119 specparam_declaration_instance14119();
    specparam_declaration14120 specparam_declaration_instance14120();
    specparam_declaration14121 specparam_declaration_instance14121();
    specparam_declaration14122 specparam_declaration_instance14122();
    specparam_declaration14123 specparam_declaration_instance14123();
    specparam_declaration14124 specparam_declaration_instance14124();
    specparam_declaration14125 specparam_declaration_instance14125();
    specparam_declaration14126 specparam_declaration_instance14126();
    specparam_declaration14127 specparam_declaration_instance14127();
    specparam_declaration14128 specparam_declaration_instance14128();
    specparam_declaration14129 specparam_declaration_instance14129();
    specparam_declaration14130 specparam_declaration_instance14130();
    specparam_declaration14131 specparam_declaration_instance14131();
    specparam_declaration14132 specparam_declaration_instance14132();
    specparam_declaration14133 specparam_declaration_instance14133();
    specparam_declaration14134 specparam_declaration_instance14134();
    specparam_declaration14135 specparam_declaration_instance14135();
    specparam_declaration14136 specparam_declaration_instance14136();
    specparam_declaration14137 specparam_declaration_instance14137();
    specparam_declaration14138 specparam_declaration_instance14138();
    specparam_declaration14139 specparam_declaration_instance14139();
    specparam_declaration14140 specparam_declaration_instance14140();
    specparam_declaration14141 specparam_declaration_instance14141();
    specparam_declaration14142 specparam_declaration_instance14142();
    specparam_declaration14143 specparam_declaration_instance14143();
    specparam_declaration14144 specparam_declaration_instance14144();
    specparam_declaration14145 specparam_declaration_instance14145();
    specparam_declaration14146 specparam_declaration_instance14146();
    specparam_declaration14147 specparam_declaration_instance14147();
    specparam_declaration14148 specparam_declaration_instance14148();
    specparam_declaration14149 specparam_declaration_instance14149();
    specparam_declaration14150 specparam_declaration_instance14150();
    specparam_declaration14151 specparam_declaration_instance14151();
    specparam_declaration14152 specparam_declaration_instance14152();
    specparam_declaration14153 specparam_declaration_instance14153();
    specparam_declaration14154 specparam_declaration_instance14154();
    specparam_declaration14155 specparam_declaration_instance14155();
    specparam_declaration14156 specparam_declaration_instance14156();
    specparam_declaration14157 specparam_declaration_instance14157();
    specparam_declaration14158 specparam_declaration_instance14158();
    specparam_declaration14159 specparam_declaration_instance14159();
    specparam_declaration14160 specparam_declaration_instance14160();
    specparam_declaration14161 specparam_declaration_instance14161();
    specparam_declaration14162 specparam_declaration_instance14162();
    specparam_declaration14163 specparam_declaration_instance14163();
    specparam_declaration14164 specparam_declaration_instance14164();
    specparam_declaration14165 specparam_declaration_instance14165();
    specparam_declaration14166 specparam_declaration_instance14166();
    specparam_declaration14167 specparam_declaration_instance14167();
    specparam_declaration14168 specparam_declaration_instance14168();
    specparam_declaration14169 specparam_declaration_instance14169();
    specparam_declaration14170 specparam_declaration_instance14170();
    specparam_declaration14171 specparam_declaration_instance14171();
    specparam_declaration14172 specparam_declaration_instance14172();
    specparam_declaration14173 specparam_declaration_instance14173();
    specparam_declaration14174 specparam_declaration_instance14174();
    specparam_declaration14175 specparam_declaration_instance14175();
    specparam_declaration14176 specparam_declaration_instance14176();
    specparam_declaration14177 specparam_declaration_instance14177();
    specparam_declaration14178 specparam_declaration_instance14178();
    specparam_declaration14179 specparam_declaration_instance14179();
    specparam_declaration14180 specparam_declaration_instance14180();
    specparam_declaration14181 specparam_declaration_instance14181();
    specparam_declaration14182 specparam_declaration_instance14182();
    specparam_declaration14183 specparam_declaration_instance14183();
    specparam_declaration14184 specparam_declaration_instance14184();
    specparam_declaration14185 specparam_declaration_instance14185();
    specparam_declaration14186 specparam_declaration_instance14186();
    specparam_declaration14187 specparam_declaration_instance14187();
    specparam_declaration14188 specparam_declaration_instance14188();
    specparam_declaration14189 specparam_declaration_instance14189();
    specparam_declaration14190 specparam_declaration_instance14190();
    specparam_declaration14191 specparam_declaration_instance14191();
    specparam_declaration14192 specparam_declaration_instance14192();
    specparam_declaration14193 specparam_declaration_instance14193();
    specparam_declaration14194 specparam_declaration_instance14194();
    specparam_declaration14195 specparam_declaration_instance14195();
    specparam_declaration14196 specparam_declaration_instance14196();
    specparam_declaration14197 specparam_declaration_instance14197();
    specparam_declaration14198 specparam_declaration_instance14198();
    specparam_declaration14199 specparam_declaration_instance14199();
    specparam_declaration14200 specparam_declaration_instance14200();
    specparam_declaration14201 specparam_declaration_instance14201();
    specparam_declaration14202 specparam_declaration_instance14202();
    specparam_declaration14203 specparam_declaration_instance14203();
    specparam_declaration14204 specparam_declaration_instance14204();
    specparam_declaration14205 specparam_declaration_instance14205();
    specparam_declaration14206 specparam_declaration_instance14206();
    specparam_declaration14207 specparam_declaration_instance14207();
    specparam_declaration14208 specparam_declaration_instance14208();
    specparam_declaration14209 specparam_declaration_instance14209();
    specparam_declaration14210 specparam_declaration_instance14210();
    specparam_declaration14211 specparam_declaration_instance14211();
    specparam_declaration14212 specparam_declaration_instance14212();
    specparam_declaration14213 specparam_declaration_instance14213();
    specparam_declaration14214 specparam_declaration_instance14214();
    specparam_declaration14215 specparam_declaration_instance14215();
    specparam_declaration14216 specparam_declaration_instance14216();
    specparam_declaration14217 specparam_declaration_instance14217();
    specparam_declaration14218 specparam_declaration_instance14218();
    specparam_declaration14219 specparam_declaration_instance14219();
    specparam_declaration14220 specparam_declaration_instance14220();
    specparam_declaration14221 specparam_declaration_instance14221();
    specparam_declaration14222 specparam_declaration_instance14222();
    specparam_declaration14223 specparam_declaration_instance14223();
    specparam_declaration14224 specparam_declaration_instance14224();
    specparam_declaration14225 specparam_declaration_instance14225();
    specparam_declaration14226 specparam_declaration_instance14226();
    specparam_declaration14227 specparam_declaration_instance14227();
    specparam_declaration14228 specparam_declaration_instance14228();
    specparam_declaration14229 specparam_declaration_instance14229();
    specparam_declaration14230 specparam_declaration_instance14230();
    specparam_declaration14231 specparam_declaration_instance14231();
    specparam_declaration14232 specparam_declaration_instance14232();
    specparam_declaration14233 specparam_declaration_instance14233();
    specparam_declaration14234 specparam_declaration_instance14234();
    specparam_declaration14235 specparam_declaration_instance14235();
    specparam_declaration14236 specparam_declaration_instance14236();
    specparam_declaration14237 specparam_declaration_instance14237();
    specparam_declaration14238 specparam_declaration_instance14238();
    specparam_declaration14239 specparam_declaration_instance14239();
    specparam_declaration14240 specparam_declaration_instance14240();
    specparam_declaration14241 specparam_declaration_instance14241();
    specparam_declaration14242 specparam_declaration_instance14242();
    specparam_declaration14243 specparam_declaration_instance14243();
    specparam_declaration14244 specparam_declaration_instance14244();
    specparam_declaration14245 specparam_declaration_instance14245();
    specparam_declaration14246 specparam_declaration_instance14246();
    specparam_declaration14247 specparam_declaration_instance14247();
    specparam_declaration14248 specparam_declaration_instance14248();
    specparam_declaration14249 specparam_declaration_instance14249();
    specparam_declaration14250 specparam_declaration_instance14250();
    specparam_declaration14251 specparam_declaration_instance14251();
    specparam_declaration14252 specparam_declaration_instance14252();
    specparam_declaration14253 specparam_declaration_instance14253();
    specparam_declaration14254 specparam_declaration_instance14254();
    specparam_declaration14255 specparam_declaration_instance14255();
    specparam_declaration14256 specparam_declaration_instance14256();
    specparam_declaration14257 specparam_declaration_instance14257();
    specparam_declaration14258 specparam_declaration_instance14258();
    specparam_declaration14259 specparam_declaration_instance14259();
    specparam_declaration14260 specparam_declaration_instance14260();
    specparam_declaration14261 specparam_declaration_instance14261();
    specparam_declaration14262 specparam_declaration_instance14262();
    specparam_declaration14263 specparam_declaration_instance14263();
    specparam_declaration14264 specparam_declaration_instance14264();
    specparam_declaration14265 specparam_declaration_instance14265();
    specparam_declaration14266 specparam_declaration_instance14266();
    specparam_declaration14267 specparam_declaration_instance14267();
    specparam_declaration14268 specparam_declaration_instance14268();
    specparam_declaration14269 specparam_declaration_instance14269();
    specparam_declaration14270 specparam_declaration_instance14270();
    specparam_declaration14271 specparam_declaration_instance14271();
    specparam_declaration14272 specparam_declaration_instance14272();
    specparam_declaration14273 specparam_declaration_instance14273();
    specparam_declaration14274 specparam_declaration_instance14274();
    specparam_declaration14275 specparam_declaration_instance14275();
    specparam_declaration14276 specparam_declaration_instance14276();
    specparam_declaration14277 specparam_declaration_instance14277();
    specparam_declaration14278 specparam_declaration_instance14278();
    specparam_declaration14279 specparam_declaration_instance14279();
    specparam_declaration14280 specparam_declaration_instance14280();
    specparam_declaration14281 specparam_declaration_instance14281();
    specparam_declaration14282 specparam_declaration_instance14282();
    specparam_declaration14283 specparam_declaration_instance14283();
    specparam_declaration14284 specparam_declaration_instance14284();
    specparam_declaration14285 specparam_declaration_instance14285();
    specparam_declaration14286 specparam_declaration_instance14286();
    specparam_declaration14287 specparam_declaration_instance14287();
    specparam_declaration14288 specparam_declaration_instance14288();
    specparam_declaration14289 specparam_declaration_instance14289();
    specparam_declaration14290 specparam_declaration_instance14290();
    specparam_declaration14291 specparam_declaration_instance14291();
    specparam_declaration14292 specparam_declaration_instance14292();
    specparam_declaration14293 specparam_declaration_instance14293();
    specparam_declaration14294 specparam_declaration_instance14294();
    specparam_declaration14295 specparam_declaration_instance14295();
    specparam_declaration14296 specparam_declaration_instance14296();
    specparam_declaration14297 specparam_declaration_instance14297();
    specparam_declaration14298 specparam_declaration_instance14298();
    specparam_declaration14299 specparam_declaration_instance14299();
    specparam_declaration14300 specparam_declaration_instance14300();
    specparam_declaration14301 specparam_declaration_instance14301();
    specparam_declaration14302 specparam_declaration_instance14302();
    specparam_declaration14303 specparam_declaration_instance14303();
    specparam_declaration14304 specparam_declaration_instance14304();
    specparam_declaration14305 specparam_declaration_instance14305();
    specparam_declaration14306 specparam_declaration_instance14306();
    specparam_declaration14307 specparam_declaration_instance14307();
    specparam_declaration14308 specparam_declaration_instance14308();
    specparam_declaration14309 specparam_declaration_instance14309();
    specparam_declaration14310 specparam_declaration_instance14310();
    specparam_declaration14311 specparam_declaration_instance14311();
    specparam_declaration14312 specparam_declaration_instance14312();
    specparam_declaration14313 specparam_declaration_instance14313();
    specparam_declaration14314 specparam_declaration_instance14314();
    specparam_declaration14315 specparam_declaration_instance14315();
    specparam_declaration14316 specparam_declaration_instance14316();
    specparam_declaration14317 specparam_declaration_instance14317();
    specparam_declaration14318 specparam_declaration_instance14318();
    specparam_declaration14319 specparam_declaration_instance14319();
    specparam_declaration14320 specparam_declaration_instance14320();
    specparam_declaration14321 specparam_declaration_instance14321();
    specparam_declaration14322 specparam_declaration_instance14322();
    specparam_declaration14323 specparam_declaration_instance14323();
    specparam_declaration14324 specparam_declaration_instance14324();
    specparam_declaration14325 specparam_declaration_instance14325();
    specparam_declaration14326 specparam_declaration_instance14326();
    specparam_declaration14327 specparam_declaration_instance14327();
    specparam_declaration14328 specparam_declaration_instance14328();
    specparam_declaration14329 specparam_declaration_instance14329();
    specparam_declaration14330 specparam_declaration_instance14330();
    specparam_declaration14331 specparam_declaration_instance14331();
    specparam_declaration14332 specparam_declaration_instance14332();
    specparam_declaration14333 specparam_declaration_instance14333();
    specparam_declaration14334 specparam_declaration_instance14334();
    specparam_declaration14335 specparam_declaration_instance14335();
    specparam_declaration14336 specparam_declaration_instance14336();
    specparam_declaration14337 specparam_declaration_instance14337();
    specparam_declaration14338 specparam_declaration_instance14338();
    specparam_declaration14339 specparam_declaration_instance14339();
    specparam_declaration14340 specparam_declaration_instance14340();
    specparam_declaration14341 specparam_declaration_instance14341();
    specparam_declaration14342 specparam_declaration_instance14342();
    specparam_declaration14343 specparam_declaration_instance14343();
    specparam_declaration14344 specparam_declaration_instance14344();
    specparam_declaration14345 specparam_declaration_instance14345();
    specparam_declaration14346 specparam_declaration_instance14346();
    specparam_declaration14347 specparam_declaration_instance14347();
    specparam_declaration14348 specparam_declaration_instance14348();
    specparam_declaration14349 specparam_declaration_instance14349();
    specparam_declaration14350 specparam_declaration_instance14350();
    specparam_declaration14351 specparam_declaration_instance14351();
    specparam_declaration14352 specparam_declaration_instance14352();
    specparam_declaration14353 specparam_declaration_instance14353();
    specparam_declaration14354 specparam_declaration_instance14354();
    specparam_declaration14355 specparam_declaration_instance14355();
    specparam_declaration14356 specparam_declaration_instance14356();
    specparam_declaration14357 specparam_declaration_instance14357();
    specparam_declaration14358 specparam_declaration_instance14358();
    specparam_declaration14359 specparam_declaration_instance14359();
    specparam_declaration14360 specparam_declaration_instance14360();
    specparam_declaration14361 specparam_declaration_instance14361();
    specparam_declaration14362 specparam_declaration_instance14362();
    specparam_declaration14363 specparam_declaration_instance14363();
    specparam_declaration14364 specparam_declaration_instance14364();
    specparam_declaration14365 specparam_declaration_instance14365();
    specparam_declaration14366 specparam_declaration_instance14366();
    specparam_declaration14367 specparam_declaration_instance14367();
    specparam_declaration14368 specparam_declaration_instance14368();
    specparam_declaration14369 specparam_declaration_instance14369();
    specparam_declaration14370 specparam_declaration_instance14370();
    specparam_declaration14371 specparam_declaration_instance14371();
    specparam_declaration14372 specparam_declaration_instance14372();
    specparam_declaration14373 specparam_declaration_instance14373();
    specparam_declaration14374 specparam_declaration_instance14374();
    specparam_declaration14375 specparam_declaration_instance14375();
    specparam_declaration14376 specparam_declaration_instance14376();
    specparam_declaration14377 specparam_declaration_instance14377();
    specparam_declaration14378 specparam_declaration_instance14378();
    specparam_declaration14379 specparam_declaration_instance14379();
    specparam_declaration14380 specparam_declaration_instance14380();
    specparam_declaration14381 specparam_declaration_instance14381();
    specparam_declaration14382 specparam_declaration_instance14382();
    specparam_declaration14383 specparam_declaration_instance14383();
    specparam_declaration14384 specparam_declaration_instance14384();
    specparam_declaration14385 specparam_declaration_instance14385();
    specparam_declaration14386 specparam_declaration_instance14386();
    specparam_declaration14387 specparam_declaration_instance14387();
    specparam_declaration14388 specparam_declaration_instance14388();
    specparam_declaration14389 specparam_declaration_instance14389();
    specparam_declaration14390 specparam_declaration_instance14390();
    specparam_declaration14391 specparam_declaration_instance14391();
    specparam_declaration14392 specparam_declaration_instance14392();
    specparam_declaration14393 specparam_declaration_instance14393();
    specparam_declaration14394 specparam_declaration_instance14394();
    specparam_declaration14395 specparam_declaration_instance14395();
    specparam_declaration14396 specparam_declaration_instance14396();
    specparam_declaration14397 specparam_declaration_instance14397();
    specparam_declaration14398 specparam_declaration_instance14398();
    specparam_declaration14399 specparam_declaration_instance14399();
    specparam_declaration14400 specparam_declaration_instance14400();
    specparam_declaration14401 specparam_declaration_instance14401();
    specparam_declaration14402 specparam_declaration_instance14402();
    specparam_declaration14403 specparam_declaration_instance14403();
    specparam_declaration14404 specparam_declaration_instance14404();
    specparam_declaration14405 specparam_declaration_instance14405();
    specparam_declaration14406 specparam_declaration_instance14406();
    specparam_declaration14407 specparam_declaration_instance14407();
    specparam_declaration14408 specparam_declaration_instance14408();
    specparam_declaration14409 specparam_declaration_instance14409();
    specparam_declaration14410 specparam_declaration_instance14410();
    specparam_declaration14411 specparam_declaration_instance14411();
    specparam_declaration14412 specparam_declaration_instance14412();
    specparam_declaration14413 specparam_declaration_instance14413();
    specparam_declaration14414 specparam_declaration_instance14414();
    specparam_declaration14415 specparam_declaration_instance14415();
    specparam_declaration14416 specparam_declaration_instance14416();
    specparam_declaration14417 specparam_declaration_instance14417();
    specparam_declaration14418 specparam_declaration_instance14418();
    specparam_declaration14419 specparam_declaration_instance14419();
    specparam_declaration14420 specparam_declaration_instance14420();
    specparam_declaration14421 specparam_declaration_instance14421();
    specparam_declaration14422 specparam_declaration_instance14422();
    specparam_declaration14423 specparam_declaration_instance14423();
    specparam_declaration14424 specparam_declaration_instance14424();
    specparam_declaration14425 specparam_declaration_instance14425();
    specparam_declaration14426 specparam_declaration_instance14426();
    specparam_declaration14427 specparam_declaration_instance14427();
    specparam_declaration14428 specparam_declaration_instance14428();
    specparam_declaration14429 specparam_declaration_instance14429();
    specparam_declaration14430 specparam_declaration_instance14430();
    specparam_declaration14431 specparam_declaration_instance14431();
    specparam_declaration14432 specparam_declaration_instance14432();
    specparam_declaration14433 specparam_declaration_instance14433();
    specparam_declaration14434 specparam_declaration_instance14434();
    specparam_declaration14435 specparam_declaration_instance14435();
    specparam_declaration14436 specparam_declaration_instance14436();
    specparam_declaration14437 specparam_declaration_instance14437();
    specparam_declaration14438 specparam_declaration_instance14438();
    specparam_declaration14439 specparam_declaration_instance14439();
    specparam_declaration14440 specparam_declaration_instance14440();
    specparam_declaration14441 specparam_declaration_instance14441();
    specparam_declaration14442 specparam_declaration_instance14442();
    specparam_declaration14443 specparam_declaration_instance14443();
    specparam_declaration14444 specparam_declaration_instance14444();
    specparam_declaration14445 specparam_declaration_instance14445();
    specparam_declaration14446 specparam_declaration_instance14446();
    specparam_declaration14447 specparam_declaration_instance14447();
    specparam_declaration14448 specparam_declaration_instance14448();
    specparam_declaration14449 specparam_declaration_instance14449();
    specparam_declaration14450 specparam_declaration_instance14450();
    specparam_declaration14451 specparam_declaration_instance14451();
    specparam_declaration14452 specparam_declaration_instance14452();
    specparam_declaration14453 specparam_declaration_instance14453();
    specparam_declaration14454 specparam_declaration_instance14454();
    specparam_declaration14455 specparam_declaration_instance14455();
    specparam_declaration14456 specparam_declaration_instance14456();
    specparam_declaration14457 specparam_declaration_instance14457();
    specparam_declaration14458 specparam_declaration_instance14458();
    specparam_declaration14459 specparam_declaration_instance14459();
    specparam_declaration14460 specparam_declaration_instance14460();
    specparam_declaration14461 specparam_declaration_instance14461();
    specparam_declaration14462 specparam_declaration_instance14462();
    specparam_declaration14463 specparam_declaration_instance14463();
    specparam_declaration14464 specparam_declaration_instance14464();
    specparam_declaration14465 specparam_declaration_instance14465();
    specparam_declaration14466 specparam_declaration_instance14466();
    specparam_declaration14467 specparam_declaration_instance14467();
    specparam_declaration14468 specparam_declaration_instance14468();
    specparam_declaration14469 specparam_declaration_instance14469();
    specparam_declaration14470 specparam_declaration_instance14470();
    specparam_declaration14471 specparam_declaration_instance14471();
    specparam_declaration14472 specparam_declaration_instance14472();
    specparam_declaration14473 specparam_declaration_instance14473();
    specparam_declaration14474 specparam_declaration_instance14474();
    specparam_declaration14475 specparam_declaration_instance14475();
    specparam_declaration14476 specparam_declaration_instance14476();
    specparam_declaration14477 specparam_declaration_instance14477();
    specparam_declaration14478 specparam_declaration_instance14478();
    specparam_declaration14479 specparam_declaration_instance14479();
    specparam_declaration14480 specparam_declaration_instance14480();
    specparam_declaration14481 specparam_declaration_instance14481();
    specparam_declaration14482 specparam_declaration_instance14482();
    specparam_declaration14483 specparam_declaration_instance14483();
    specparam_declaration14484 specparam_declaration_instance14484();
    specparam_declaration14485 specparam_declaration_instance14485();
    specparam_declaration14486 specparam_declaration_instance14486();
    specparam_declaration14487 specparam_declaration_instance14487();
    specparam_declaration14488 specparam_declaration_instance14488();
    specparam_declaration14489 specparam_declaration_instance14489();
    specparam_declaration14490 specparam_declaration_instance14490();
    specparam_declaration14491 specparam_declaration_instance14491();
    specparam_declaration14492 specparam_declaration_instance14492();
    specparam_declaration14493 specparam_declaration_instance14493();
    specparam_declaration14494 specparam_declaration_instance14494();
    specparam_declaration14495 specparam_declaration_instance14495();
    specparam_declaration14496 specparam_declaration_instance14496();
    specparam_declaration14497 specparam_declaration_instance14497();
    specparam_declaration14498 specparam_declaration_instance14498();
    specparam_declaration14499 specparam_declaration_instance14499();
    specparam_declaration14500 specparam_declaration_instance14500();
    specparam_declaration14501 specparam_declaration_instance14501();
    specparam_declaration14502 specparam_declaration_instance14502();
    specparam_declaration14503 specparam_declaration_instance14503();
    specparam_declaration14504 specparam_declaration_instance14504();
    specparam_declaration14505 specparam_declaration_instance14505();
    specparam_declaration14506 specparam_declaration_instance14506();
    specparam_declaration14507 specparam_declaration_instance14507();
    specparam_declaration14508 specparam_declaration_instance14508();
    specparam_declaration14509 specparam_declaration_instance14509();
    specparam_declaration14510 specparam_declaration_instance14510();
    specparam_declaration14511 specparam_declaration_instance14511();
    specparam_declaration14512 specparam_declaration_instance14512();
    specparam_declaration14513 specparam_declaration_instance14513();
    specparam_declaration14514 specparam_declaration_instance14514();
    specparam_declaration14515 specparam_declaration_instance14515();
    specparam_declaration14516 specparam_declaration_instance14516();
    specparam_declaration14517 specparam_declaration_instance14517();
    specparam_declaration14518 specparam_declaration_instance14518();
    specparam_declaration14519 specparam_declaration_instance14519();
    specparam_declaration14520 specparam_declaration_instance14520();
    specparam_declaration14521 specparam_declaration_instance14521();
    specparam_declaration14522 specparam_declaration_instance14522();
    specparam_declaration14523 specparam_declaration_instance14523();
    specparam_declaration14524 specparam_declaration_instance14524();
    specparam_declaration14525 specparam_declaration_instance14525();
    specparam_declaration14526 specparam_declaration_instance14526();
    specparam_declaration14527 specparam_declaration_instance14527();
    specparam_declaration14528 specparam_declaration_instance14528();
    specparam_declaration14529 specparam_declaration_instance14529();
    specparam_declaration14530 specparam_declaration_instance14530();
    specparam_declaration14531 specparam_declaration_instance14531();
    specparam_declaration14532 specparam_declaration_instance14532();
    specparam_declaration14533 specparam_declaration_instance14533();
    specparam_declaration14534 specparam_declaration_instance14534();
    specparam_declaration14535 specparam_declaration_instance14535();
    specparam_declaration14536 specparam_declaration_instance14536();
    specparam_declaration14537 specparam_declaration_instance14537();
    specparam_declaration14538 specparam_declaration_instance14538();
    specparam_declaration14539 specparam_declaration_instance14539();
    specparam_declaration14540 specparam_declaration_instance14540();
    specparam_declaration14541 specparam_declaration_instance14541();
    specparam_declaration14542 specparam_declaration_instance14542();
    specparam_declaration14543 specparam_declaration_instance14543();
    specparam_declaration14544 specparam_declaration_instance14544();
    specparam_declaration14545 specparam_declaration_instance14545();
    specparam_declaration14546 specparam_declaration_instance14546();
    specparam_declaration14547 specparam_declaration_instance14547();
    specparam_declaration14548 specparam_declaration_instance14548();
    specparam_declaration14549 specparam_declaration_instance14549();
    specparam_declaration14550 specparam_declaration_instance14550();
    specparam_declaration14551 specparam_declaration_instance14551();
    specparam_declaration14552 specparam_declaration_instance14552();
    specparam_declaration14553 specparam_declaration_instance14553();
    specparam_declaration14554 specparam_declaration_instance14554();
    specparam_declaration14555 specparam_declaration_instance14555();
    specparam_declaration14556 specparam_declaration_instance14556();
    specparam_declaration14557 specparam_declaration_instance14557();
    specparam_declaration14558 specparam_declaration_instance14558();
    specparam_declaration14559 specparam_declaration_instance14559();
    specparam_declaration14560 specparam_declaration_instance14560();
    specparam_declaration14561 specparam_declaration_instance14561();
    specparam_declaration14562 specparam_declaration_instance14562();
    specparam_declaration14563 specparam_declaration_instance14563();
    specparam_declaration14564 specparam_declaration_instance14564();
    specparam_declaration14565 specparam_declaration_instance14565();
    specparam_declaration14566 specparam_declaration_instance14566();
    specparam_declaration14567 specparam_declaration_instance14567();
    specparam_declaration14568 specparam_declaration_instance14568();
    specparam_declaration14569 specparam_declaration_instance14569();
    specparam_declaration14570 specparam_declaration_instance14570();
    specparam_declaration14571 specparam_declaration_instance14571();
    specparam_declaration14572 specparam_declaration_instance14572();
    specparam_declaration14573 specparam_declaration_instance14573();
    specparam_declaration14574 specparam_declaration_instance14574();
    specparam_declaration14575 specparam_declaration_instance14575();
    specparam_declaration14576 specparam_declaration_instance14576();
    specparam_declaration14577 specparam_declaration_instance14577();
    specparam_declaration14578 specparam_declaration_instance14578();
    specparam_declaration14579 specparam_declaration_instance14579();
    specparam_declaration14580 specparam_declaration_instance14580();
    specparam_declaration14581 specparam_declaration_instance14581();
    specparam_declaration14582 specparam_declaration_instance14582();
    specparam_declaration14583 specparam_declaration_instance14583();
    specparam_declaration14584 specparam_declaration_instance14584();
    specparam_declaration14585 specparam_declaration_instance14585();
    specparam_declaration14586 specparam_declaration_instance14586();
    specparam_declaration14587 specparam_declaration_instance14587();
    specparam_declaration14588 specparam_declaration_instance14588();
    specparam_declaration14589 specparam_declaration_instance14589();
    specparam_declaration14590 specparam_declaration_instance14590();
    specparam_declaration14591 specparam_declaration_instance14591();
    specparam_declaration14592 specparam_declaration_instance14592();
    specparam_declaration14593 specparam_declaration_instance14593();
    specparam_declaration14594 specparam_declaration_instance14594();
    specparam_declaration14595 specparam_declaration_instance14595();
    specparam_declaration14596 specparam_declaration_instance14596();
    specparam_declaration14597 specparam_declaration_instance14597();
    specparam_declaration14598 specparam_declaration_instance14598();
    specparam_declaration14599 specparam_declaration_instance14599();
    specparam_declaration14600 specparam_declaration_instance14600();
    specparam_declaration14601 specparam_declaration_instance14601();
    specparam_declaration14602 specparam_declaration_instance14602();
    specparam_declaration14603 specparam_declaration_instance14603();
    specparam_declaration14604 specparam_declaration_instance14604();
    specparam_declaration14605 specparam_declaration_instance14605();
    specparam_declaration14606 specparam_declaration_instance14606();
    specparam_declaration14607 specparam_declaration_instance14607();
    specparam_declaration14608 specparam_declaration_instance14608();
    specparam_declaration14609 specparam_declaration_instance14609();
    specparam_declaration14610 specparam_declaration_instance14610();
    specparam_declaration14611 specparam_declaration_instance14611();
    specparam_declaration14612 specparam_declaration_instance14612();
    specparam_declaration14613 specparam_declaration_instance14613();
    specparam_declaration14614 specparam_declaration_instance14614();
    specparam_declaration14615 specparam_declaration_instance14615();
    specparam_declaration14616 specparam_declaration_instance14616();
    specparam_declaration14617 specparam_declaration_instance14617();
    specparam_declaration14618 specparam_declaration_instance14618();
    specparam_declaration14619 specparam_declaration_instance14619();
    specparam_declaration14620 specparam_declaration_instance14620();
    specparam_declaration14621 specparam_declaration_instance14621();
    specparam_declaration14622 specparam_declaration_instance14622();
    specparam_declaration14623 specparam_declaration_instance14623();
    specparam_declaration14624 specparam_declaration_instance14624();
    specparam_declaration14625 specparam_declaration_instance14625();
    specparam_declaration14626 specparam_declaration_instance14626();
    specparam_declaration14627 specparam_declaration_instance14627();
    specparam_declaration14628 specparam_declaration_instance14628();
    specparam_declaration14629 specparam_declaration_instance14629();
    specparam_declaration14630 specparam_declaration_instance14630();
    specparam_declaration14631 specparam_declaration_instance14631();
    specparam_declaration14632 specparam_declaration_instance14632();
    specparam_declaration14633 specparam_declaration_instance14633();
    specparam_declaration14634 specparam_declaration_instance14634();
    specparam_declaration14635 specparam_declaration_instance14635();
    specparam_declaration14636 specparam_declaration_instance14636();
    specparam_declaration14637 specparam_declaration_instance14637();
    specparam_declaration14638 specparam_declaration_instance14638();
    specparam_declaration14639 specparam_declaration_instance14639();
    specparam_declaration14640 specparam_declaration_instance14640();
    specparam_declaration14641 specparam_declaration_instance14641();
    specparam_declaration14642 specparam_declaration_instance14642();
    specparam_declaration14643 specparam_declaration_instance14643();
    specparam_declaration14644 specparam_declaration_instance14644();
    specparam_declaration14645 specparam_declaration_instance14645();
    specparam_declaration14646 specparam_declaration_instance14646();
    specparam_declaration14647 specparam_declaration_instance14647();
    specparam_declaration14648 specparam_declaration_instance14648();
    specparam_declaration14649 specparam_declaration_instance14649();
    specparam_declaration14650 specparam_declaration_instance14650();
    specparam_declaration14651 specparam_declaration_instance14651();
    specparam_declaration14652 specparam_declaration_instance14652();
    specparam_declaration14653 specparam_declaration_instance14653();
    specparam_declaration14654 specparam_declaration_instance14654();
    specparam_declaration14655 specparam_declaration_instance14655();
    specparam_declaration14656 specparam_declaration_instance14656();
    specparam_declaration14657 specparam_declaration_instance14657();
    specparam_declaration14658 specparam_declaration_instance14658();
    specparam_declaration14659 specparam_declaration_instance14659();
    specparam_declaration14660 specparam_declaration_instance14660();
    specparam_declaration14661 specparam_declaration_instance14661();
    specparam_declaration14662 specparam_declaration_instance14662();
    specparam_declaration14663 specparam_declaration_instance14663();
    specparam_declaration14664 specparam_declaration_instance14664();
    specparam_declaration14665 specparam_declaration_instance14665();
    specparam_declaration14666 specparam_declaration_instance14666();
    specparam_declaration14667 specparam_declaration_instance14667();
    specparam_declaration14668 specparam_declaration_instance14668();
    specparam_declaration14669 specparam_declaration_instance14669();
    specparam_declaration14670 specparam_declaration_instance14670();
    specparam_declaration14671 specparam_declaration_instance14671();
    specparam_declaration14672 specparam_declaration_instance14672();
    specparam_declaration14673 specparam_declaration_instance14673();
    specparam_declaration14674 specparam_declaration_instance14674();
    specparam_declaration14675 specparam_declaration_instance14675();
    specparam_declaration14676 specparam_declaration_instance14676();
    specparam_declaration14677 specparam_declaration_instance14677();
    specparam_declaration14678 specparam_declaration_instance14678();
    specparam_declaration14679 specparam_declaration_instance14679();
    specparam_declaration14680 specparam_declaration_instance14680();
    specparam_declaration14681 specparam_declaration_instance14681();
    specparam_declaration14682 specparam_declaration_instance14682();
    specparam_declaration14683 specparam_declaration_instance14683();
    specparam_declaration14684 specparam_declaration_instance14684();
    specparam_declaration14685 specparam_declaration_instance14685();
    specparam_declaration14686 specparam_declaration_instance14686();
    specparam_declaration14687 specparam_declaration_instance14687();
    specparam_declaration14688 specparam_declaration_instance14688();
    specparam_declaration14689 specparam_declaration_instance14689();
    specparam_declaration14690 specparam_declaration_instance14690();
    specparam_declaration14691 specparam_declaration_instance14691();
    specparam_declaration14692 specparam_declaration_instance14692();
    specparam_declaration14693 specparam_declaration_instance14693();
    specparam_declaration14694 specparam_declaration_instance14694();
    specparam_declaration14695 specparam_declaration_instance14695();
    specparam_declaration14696 specparam_declaration_instance14696();
    specparam_declaration14697 specparam_declaration_instance14697();
    specparam_declaration14698 specparam_declaration_instance14698();
    specparam_declaration14699 specparam_declaration_instance14699();
    specparam_declaration14700 specparam_declaration_instance14700();
    specparam_declaration14701 specparam_declaration_instance14701();
    specparam_declaration14702 specparam_declaration_instance14702();
    specparam_declaration14703 specparam_declaration_instance14703();
    specparam_declaration14704 specparam_declaration_instance14704();
    specparam_declaration14705 specparam_declaration_instance14705();
    specparam_declaration14706 specparam_declaration_instance14706();
    specparam_declaration14707 specparam_declaration_instance14707();
    specparam_declaration14708 specparam_declaration_instance14708();
    specparam_declaration14709 specparam_declaration_instance14709();
    specparam_declaration14710 specparam_declaration_instance14710();
    specparam_declaration14711 specparam_declaration_instance14711();
    specparam_declaration14712 specparam_declaration_instance14712();
    specparam_declaration14713 specparam_declaration_instance14713();
    specparam_declaration14714 specparam_declaration_instance14714();
    specparam_declaration14715 specparam_declaration_instance14715();
    specparam_declaration14716 specparam_declaration_instance14716();
    specparam_declaration14717 specparam_declaration_instance14717();
    specparam_declaration14718 specparam_declaration_instance14718();
    specparam_declaration14719 specparam_declaration_instance14719();
    specparam_declaration14720 specparam_declaration_instance14720();
    specparam_declaration14721 specparam_declaration_instance14721();
    specparam_declaration14722 specparam_declaration_instance14722();
    specparam_declaration14723 specparam_declaration_instance14723();
    specparam_declaration14724 specparam_declaration_instance14724();
    specparam_declaration14725 specparam_declaration_instance14725();
    specparam_declaration14726 specparam_declaration_instance14726();
    specparam_declaration14727 specparam_declaration_instance14727();
    specparam_declaration14728 specparam_declaration_instance14728();
    specparam_declaration14729 specparam_declaration_instance14729();
    specparam_declaration14730 specparam_declaration_instance14730();
    specparam_declaration14731 specparam_declaration_instance14731();
    specparam_declaration14732 specparam_declaration_instance14732();
    specparam_declaration14733 specparam_declaration_instance14733();
    specparam_declaration14734 specparam_declaration_instance14734();
    specparam_declaration14735 specparam_declaration_instance14735();
    specparam_declaration14736 specparam_declaration_instance14736();
    specparam_declaration14737 specparam_declaration_instance14737();
    specparam_declaration14738 specparam_declaration_instance14738();
    specparam_declaration14739 specparam_declaration_instance14739();
    specparam_declaration14740 specparam_declaration_instance14740();
    specparam_declaration14741 specparam_declaration_instance14741();
    specparam_declaration14742 specparam_declaration_instance14742();
    specparam_declaration14743 specparam_declaration_instance14743();
    specparam_declaration14744 specparam_declaration_instance14744();
    specparam_declaration14745 specparam_declaration_instance14745();
    specparam_declaration14746 specparam_declaration_instance14746();
    specparam_declaration14747 specparam_declaration_instance14747();
    specparam_declaration14748 specparam_declaration_instance14748();
    specparam_declaration14749 specparam_declaration_instance14749();
    specparam_declaration14750 specparam_declaration_instance14750();
    specparam_declaration14751 specparam_declaration_instance14751();
    specparam_declaration14752 specparam_declaration_instance14752();
    specparam_declaration14753 specparam_declaration_instance14753();
    specparam_declaration14754 specparam_declaration_instance14754();
    specparam_declaration14755 specparam_declaration_instance14755();
    specparam_declaration14756 specparam_declaration_instance14756();
    specparam_declaration14757 specparam_declaration_instance14757();
    specparam_declaration14758 specparam_declaration_instance14758();
    specparam_declaration14759 specparam_declaration_instance14759();
    specparam_declaration14760 specparam_declaration_instance14760();
    specparam_declaration14761 specparam_declaration_instance14761();
    specparam_declaration14762 specparam_declaration_instance14762();
    specparam_declaration14763 specparam_declaration_instance14763();
    specparam_declaration14764 specparam_declaration_instance14764();
    specparam_declaration14765 specparam_declaration_instance14765();
    specparam_declaration14766 specparam_declaration_instance14766();
    specparam_declaration14767 specparam_declaration_instance14767();
    specparam_declaration14768 specparam_declaration_instance14768();
    specparam_declaration14769 specparam_declaration_instance14769();
    specparam_declaration14770 specparam_declaration_instance14770();
    specparam_declaration14771 specparam_declaration_instance14771();
    specparam_declaration14772 specparam_declaration_instance14772();
    specparam_declaration14773 specparam_declaration_instance14773();
    specparam_declaration14774 specparam_declaration_instance14774();
    specparam_declaration14775 specparam_declaration_instance14775();
    specparam_declaration14776 specparam_declaration_instance14776();
    specparam_declaration14777 specparam_declaration_instance14777();
    specparam_declaration14778 specparam_declaration_instance14778();
    specparam_declaration14779 specparam_declaration_instance14779();
    specparam_declaration14780 specparam_declaration_instance14780();
    specparam_declaration14781 specparam_declaration_instance14781();
    specparam_declaration14782 specparam_declaration_instance14782();
    specparam_declaration14783 specparam_declaration_instance14783();
    specparam_declaration14784 specparam_declaration_instance14784();
    specparam_declaration14785 specparam_declaration_instance14785();
    specparam_declaration14786 specparam_declaration_instance14786();
    specparam_declaration14787 specparam_declaration_instance14787();
    specparam_declaration14788 specparam_declaration_instance14788();
    specparam_declaration14789 specparam_declaration_instance14789();
    specparam_declaration14790 specparam_declaration_instance14790();
    specparam_declaration14791 specparam_declaration_instance14791();
    specparam_declaration14792 specparam_declaration_instance14792();
    specparam_declaration14793 specparam_declaration_instance14793();
    specparam_declaration14794 specparam_declaration_instance14794();
    specparam_declaration14795 specparam_declaration_instance14795();
    specparam_declaration14796 specparam_declaration_instance14796();
    specparam_declaration14797 specparam_declaration_instance14797();
    specparam_declaration14798 specparam_declaration_instance14798();
    specparam_declaration14799 specparam_declaration_instance14799();
    specparam_declaration14800 specparam_declaration_instance14800();
    specparam_declaration14801 specparam_declaration_instance14801();
    specparam_declaration14802 specparam_declaration_instance14802();
    specparam_declaration14803 specparam_declaration_instance14803();
    specparam_declaration14804 specparam_declaration_instance14804();
    specparam_declaration14805 specparam_declaration_instance14805();
    specparam_declaration14806 specparam_declaration_instance14806();
    specparam_declaration14807 specparam_declaration_instance14807();
    specparam_declaration14808 specparam_declaration_instance14808();
    specparam_declaration14809 specparam_declaration_instance14809();
    specparam_declaration14810 specparam_declaration_instance14810();
    specparam_declaration14811 specparam_declaration_instance14811();
    specparam_declaration14812 specparam_declaration_instance14812();
    specparam_declaration14813 specparam_declaration_instance14813();
    specparam_declaration14814 specparam_declaration_instance14814();
    specparam_declaration14815 specparam_declaration_instance14815();
    specparam_declaration14816 specparam_declaration_instance14816();
    specparam_declaration14817 specparam_declaration_instance14817();
    specparam_declaration14818 specparam_declaration_instance14818();
    specparam_declaration14819 specparam_declaration_instance14819();
    specparam_declaration14820 specparam_declaration_instance14820();
    specparam_declaration14821 specparam_declaration_instance14821();
    specparam_declaration14822 specparam_declaration_instance14822();
    specparam_declaration14823 specparam_declaration_instance14823();
    specparam_declaration14824 specparam_declaration_instance14824();
    specparam_declaration14825 specparam_declaration_instance14825();
    specparam_declaration14826 specparam_declaration_instance14826();
    specparam_declaration14827 specparam_declaration_instance14827();
    specparam_declaration14828 specparam_declaration_instance14828();
    specparam_declaration14829 specparam_declaration_instance14829();
    specparam_declaration14830 specparam_declaration_instance14830();
    specparam_declaration14831 specparam_declaration_instance14831();
    specparam_declaration14832 specparam_declaration_instance14832();
    specparam_declaration14833 specparam_declaration_instance14833();
    specparam_declaration14834 specparam_declaration_instance14834();
    specparam_declaration14835 specparam_declaration_instance14835();
    specparam_declaration14836 specparam_declaration_instance14836();
    specparam_declaration14837 specparam_declaration_instance14837();
    specparam_declaration14838 specparam_declaration_instance14838();
    specparam_declaration14839 specparam_declaration_instance14839();
    specparam_declaration14840 specparam_declaration_instance14840();
    specparam_declaration14841 specparam_declaration_instance14841();
    specparam_declaration14842 specparam_declaration_instance14842();
    specparam_declaration14843 specparam_declaration_instance14843();
    specparam_declaration14844 specparam_declaration_instance14844();
    specparam_declaration14845 specparam_declaration_instance14845();
    specparam_declaration14846 specparam_declaration_instance14846();
    specparam_declaration14847 specparam_declaration_instance14847();
    specparam_declaration14848 specparam_declaration_instance14848();
    specparam_declaration14849 specparam_declaration_instance14849();
    specparam_declaration14850 specparam_declaration_instance14850();
    specparam_declaration14851 specparam_declaration_instance14851();
    specparam_declaration14852 specparam_declaration_instance14852();
    specparam_declaration14853 specparam_declaration_instance14853();
    specparam_declaration14854 specparam_declaration_instance14854();
    specparam_declaration14855 specparam_declaration_instance14855();
    specparam_declaration14856 specparam_declaration_instance14856();
    specparam_declaration14857 specparam_declaration_instance14857();
    specparam_declaration14858 specparam_declaration_instance14858();
    specparam_declaration14859 specparam_declaration_instance14859();
    specparam_declaration14860 specparam_declaration_instance14860();
    specparam_declaration14861 specparam_declaration_instance14861();
    specparam_declaration14862 specparam_declaration_instance14862();
    specparam_declaration14863 specparam_declaration_instance14863();
    specparam_declaration14864 specparam_declaration_instance14864();
    specparam_declaration14865 specparam_declaration_instance14865();
    specparam_declaration14866 specparam_declaration_instance14866();
    specparam_declaration14867 specparam_declaration_instance14867();
    specparam_declaration14868 specparam_declaration_instance14868();
    specparam_declaration14869 specparam_declaration_instance14869();
    specparam_declaration14870 specparam_declaration_instance14870();
    specparam_declaration14871 specparam_declaration_instance14871();
    specparam_declaration14872 specparam_declaration_instance14872();
    specparam_declaration14873 specparam_declaration_instance14873();
    specparam_declaration14874 specparam_declaration_instance14874();
    specparam_declaration14875 specparam_declaration_instance14875();
    specparam_declaration14876 specparam_declaration_instance14876();
    specparam_declaration14877 specparam_declaration_instance14877();
    specparam_declaration14878 specparam_declaration_instance14878();
    specparam_declaration14879 specparam_declaration_instance14879();
    specparam_declaration14880 specparam_declaration_instance14880();
    specparam_declaration14881 specparam_declaration_instance14881();
    specparam_declaration14882 specparam_declaration_instance14882();
    specparam_declaration14883 specparam_declaration_instance14883();
    specparam_declaration14884 specparam_declaration_instance14884();
    specparam_declaration14885 specparam_declaration_instance14885();
    specparam_declaration14886 specparam_declaration_instance14886();
    specparam_declaration14887 specparam_declaration_instance14887();
    specparam_declaration14888 specparam_declaration_instance14888();
    specparam_declaration14889 specparam_declaration_instance14889();
    specparam_declaration14890 specparam_declaration_instance14890();
    specparam_declaration14891 specparam_declaration_instance14891();
    specparam_declaration14892 specparam_declaration_instance14892();
    specparam_declaration14893 specparam_declaration_instance14893();
    specparam_declaration14894 specparam_declaration_instance14894();
    specparam_declaration14895 specparam_declaration_instance14895();
    specparam_declaration14896 specparam_declaration_instance14896();
    specparam_declaration14897 specparam_declaration_instance14897();
    specparam_declaration14898 specparam_declaration_instance14898();
    specparam_declaration14899 specparam_declaration_instance14899();
    specparam_declaration14900 specparam_declaration_instance14900();
    specparam_declaration14901 specparam_declaration_instance14901();
    specparam_declaration14902 specparam_declaration_instance14902();
    specparam_declaration14903 specparam_declaration_instance14903();
    specparam_declaration14904 specparam_declaration_instance14904();
    specparam_declaration14905 specparam_declaration_instance14905();
    specparam_declaration14906 specparam_declaration_instance14906();
    specparam_declaration14907 specparam_declaration_instance14907();
    specparam_declaration14908 specparam_declaration_instance14908();
    specparam_declaration14909 specparam_declaration_instance14909();
    specparam_declaration14910 specparam_declaration_instance14910();
    specparam_declaration14911 specparam_declaration_instance14911();
    specparam_declaration14912 specparam_declaration_instance14912();
    specparam_declaration14913 specparam_declaration_instance14913();
    specparam_declaration14914 specparam_declaration_instance14914();
    specparam_declaration14915 specparam_declaration_instance14915();
    specparam_declaration14916 specparam_declaration_instance14916();
    specparam_declaration14917 specparam_declaration_instance14917();
    specparam_declaration14918 specparam_declaration_instance14918();
    specparam_declaration14919 specparam_declaration_instance14919();
    specparam_declaration14920 specparam_declaration_instance14920();
    specparam_declaration14921 specparam_declaration_instance14921();
    specparam_declaration14922 specparam_declaration_instance14922();
    specparam_declaration14923 specparam_declaration_instance14923();
    specparam_declaration14924 specparam_declaration_instance14924();
    specparam_declaration14925 specparam_declaration_instance14925();
    specparam_declaration14926 specparam_declaration_instance14926();
    specparam_declaration14927 specparam_declaration_instance14927();
    specparam_declaration14928 specparam_declaration_instance14928();
    specparam_declaration14929 specparam_declaration_instance14929();
    specparam_declaration14930 specparam_declaration_instance14930();
    specparam_declaration14931 specparam_declaration_instance14931();
    specparam_declaration14932 specparam_declaration_instance14932();
    specparam_declaration14933 specparam_declaration_instance14933();
    specparam_declaration14934 specparam_declaration_instance14934();
    specparam_declaration14935 specparam_declaration_instance14935();
    specparam_declaration14936 specparam_declaration_instance14936();
    specparam_declaration14937 specparam_declaration_instance14937();
    specparam_declaration14938 specparam_declaration_instance14938();
    specparam_declaration14939 specparam_declaration_instance14939();
    specparam_declaration14940 specparam_declaration_instance14940();
    specparam_declaration14941 specparam_declaration_instance14941();
    specparam_declaration14942 specparam_declaration_instance14942();
    specparam_declaration14943 specparam_declaration_instance14943();
    specparam_declaration14944 specparam_declaration_instance14944();
    specparam_declaration14945 specparam_declaration_instance14945();
    specparam_declaration14946 specparam_declaration_instance14946();
    specparam_declaration14947 specparam_declaration_instance14947();
    specparam_declaration14948 specparam_declaration_instance14948();
    specparam_declaration14949 specparam_declaration_instance14949();
    specparam_declaration14950 specparam_declaration_instance14950();
    specparam_declaration14951 specparam_declaration_instance14951();
    specparam_declaration14952 specparam_declaration_instance14952();
    specparam_declaration14953 specparam_declaration_instance14953();
    specparam_declaration14954 specparam_declaration_instance14954();
    specparam_declaration14955 specparam_declaration_instance14955();
    specparam_declaration14956 specparam_declaration_instance14956();
    specparam_declaration14957 specparam_declaration_instance14957();
    specparam_declaration14958 specparam_declaration_instance14958();
    specparam_declaration14959 specparam_declaration_instance14959();
    specparam_declaration14960 specparam_declaration_instance14960();
    specparam_declaration14961 specparam_declaration_instance14961();
    specparam_declaration14962 specparam_declaration_instance14962();
    specparam_declaration14963 specparam_declaration_instance14963();
    specparam_declaration14964 specparam_declaration_instance14964();
    specparam_declaration14965 specparam_declaration_instance14965();
    specparam_declaration14966 specparam_declaration_instance14966();
    specparam_declaration14967 specparam_declaration_instance14967();
    specparam_declaration14968 specparam_declaration_instance14968();
    specparam_declaration14969 specparam_declaration_instance14969();
    specparam_declaration14970 specparam_declaration_instance14970();
    specparam_declaration14971 specparam_declaration_instance14971();
    specparam_declaration14972 specparam_declaration_instance14972();
    specparam_declaration14973 specparam_declaration_instance14973();
    specparam_declaration14974 specparam_declaration_instance14974();
    specparam_declaration14975 specparam_declaration_instance14975();
    specparam_declaration14976 specparam_declaration_instance14976();
    specparam_declaration14977 specparam_declaration_instance14977();
    specparam_declaration14978 specparam_declaration_instance14978();
    specparam_declaration14979 specparam_declaration_instance14979();
    specparam_declaration14980 specparam_declaration_instance14980();
    specparam_declaration14981 specparam_declaration_instance14981();
    specparam_declaration14982 specparam_declaration_instance14982();
    specparam_declaration14983 specparam_declaration_instance14983();
    specparam_declaration14984 specparam_declaration_instance14984();
    specparam_declaration14985 specparam_declaration_instance14985();
    specparam_declaration14986 specparam_declaration_instance14986();
    specparam_declaration14987 specparam_declaration_instance14987();
    specparam_declaration14988 specparam_declaration_instance14988();
    specparam_declaration14989 specparam_declaration_instance14989();
    specparam_declaration14990 specparam_declaration_instance14990();
    specparam_declaration14991 specparam_declaration_instance14991();
    specparam_declaration14992 specparam_declaration_instance14992();
    specparam_declaration14993 specparam_declaration_instance14993();
    specparam_declaration14994 specparam_declaration_instance14994();
    specparam_declaration14995 specparam_declaration_instance14995();
    specparam_declaration14996 specparam_declaration_instance14996();
    specparam_declaration14997 specparam_declaration_instance14997();
    specparam_declaration14998 specparam_declaration_instance14998();
    specparam_declaration14999 specparam_declaration_instance14999();
    specparam_declaration15000 specparam_declaration_instance15000();
    specparam_declaration15001 specparam_declaration_instance15001();
    specparam_declaration15002 specparam_declaration_instance15002();
    specparam_declaration15003 specparam_declaration_instance15003();
    specparam_declaration15004 specparam_declaration_instance15004();
    specparam_declaration15005 specparam_declaration_instance15005();
    specparam_declaration15006 specparam_declaration_instance15006();
    specparam_declaration15007 specparam_declaration_instance15007();
    specparam_declaration15008 specparam_declaration_instance15008();
    specparam_declaration15009 specparam_declaration_instance15009();
    specparam_declaration15010 specparam_declaration_instance15010();
    specparam_declaration15011 specparam_declaration_instance15011();
    specparam_declaration15012 specparam_declaration_instance15012();
    specparam_declaration15013 specparam_declaration_instance15013();
    specparam_declaration15014 specparam_declaration_instance15014();
    specparam_declaration15015 specparam_declaration_instance15015();
    specparam_declaration15016 specparam_declaration_instance15016();
    specparam_declaration15017 specparam_declaration_instance15017();
    specparam_declaration15018 specparam_declaration_instance15018();
    specparam_declaration15019 specparam_declaration_instance15019();
    specparam_declaration15020 specparam_declaration_instance15020();
    specparam_declaration15021 specparam_declaration_instance15021();
    specparam_declaration15022 specparam_declaration_instance15022();
    specparam_declaration15023 specparam_declaration_instance15023();
    specparam_declaration15024 specparam_declaration_instance15024();
    specparam_declaration15025 specparam_declaration_instance15025();
    specparam_declaration15026 specparam_declaration_instance15026();
    specparam_declaration15027 specparam_declaration_instance15027();
    specparam_declaration15028 specparam_declaration_instance15028();
    specparam_declaration15029 specparam_declaration_instance15029();
    specparam_declaration15030 specparam_declaration_instance15030();
    specparam_declaration15031 specparam_declaration_instance15031();
    specparam_declaration15032 specparam_declaration_instance15032();
    specparam_declaration15033 specparam_declaration_instance15033();
    specparam_declaration15034 specparam_declaration_instance15034();
    specparam_declaration15035 specparam_declaration_instance15035();
    specparam_declaration15036 specparam_declaration_instance15036();
    specparam_declaration15037 specparam_declaration_instance15037();
    specparam_declaration15038 specparam_declaration_instance15038();
    specparam_declaration15039 specparam_declaration_instance15039();
    specparam_declaration15040 specparam_declaration_instance15040();
    specparam_declaration15041 specparam_declaration_instance15041();
    specparam_declaration15042 specparam_declaration_instance15042();
    specparam_declaration15043 specparam_declaration_instance15043();
    specparam_declaration15044 specparam_declaration_instance15044();
    specparam_declaration15045 specparam_declaration_instance15045();
    specparam_declaration15046 specparam_declaration_instance15046();
    specparam_declaration15047 specparam_declaration_instance15047();
    specparam_declaration15048 specparam_declaration_instance15048();
    specparam_declaration15049 specparam_declaration_instance15049();
    specparam_declaration15050 specparam_declaration_instance15050();
    specparam_declaration15051 specparam_declaration_instance15051();
    specparam_declaration15052 specparam_declaration_instance15052();
    specparam_declaration15053 specparam_declaration_instance15053();
    specparam_declaration15054 specparam_declaration_instance15054();
    specparam_declaration15055 specparam_declaration_instance15055();
    specparam_declaration15056 specparam_declaration_instance15056();
    specparam_declaration15057 specparam_declaration_instance15057();
    specparam_declaration15058 specparam_declaration_instance15058();
    specparam_declaration15059 specparam_declaration_instance15059();
    specparam_declaration15060 specparam_declaration_instance15060();
    specparam_declaration15061 specparam_declaration_instance15061();
    specparam_declaration15062 specparam_declaration_instance15062();
    specparam_declaration15063 specparam_declaration_instance15063();
    specparam_declaration15064 specparam_declaration_instance15064();
    specparam_declaration15065 specparam_declaration_instance15065();
    specparam_declaration15066 specparam_declaration_instance15066();
    specparam_declaration15067 specparam_declaration_instance15067();
    specparam_declaration15068 specparam_declaration_instance15068();
    specparam_declaration15069 specparam_declaration_instance15069();
    specparam_declaration15070 specparam_declaration_instance15070();
    specparam_declaration15071 specparam_declaration_instance15071();
    specparam_declaration15072 specparam_declaration_instance15072();
    specparam_declaration15073 specparam_declaration_instance15073();
    specparam_declaration15074 specparam_declaration_instance15074();
    specparam_declaration15075 specparam_declaration_instance15075();
    specparam_declaration15076 specparam_declaration_instance15076();
    specparam_declaration15077 specparam_declaration_instance15077();
    specparam_declaration15078 specparam_declaration_instance15078();
    specparam_declaration15079 specparam_declaration_instance15079();
    specparam_declaration15080 specparam_declaration_instance15080();
    specparam_declaration15081 specparam_declaration_instance15081();
    specparam_declaration15082 specparam_declaration_instance15082();
    specparam_declaration15083 specparam_declaration_instance15083();
    specparam_declaration15084 specparam_declaration_instance15084();
    specparam_declaration15085 specparam_declaration_instance15085();
    specparam_declaration15086 specparam_declaration_instance15086();
    specparam_declaration15087 specparam_declaration_instance15087();
    specparam_declaration15088 specparam_declaration_instance15088();
    specparam_declaration15089 specparam_declaration_instance15089();
    specparam_declaration15090 specparam_declaration_instance15090();
    specparam_declaration15091 specparam_declaration_instance15091();
    specparam_declaration15092 specparam_declaration_instance15092();
    specparam_declaration15093 specparam_declaration_instance15093();
    specparam_declaration15094 specparam_declaration_instance15094();
    specparam_declaration15095 specparam_declaration_instance15095();
    specparam_declaration15096 specparam_declaration_instance15096();
    specparam_declaration15097 specparam_declaration_instance15097();
    specparam_declaration15098 specparam_declaration_instance15098();
    specparam_declaration15099 specparam_declaration_instance15099();
    specparam_declaration15100 specparam_declaration_instance15100();
    specparam_declaration15101 specparam_declaration_instance15101();
    specparam_declaration15102 specparam_declaration_instance15102();
    specparam_declaration15103 specparam_declaration_instance15103();
    specparam_declaration15104 specparam_declaration_instance15104();
    specparam_declaration15105 specparam_declaration_instance15105();
    specparam_declaration15106 specparam_declaration_instance15106();
    specparam_declaration15107 specparam_declaration_instance15107();
    specparam_declaration15108 specparam_declaration_instance15108();
    specparam_declaration15109 specparam_declaration_instance15109();
    specparam_declaration15110 specparam_declaration_instance15110();
    specparam_declaration15111 specparam_declaration_instance15111();
    specparam_declaration15112 specparam_declaration_instance15112();
    specparam_declaration15113 specparam_declaration_instance15113();
    specparam_declaration15114 specparam_declaration_instance15114();
    specparam_declaration15115 specparam_declaration_instance15115();
    specparam_declaration15116 specparam_declaration_instance15116();
    specparam_declaration15117 specparam_declaration_instance15117();
    specparam_declaration15118 specparam_declaration_instance15118();
    specparam_declaration15119 specparam_declaration_instance15119();
    specparam_declaration15120 specparam_declaration_instance15120();
    specparam_declaration15121 specparam_declaration_instance15121();
    specparam_declaration15122 specparam_declaration_instance15122();
    specparam_declaration15123 specparam_declaration_instance15123();
    specparam_declaration15124 specparam_declaration_instance15124();
    specparam_declaration15125 specparam_declaration_instance15125();
    specparam_declaration15126 specparam_declaration_instance15126();
    specparam_declaration15127 specparam_declaration_instance15127();
    specparam_declaration15128 specparam_declaration_instance15128();
    specparam_declaration15129 specparam_declaration_instance15129();
    specparam_declaration15130 specparam_declaration_instance15130();
    specparam_declaration15131 specparam_declaration_instance15131();
    specparam_declaration15132 specparam_declaration_instance15132();
    specparam_declaration15133 specparam_declaration_instance15133();
    specparam_declaration15134 specparam_declaration_instance15134();
    specparam_declaration15135 specparam_declaration_instance15135();
    specparam_declaration15136 specparam_declaration_instance15136();
    specparam_declaration15137 specparam_declaration_instance15137();
    specparam_declaration15138 specparam_declaration_instance15138();
    specparam_declaration15139 specparam_declaration_instance15139();
    specparam_declaration15140 specparam_declaration_instance15140();
    specparam_declaration15141 specparam_declaration_instance15141();
    specparam_declaration15142 specparam_declaration_instance15142();
    specparam_declaration15143 specparam_declaration_instance15143();
    specparam_declaration15144 specparam_declaration_instance15144();
    specparam_declaration15145 specparam_declaration_instance15145();
    specparam_declaration15146 specparam_declaration_instance15146();
    specparam_declaration15147 specparam_declaration_instance15147();
    specparam_declaration15148 specparam_declaration_instance15148();
    specparam_declaration15149 specparam_declaration_instance15149();
    specparam_declaration15150 specparam_declaration_instance15150();
    specparam_declaration15151 specparam_declaration_instance15151();
    specparam_declaration15152 specparam_declaration_instance15152();
    specparam_declaration15153 specparam_declaration_instance15153();
    specparam_declaration15154 specparam_declaration_instance15154();
    specparam_declaration15155 specparam_declaration_instance15155();
    specparam_declaration15156 specparam_declaration_instance15156();
    specparam_declaration15157 specparam_declaration_instance15157();
    specparam_declaration15158 specparam_declaration_instance15158();
    specparam_declaration15159 specparam_declaration_instance15159();
    specparam_declaration15160 specparam_declaration_instance15160();
    specparam_declaration15161 specparam_declaration_instance15161();
    specparam_declaration15162 specparam_declaration_instance15162();
    specparam_declaration15163 specparam_declaration_instance15163();
    specparam_declaration15164 specparam_declaration_instance15164();
    specparam_declaration15165 specparam_declaration_instance15165();
    specparam_declaration15166 specparam_declaration_instance15166();
    specparam_declaration15167 specparam_declaration_instance15167();
    specparam_declaration15168 specparam_declaration_instance15168();
    specparam_declaration15169 specparam_declaration_instance15169();
    specparam_declaration15170 specparam_declaration_instance15170();
    specparam_declaration15171 specparam_declaration_instance15171();
    specparam_declaration15172 specparam_declaration_instance15172();
    specparam_declaration15173 specparam_declaration_instance15173();
    specparam_declaration15174 specparam_declaration_instance15174();
    specparam_declaration15175 specparam_declaration_instance15175();
    specparam_declaration15176 specparam_declaration_instance15176();
    specparam_declaration15177 specparam_declaration_instance15177();
    specparam_declaration15178 specparam_declaration_instance15178();
    specparam_declaration15179 specparam_declaration_instance15179();
    specparam_declaration15180 specparam_declaration_instance15180();
    specparam_declaration15181 specparam_declaration_instance15181();
    specparam_declaration15182 specparam_declaration_instance15182();
    specparam_declaration15183 specparam_declaration_instance15183();
    specparam_declaration15184 specparam_declaration_instance15184();
    specparam_declaration15185 specparam_declaration_instance15185();
    specparam_declaration15186 specparam_declaration_instance15186();
    specparam_declaration15187 specparam_declaration_instance15187();
    specparam_declaration15188 specparam_declaration_instance15188();
    specparam_declaration15189 specparam_declaration_instance15189();
    specparam_declaration15190 specparam_declaration_instance15190();
    specparam_declaration15191 specparam_declaration_instance15191();
    specparam_declaration15192 specparam_declaration_instance15192();
    specparam_declaration15193 specparam_declaration_instance15193();
    specparam_declaration15194 specparam_declaration_instance15194();
    specparam_declaration15195 specparam_declaration_instance15195();
    specparam_declaration15196 specparam_declaration_instance15196();
    specparam_declaration15197 specparam_declaration_instance15197();
    specparam_declaration15198 specparam_declaration_instance15198();
    specparam_declaration15199 specparam_declaration_instance15199();
    specparam_declaration15200 specparam_declaration_instance15200();
    specparam_declaration15201 specparam_declaration_instance15201();
    specparam_declaration15202 specparam_declaration_instance15202();
    specparam_declaration15203 specparam_declaration_instance15203();
    specparam_declaration15204 specparam_declaration_instance15204();
    specparam_declaration15205 specparam_declaration_instance15205();
    specparam_declaration15206 specparam_declaration_instance15206();
    specparam_declaration15207 specparam_declaration_instance15207();
    specparam_declaration15208 specparam_declaration_instance15208();
    specparam_declaration15209 specparam_declaration_instance15209();
    specparam_declaration15210 specparam_declaration_instance15210();
    specparam_declaration15211 specparam_declaration_instance15211();
    specparam_declaration15212 specparam_declaration_instance15212();
    specparam_declaration15213 specparam_declaration_instance15213();
    specparam_declaration15214 specparam_declaration_instance15214();
    specparam_declaration15215 specparam_declaration_instance15215();
    specparam_declaration15216 specparam_declaration_instance15216();
    specparam_declaration15217 specparam_declaration_instance15217();
    specparam_declaration15218 specparam_declaration_instance15218();
    specparam_declaration15219 specparam_declaration_instance15219();
    specparam_declaration15220 specparam_declaration_instance15220();
    specparam_declaration15221 specparam_declaration_instance15221();
    specparam_declaration15222 specparam_declaration_instance15222();
    specparam_declaration15223 specparam_declaration_instance15223();
    specparam_declaration15224 specparam_declaration_instance15224();
    specparam_declaration15225 specparam_declaration_instance15225();
    specparam_declaration15226 specparam_declaration_instance15226();
    specparam_declaration15227 specparam_declaration_instance15227();
    specparam_declaration15228 specparam_declaration_instance15228();
    specparam_declaration15229 specparam_declaration_instance15229();
    specparam_declaration15230 specparam_declaration_instance15230();
    specparam_declaration15231 specparam_declaration_instance15231();
    specparam_declaration15232 specparam_declaration_instance15232();
    specparam_declaration15233 specparam_declaration_instance15233();
    specparam_declaration15234 specparam_declaration_instance15234();
    specparam_declaration15235 specparam_declaration_instance15235();
    specparam_declaration15236 specparam_declaration_instance15236();
    specparam_declaration15237 specparam_declaration_instance15237();
    specparam_declaration15238 specparam_declaration_instance15238();
    specparam_declaration15239 specparam_declaration_instance15239();
    specparam_declaration15240 specparam_declaration_instance15240();
    specparam_declaration15241 specparam_declaration_instance15241();
    specparam_declaration15242 specparam_declaration_instance15242();
    specparam_declaration15243 specparam_declaration_instance15243();
    specparam_declaration15244 specparam_declaration_instance15244();
    specparam_declaration15245 specparam_declaration_instance15245();
    specparam_declaration15246 specparam_declaration_instance15246();
    specparam_declaration15247 specparam_declaration_instance15247();
    specparam_declaration15248 specparam_declaration_instance15248();
    specparam_declaration15249 specparam_declaration_instance15249();
    specparam_declaration15250 specparam_declaration_instance15250();
    specparam_declaration15251 specparam_declaration_instance15251();
    specparam_declaration15252 specparam_declaration_instance15252();
    specparam_declaration15253 specparam_declaration_instance15253();
    specparam_declaration15254 specparam_declaration_instance15254();
    specparam_declaration15255 specparam_declaration_instance15255();
    specparam_declaration15256 specparam_declaration_instance15256();
    specparam_declaration15257 specparam_declaration_instance15257();
    specparam_declaration15258 specparam_declaration_instance15258();
    specparam_declaration15259 specparam_declaration_instance15259();
    specparam_declaration15260 specparam_declaration_instance15260();
    specparam_declaration15261 specparam_declaration_instance15261();
    specparam_declaration15262 specparam_declaration_instance15262();
    specparam_declaration15263 specparam_declaration_instance15263();
    specparam_declaration15264 specparam_declaration_instance15264();
    specparam_declaration15265 specparam_declaration_instance15265();
    specparam_declaration15266 specparam_declaration_instance15266();
    specparam_declaration15267 specparam_declaration_instance15267();
    specparam_declaration15268 specparam_declaration_instance15268();
    specparam_declaration15269 specparam_declaration_instance15269();
    specparam_declaration15270 specparam_declaration_instance15270();
    specparam_declaration15271 specparam_declaration_instance15271();
    specparam_declaration15272 specparam_declaration_instance15272();
    specparam_declaration15273 specparam_declaration_instance15273();
    specparam_declaration15274 specparam_declaration_instance15274();
    specparam_declaration15275 specparam_declaration_instance15275();
    specparam_declaration15276 specparam_declaration_instance15276();
    specparam_declaration15277 specparam_declaration_instance15277();
    specparam_declaration15278 specparam_declaration_instance15278();
    specparam_declaration15279 specparam_declaration_instance15279();
    specparam_declaration15280 specparam_declaration_instance15280();
    specparam_declaration15281 specparam_declaration_instance15281();
    specparam_declaration15282 specparam_declaration_instance15282();
    specparam_declaration15283 specparam_declaration_instance15283();
    specparam_declaration15284 specparam_declaration_instance15284();
    specparam_declaration15285 specparam_declaration_instance15285();
    specparam_declaration15286 specparam_declaration_instance15286();
    specparam_declaration15287 specparam_declaration_instance15287();
endmodule
//@
//author : andreib
module specparam_declaration0(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration1(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration16(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration17(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration18(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration19(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration20(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration21(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration22(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration23(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration24(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration25(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration26(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration27(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration28(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration29(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration30(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration31(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration32(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration33(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration34(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration35(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration36(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration37(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration38(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration39(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration40(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration41(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration42(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration43(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration44(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration45(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration46(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration47(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration48(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration49(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration50(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration51(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration52(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration53(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration54(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration55(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration56(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration57(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration58(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration59(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration60(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration61(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration62(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration63(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration64(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration65(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration66(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration67(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration68(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration69(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration70(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration71(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration72(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration73(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration74(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration75(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration76(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration77(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration78(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration79(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration80(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration81(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration82(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration83(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration84(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration85(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration86(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration87(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration88(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration89(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration90(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration91(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration92(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration93(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration94(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration95(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration96(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration97(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration98(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration99(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration100(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration101(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration102(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration103(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration104(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration105(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration106(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration107(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration108(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration109(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration110(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration111(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration112(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration113(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration114(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration115(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration116(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration117(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration118(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration119(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration120(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration121(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration122(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration123(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration124(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration125(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration126(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration127(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration128(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration129(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration130(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration131(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration132(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration133(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration134(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration135(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration136(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration137(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration138(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration139(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration140(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration141(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration142(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration143(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration144(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration145(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration146(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration147(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration148(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration149(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration150(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration151(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration152(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration153(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration154(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration155(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration156(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration157(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration158(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration159(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration160(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration161(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration162(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration163(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration164(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration165(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration166(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration167(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration168(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration169(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration170(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration171(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration172(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration173(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration174(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration175(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration176(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration177(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration178(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration179(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration180(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration181(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration182(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration183(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration184(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration185(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration186(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration187(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration188(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration189(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration190(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration191(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration192(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration193(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration194(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration195(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration196(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration197(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration198(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration199(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration200(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration201(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration202(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration203(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration204(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration205(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration206(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration207(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration208(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration209(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration210(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration211(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration212(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration213(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration214(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration215(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration216(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration217(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration218(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration219(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration220(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration221(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration222(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration223(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration224(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration225(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration226(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration227(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration228(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration229(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration230(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration231(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration232(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration233(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration234(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration235(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration236(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration237(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration238(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration239(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration240(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration241(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration242(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration243(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration244(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration245(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration246(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration247(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration248(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration249(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration250(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration251(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration252(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration253(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration254(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration255(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration256(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration257(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration258(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration259(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration260(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration261(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration262(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration263(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration264(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration265(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration266(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration267(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration268(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration269(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration270(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration271(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration272(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration273(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration274(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration275(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration276(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration277(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration278(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration279(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration280(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration281(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration282(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration283(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration284(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration285(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration286(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration287(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration288(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration289(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration290(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration291(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration292(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration293(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration294(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration295(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration296(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration297(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration298(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration299(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration300(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration301(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration302(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration303(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration304(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration305(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration306(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration307(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration308(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration309(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration310(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration311(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration312(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration313(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration314(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration315(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration316(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration317(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration318(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration319(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration320(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration321(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration322(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration323(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration324(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration325(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration326(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration327(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration328(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration329(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration330(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration331(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration332(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration333(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration334(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration335(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration336(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration337(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration338(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration339(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration340(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration341(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration342(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration343(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration344(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration345(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration346(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration347(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration348(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration349(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration350(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration351(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration352(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration353(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration354(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration355(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration356(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration357(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration358(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration359(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration360(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration361(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration362(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration363(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration364(clk,q);
input clk;
output q;
    specparam test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration365(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration366(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration367(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration368(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration369(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration370(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration371(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration372(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration373(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration374(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration375(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration376(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration377(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration378(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration379(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration380(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration381(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration382(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration383(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration384(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration385(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration386(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration387(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration388(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration389(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration390(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration391(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration392(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration393(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration394(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration395(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration396(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration397(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration398(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration399(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration400(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration401(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration402(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration403(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration404(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration405(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration406(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration407(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration408(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration409(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration410(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration411(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration412(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration413(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration414(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration415(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration416(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration417(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration418(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration419(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration420(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration421(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration422(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration423(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration424(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration425(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration426(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration427(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration428(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration429(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration430(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration431(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration432(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration433(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration434(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration435(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration436(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration437(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration438(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration439(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration440(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration441(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration442(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration443(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration444(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration445(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration446(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration447(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration448(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration449(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration450(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration451(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration452(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration453(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration454(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration455(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration456(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration457(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration458(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration459(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration460(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration461(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration462(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration463(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration464(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration465(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration466(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration467(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration468(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration469(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration470(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration471(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration472(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration473(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration474(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration475(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration476(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration477(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration478(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration479(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration480(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration481(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration482(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration483(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration484(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration485(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration486(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration487(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration488(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration489(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration490(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration491(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration492(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration493(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration494(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration495(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration496(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration497(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration498(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration499(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration500(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration501(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration502(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration503(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration504(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration505(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration506(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration507(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration508(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration509(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration510(clk,q);
input clk;
output q;
    specparam test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration511(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration512(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration513(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration514(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration515(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration516(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration517(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration518(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration519(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration520(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration521(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration522(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration523(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration524(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration525(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration526(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration527(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration528(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration529(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration530(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration531(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration532(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration533(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration534(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration535(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration536(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration537(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration538(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration539(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration540(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration541(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration542(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration543(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration544(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration545(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration546(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration547(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration548(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration549(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration550(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration551(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration552(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration553(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration554(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration555(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration556(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration557(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration558(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration559(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration560(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration561(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration562(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration563(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration564(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration565(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration566(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration567(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration568(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration569(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration570(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration571(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration572(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration573(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration574(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration575(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration576(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration577(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration578(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration579(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration580(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration581(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration582(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration583(clk,q);
input clk;
output q;
    specparam test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration584(clk,q);
input clk;
output q;
    specparam PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration585(clk,q);
input clk;
output q;
    specparam PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration586(clk,q);
input clk;
output q;
    specparam PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration587(clk,q);
input clk;
output q;
    specparam PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration588(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration589(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration590(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration591(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration592(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration593(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration594(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration595(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration596(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration597(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration598(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration599(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration600(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration601(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration602(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration603(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration604(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration605(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration606(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration607(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration608(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration609(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration610(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration611(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration612(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration613(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration614(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration615(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration616(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration617(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration618(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration619(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration620(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration621(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration622(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration623(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration624(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration625(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration626(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration627(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration628(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration629(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration630(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration631(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration632(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration633(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration634(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration635(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration636(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration637(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration638(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration639(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration640(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration641(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration642(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration643(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration644(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration645(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration646(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration647(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration648(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration649(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration650(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration651(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration652(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration653(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration654(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration655(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration656(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration657(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration658(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration659(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration660(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration661(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration662(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration663(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration664(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration665(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration666(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration667(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration668(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration669(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration670(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration671(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration672(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration673(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration674(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration675(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration676(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration677(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration678(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration679(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration680(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration681(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration682(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration683(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration684(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration685(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration686(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration687(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration688(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration689(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration690(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration691(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration692(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration693(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration694(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration695(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration696(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration697(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration698(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration699(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration700(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration701(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration702(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration703(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration704(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration705(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration706(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration707(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration708(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration709(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration710(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration711(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration712(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration713(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration714(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration715(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration716(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration717(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration718(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration719(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration720(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration721(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration722(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration723(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration724(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration725(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration726(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration727(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration728(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration729(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration730(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration731(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration732(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration733(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration734(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration735(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration736(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration737(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration738(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration739(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration740(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration741(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration742(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration743(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration744(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration745(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration746(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration747(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration748(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration749(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration750(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration751(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration752(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration753(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration754(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration755(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration756(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration757(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration758(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration759(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration760(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration761(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration762(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration763(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration764(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration765(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration766(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration767(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration768(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration769(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration770(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration771(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration772(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration773(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration774(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration775(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration776(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration777(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration778(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration779(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration780(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration781(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration782(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration783(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration784(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration785(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration786(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration787(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration788(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration789(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration790(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration791(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration792(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration793(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration794(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration795(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration796(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration797(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration798(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration799(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration800(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration801(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration802(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration803(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration804(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration805(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration806(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration807(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration808(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration809(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration810(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration811(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration812(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration813(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration814(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration815(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration816(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration817(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration818(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration819(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration820(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration821(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration822(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration823(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration824(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration825(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration826(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration827(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration828(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration829(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration830(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration831(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration832(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration833(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration834(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration835(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration836(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration837(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration838(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration839(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration840(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration841(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration842(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration843(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration844(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration845(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration846(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration847(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration848(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration849(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration850(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration851(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration852(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration853(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration854(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration855(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration856(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration857(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration858(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration859(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration860(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration861(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration862(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration863(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration864(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration865(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration866(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration867(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration868(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration869(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration870(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration871(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration872(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration873(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration874(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration875(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration876(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration877(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration878(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration879(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration880(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration881(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration882(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration883(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration884(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration885(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration886(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration887(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration888(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration889(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration890(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration891(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration892(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration893(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration894(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration895(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration896(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration897(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration898(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration899(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration900(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration901(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration902(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration903(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration904(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration905(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration906(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration907(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration908(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration909(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration910(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration911(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration912(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration913(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration914(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration915(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration916(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration917(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration918(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration919(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration920(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration921(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration922(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration923(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration924(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration925(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration926(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration927(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration928(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration929(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration930(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration931(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration932(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration933(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration934(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration935(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration936(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration937(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration938(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration939(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration940(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration941(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration942(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration943(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration944(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration945(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration946(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration947(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration948(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration949(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration950(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration951(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration952(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration953(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration954(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration955(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration956(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration957(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration958(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration959(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration960(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration961(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration962(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration963(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration964(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration965(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration966(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration967(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration968(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration969(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration970(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration971(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration972(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration973(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration974(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration975(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration976(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration977(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration978(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration979(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration980(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration981(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration982(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration983(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration984(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration985(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration986(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration987(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration988(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration989(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration990(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration991(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration992(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration993(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration994(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration995(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration996(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration997(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration998(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration999(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1000(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1001(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1002(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1003(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1004(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1005(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1006(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1007(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1008(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1009(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1010(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1011(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1012(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1013(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1014(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1015(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1016(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1017(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1018(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1019(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1020(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1021(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1022(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1023(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1024(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1025(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1026(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1027(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1028(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1029(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1030(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1031(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1032(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1033(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1034(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1035(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1036(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1037(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1038(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1039(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1040(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1041(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1042(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1043(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1044(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1045(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1046(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1047(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1048(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1049(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1050(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1051(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1052(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1053(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1054(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1055(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1056(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1057(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1058(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1059(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1060(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1061(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1062(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1063(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1064(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1065(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1066(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1067(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1068(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1069(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1070(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1071(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1072(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1073(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1074(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1075(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1076(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1077(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1078(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1079(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1080(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1081(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1082(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1083(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1084(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1085(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1086(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1087(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1088(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1089(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1090(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1091(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1092(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1093(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1094(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1095(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1096(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1097(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1098(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1099(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1100(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1101(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1102(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1103(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1104(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1105(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1106(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1107(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1108(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1109(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1110(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1111(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1112(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1113(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1114(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1115(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1116(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1117(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1118(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1119(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1120(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1121(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1122(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1123(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1124(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1125(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1126(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1127(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1128(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1129(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1130(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1131(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1132(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1133(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1134(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1135(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1136(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1137(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1138(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1139(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1140(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1141(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1142(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1143(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1144(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1145(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1146(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1147(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1148(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1149(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1150(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1151(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1152(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1153(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1154(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1155(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1156(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1157(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1158(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1159(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1160(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1161(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1162(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1163(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1164(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1165(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1166(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1167(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1168(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1169(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1170(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1171(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1172(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration1173(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration1174(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration1175(clk,q);
input clk;
output q;
    specparam [ 2 : 1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration1176(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration1177(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1178(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1179(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1180(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1181(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1182(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1183(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1184(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1185(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1186(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1187(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1188(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1189(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1190(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1191(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1192(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1193(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1194(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1195(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1196(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1197(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1198(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1199(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1200(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1201(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1202(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1203(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1204(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1205(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1206(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1207(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1208(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1209(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1210(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1211(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1212(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1213(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1214(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1215(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1216(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1217(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1218(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1219(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1220(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1221(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1222(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1223(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1224(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1225(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1226(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1227(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1228(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1229(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1230(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1231(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1232(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1233(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1234(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1235(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1236(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1237(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1238(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1239(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1240(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1241(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1242(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1243(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1244(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1245(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1246(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1247(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1248(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1249(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration1250(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1251(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1252(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1253(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1254(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1255(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1256(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1257(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1258(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1259(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1260(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1261(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1262(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1263(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1264(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1265(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1266(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1267(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1268(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1269(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1270(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1271(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1272(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1273(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1274(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1275(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1276(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1277(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1278(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1279(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1280(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1281(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1282(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1283(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1284(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1285(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1286(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1287(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1288(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1289(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1290(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1291(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1292(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1293(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1294(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1295(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1296(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1297(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1298(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1299(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1300(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1301(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1302(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1303(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1304(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1305(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1306(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1307(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1308(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1309(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1310(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1311(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1312(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1313(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1314(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1315(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1316(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1317(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1318(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1319(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1320(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1321(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1322(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration1323(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1324(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1325(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1326(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1327(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1328(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1329(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1330(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1331(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1332(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1333(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1334(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1335(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1336(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1337(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1338(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1339(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1340(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1341(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1342(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1343(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1344(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1345(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1346(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1347(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1348(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1349(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1350(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1351(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1352(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1353(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1354(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1355(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1356(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1357(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1358(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1359(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1360(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1361(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1362(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1363(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1364(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1365(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1366(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1367(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1368(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1369(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1370(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1371(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1372(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1373(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1374(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1375(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1376(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1377(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1378(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1379(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1380(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1381(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1382(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1383(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1384(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1385(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1386(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1387(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1388(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1389(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1390(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1391(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1392(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1393(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1394(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1395(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1396(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1397(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1398(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1399(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1400(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1401(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1402(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1403(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1404(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1405(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1406(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1407(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1408(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1409(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1410(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1411(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1412(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1413(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1414(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1415(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1416(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1417(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1418(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1419(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1420(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1421(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1422(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1423(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1424(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1425(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1426(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1427(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1428(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1429(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1430(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1431(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1432(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1433(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1434(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1435(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1436(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1437(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1438(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1439(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1440(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1441(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1442(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1443(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1444(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1445(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1446(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1447(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1448(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1449(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1450(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1451(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1452(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1453(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1454(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1455(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1456(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1457(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1458(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1459(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1460(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1461(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1462(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1463(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1464(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1465(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1466(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1467(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1468(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration1469(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1470(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1471(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1472(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1473(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1474(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1475(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1476(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1477(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1478(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1479(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1480(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1481(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1482(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1483(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1484(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1485(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1486(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1487(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1488(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1489(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1490(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1491(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1492(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1493(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1494(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1495(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1496(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1497(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1498(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1499(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1500(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1501(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1502(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1503(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1504(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1505(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1506(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1507(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1508(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1509(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1510(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1511(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1512(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1513(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1514(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1515(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1516(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1517(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1518(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1519(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1520(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1521(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1522(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1523(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1524(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1525(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1526(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1527(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1528(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1529(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1530(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1531(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1532(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1533(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1534(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1535(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1536(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1537(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1538(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1539(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1540(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1541(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1542(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1543(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1544(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1545(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1546(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1547(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1548(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1549(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1550(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1551(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1552(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1553(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1554(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1555(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1556(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1557(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1558(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1559(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1560(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1561(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1562(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1563(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1564(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1565(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1566(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1567(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1568(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1569(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1570(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1571(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1572(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1573(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1574(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1575(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1576(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1577(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1578(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1579(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1580(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1581(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1582(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1583(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1584(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1585(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1586(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1587(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1588(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1589(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1590(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1591(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1592(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1593(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1594(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1595(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1596(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1597(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1598(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1599(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1600(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1601(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1602(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1603(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1604(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1605(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1606(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1607(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1608(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1609(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1610(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1611(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1612(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1613(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1614(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1615(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1616(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1617(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1618(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1619(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1620(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1621(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1622(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1623(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1624(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1625(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1626(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1627(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1628(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1629(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1630(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1631(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1632(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1633(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1634(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1635(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1636(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1637(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1638(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1639(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1640(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1641(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1642(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1643(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1644(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1645(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1646(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1647(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1648(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1649(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1650(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1651(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1652(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1653(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1654(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1655(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1656(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1657(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1658(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1659(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1660(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1661(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1662(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1663(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1664(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1665(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1666(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1667(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1668(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1669(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1670(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1671(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1672(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1673(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1674(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1675(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1676(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1677(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1678(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1679(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1680(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1681(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1682(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1683(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1684(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1685(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1686(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1687(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1688(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1689(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1690(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1691(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1692(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1693(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1694(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1695(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1696(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1697(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1698(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1699(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1700(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1701(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1702(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1703(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1704(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1705(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1706(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1707(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1708(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1709(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1710(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1711(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1712(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1713(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1714(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1715(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1716(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1717(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1718(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1719(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1720(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1721(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1722(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1723(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1724(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1725(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1726(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1727(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1728(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1729(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1730(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1731(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1732(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1733(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1734(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1735(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1736(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1737(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1738(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1739(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1740(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1741(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1742(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1743(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1744(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1745(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1746(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1747(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1748(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1749(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1750(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1751(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1752(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1753(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1754(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1755(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1756(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1757(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1758(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1759(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1760(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration1761(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration1762(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration1763(clk,q);
input clk;
output q;
    specparam [ 2 : +1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration1764(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration1765(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1766(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1767(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1768(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1769(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1770(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1771(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1772(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1773(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1774(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1775(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1776(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1777(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1778(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1779(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1780(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1781(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1782(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1783(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1784(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1785(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1786(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1787(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1788(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1789(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1790(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1791(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1792(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1793(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1794(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1795(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1796(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1797(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1798(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1799(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1800(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1801(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1802(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1803(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1804(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1805(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1806(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1807(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1808(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1809(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1810(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1811(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1812(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1813(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1814(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1815(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1816(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1817(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1818(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1819(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1820(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1821(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1822(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1823(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1824(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1825(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1826(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1827(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1828(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1829(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1830(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1831(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1832(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1833(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1834(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1835(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1836(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1837(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration1838(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1839(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1840(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1841(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1842(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1843(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1844(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1845(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1846(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1847(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1848(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1849(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1850(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1851(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1852(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1853(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1854(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1855(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1856(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1857(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1858(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1859(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1860(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1861(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1862(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1863(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1864(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1865(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1866(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1867(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1868(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1869(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1870(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1871(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1872(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1873(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1874(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1875(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1876(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1877(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1878(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1879(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1880(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1881(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1882(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1883(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1884(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1885(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1886(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1887(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1888(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1889(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1890(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1891(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1892(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1893(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1894(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1895(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1896(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1897(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1898(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1899(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1900(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1901(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1902(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1903(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1904(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1905(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1906(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1907(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1908(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1909(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1910(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration1911(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1912(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1913(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1914(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1915(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1916(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1917(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1918(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1919(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1920(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1921(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1922(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1923(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1924(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1925(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1926(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1927(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1928(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1929(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1930(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1931(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1932(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1933(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1934(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1935(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1936(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1937(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1938(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1939(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1940(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1941(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1942(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1943(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1944(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1945(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1946(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1947(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1948(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1949(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1950(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1951(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1952(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1953(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1954(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1955(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1956(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1957(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1958(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1959(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1960(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1961(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1962(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1963(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1964(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1965(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1966(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1967(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1968(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1969(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1970(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1971(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1972(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1973(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1974(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1975(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1976(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1977(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1978(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1979(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1980(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1981(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1982(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1983(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1984(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1985(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1986(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1987(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1988(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1989(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1990(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1991(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration1992(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration1993(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration1994(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration1995(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration1996(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration1997(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration1998(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration1999(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2000(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2001(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2002(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2003(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2004(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2005(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2006(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2007(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2008(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2009(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2010(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2011(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2012(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2013(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2014(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2015(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2016(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2017(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2018(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2019(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2020(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2021(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2022(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2023(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2024(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2025(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2026(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2027(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2028(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2029(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2030(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2031(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2032(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2033(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2034(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2035(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2036(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2037(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2038(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2039(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2040(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2041(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2042(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2043(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2044(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2045(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2046(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2047(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2048(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2049(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2050(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2051(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2052(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2053(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2054(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2055(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2056(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration2057(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2058(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2059(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2060(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2061(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2062(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2063(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2064(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2065(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2066(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2067(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2068(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2069(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2070(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2071(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2072(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2073(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2074(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2075(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2076(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2077(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2078(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2079(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2080(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2081(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2082(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2083(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2084(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2085(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2086(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2087(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2088(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2089(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2090(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2091(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2092(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2093(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2094(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2095(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2096(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2097(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2098(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2099(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2100(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2101(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2102(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2103(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2104(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2105(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2106(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2107(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2108(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2109(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2110(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2111(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2112(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2113(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2114(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2115(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2116(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2117(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2118(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2119(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2120(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2121(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2122(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2123(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2124(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2125(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2126(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2127(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2128(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2129(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2130(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2131(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2132(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2133(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2134(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2135(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2136(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2137(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2138(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2139(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2140(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2141(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2142(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2143(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2144(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2145(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2146(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2147(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2148(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2149(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2150(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2151(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2152(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2153(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2154(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2155(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2156(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2157(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2158(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2159(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2160(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2161(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2162(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2163(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2164(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2165(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2166(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2167(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2168(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2169(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2170(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2171(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2172(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2173(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2174(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2175(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2176(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2177(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2178(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2179(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2180(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2181(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2182(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2183(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2184(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2185(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2186(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2187(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2188(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2189(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2190(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2191(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2192(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2193(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2194(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2195(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2196(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2197(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2198(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2199(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2200(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2201(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2202(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2203(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2204(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2205(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2206(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2207(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2208(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2209(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2210(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2211(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2212(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2213(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2214(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2215(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2216(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2217(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2218(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2219(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2220(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2221(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2222(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2223(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2224(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2225(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2226(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2227(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2228(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2229(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2230(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2231(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2232(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2233(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2234(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2235(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2236(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2237(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2238(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2239(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2240(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2241(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2242(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2243(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2244(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2245(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2246(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2247(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2248(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2249(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2250(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2251(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2252(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2253(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2254(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2255(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2256(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2257(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2258(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2259(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2260(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2261(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2262(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2263(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2264(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2265(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2266(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2267(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2268(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2269(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2270(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2271(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2272(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2273(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2274(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2275(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2276(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2277(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2278(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2279(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2280(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2281(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2282(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2283(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2284(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2285(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2286(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2287(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2288(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2289(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2290(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2291(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2292(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2293(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2294(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2295(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2296(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2297(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2298(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2299(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2300(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2301(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2302(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2303(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2304(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2305(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2306(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2307(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2308(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2309(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2310(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2311(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2312(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2313(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2314(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2315(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2316(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2317(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2318(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2319(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2320(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2321(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2322(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2323(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2324(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2325(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2326(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2327(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2328(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2329(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2330(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2331(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2332(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2333(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2334(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2335(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2336(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2337(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2338(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2339(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2340(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2341(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2342(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2343(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2344(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2345(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2346(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2347(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2348(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration2349(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration2350(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration2351(clk,q);
input clk;
output q;
    specparam [ 2 : 2-1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration2352(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration2353(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2354(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2355(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2356(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2357(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2358(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2359(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2360(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2361(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2362(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2363(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2364(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2365(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2366(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2367(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2368(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2369(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2370(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2371(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2372(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2373(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2374(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2375(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2376(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2377(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2378(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2379(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2380(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2381(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2382(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2383(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2384(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2385(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2386(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2387(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2388(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2389(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2390(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2391(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2392(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2393(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2394(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2395(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2396(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2397(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2398(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2399(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2400(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2401(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2402(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2403(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2404(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2405(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2406(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2407(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2408(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2409(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2410(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2411(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2412(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2413(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2414(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2415(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2416(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2417(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2418(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2419(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2420(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2421(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2422(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2423(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2424(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2425(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration2426(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2427(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2428(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2429(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2430(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2431(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2432(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2433(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2434(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2435(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2436(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2437(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2438(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2439(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2440(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2441(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2442(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2443(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2444(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2445(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2446(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2447(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2448(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2449(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2450(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2451(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2452(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2453(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2454(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2455(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2456(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2457(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2458(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2459(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2460(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2461(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2462(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2463(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2464(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2465(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2466(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2467(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2468(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2469(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2470(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2471(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2472(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2473(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2474(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2475(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2476(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2477(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2478(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2479(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2480(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2481(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2482(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2483(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2484(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2485(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2486(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2487(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2488(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2489(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2490(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2491(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2492(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2493(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2494(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2495(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2496(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2497(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2498(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration2499(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2500(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2501(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2502(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2503(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2504(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2505(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2506(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2507(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2508(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2509(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2510(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2511(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2512(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2513(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2514(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2515(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2516(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2517(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2518(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2519(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2520(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2521(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2522(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2523(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2524(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2525(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2526(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2527(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2528(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2529(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2530(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2531(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2532(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2533(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2534(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2535(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2536(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2537(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2538(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2539(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2540(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2541(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2542(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2543(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2544(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2545(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2546(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2547(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2548(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2549(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2550(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2551(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2552(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2553(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2554(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2555(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2556(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2557(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2558(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2559(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2560(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2561(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2562(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2563(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2564(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2565(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2566(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2567(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2568(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2569(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2570(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2571(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2572(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2573(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2574(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2575(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2576(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2577(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2578(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2579(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2580(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2581(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2582(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2583(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2584(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2585(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2586(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2587(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2588(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2589(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2590(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2591(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2592(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2593(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2594(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2595(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2596(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2597(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2598(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2599(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2600(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2601(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2602(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2603(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2604(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2605(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2606(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2607(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2608(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2609(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2610(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2611(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2612(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2613(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2614(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2615(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2616(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2617(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2618(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2619(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2620(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2621(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2622(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2623(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2624(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2625(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2626(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2627(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2628(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2629(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2630(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2631(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2632(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2633(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2634(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2635(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2636(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2637(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2638(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2639(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2640(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2641(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2642(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2643(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2644(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration2645(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2646(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2647(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2648(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2649(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2650(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2651(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2652(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2653(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2654(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2655(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2656(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2657(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2658(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2659(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2660(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2661(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2662(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2663(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2664(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2665(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2666(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2667(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2668(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2669(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2670(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2671(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2672(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2673(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2674(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2675(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2676(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2677(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2678(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2679(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2680(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2681(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2682(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2683(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2684(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2685(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2686(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2687(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2688(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2689(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2690(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2691(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2692(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2693(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2694(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2695(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2696(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2697(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2698(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2699(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2700(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2701(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2702(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2703(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2704(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2705(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2706(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2707(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2708(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2709(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2710(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2711(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2712(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2713(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2714(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2715(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2716(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2717(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2718(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2719(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2720(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2721(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2722(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2723(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2724(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2725(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2726(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2727(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2728(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2729(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2730(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2731(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2732(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2733(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2734(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2735(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2736(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2737(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2738(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2739(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2740(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2741(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2742(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2743(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2744(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2745(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2746(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2747(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2748(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2749(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2750(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2751(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2752(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2753(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2754(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2755(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2756(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2757(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2758(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2759(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2760(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2761(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2762(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2763(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2764(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2765(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2766(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2767(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2768(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2769(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2770(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2771(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2772(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2773(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2774(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2775(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2776(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2777(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2778(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2779(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2780(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2781(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2782(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2783(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2784(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2785(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2786(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2787(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2788(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2789(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2790(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2791(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2792(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2793(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2794(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2795(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2796(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2797(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2798(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2799(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2800(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2801(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2802(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2803(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2804(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2805(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2806(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2807(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2808(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2809(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2810(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2811(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2812(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2813(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2814(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2815(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2816(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2817(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2818(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2819(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2820(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2821(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2822(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2823(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2824(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2825(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2826(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2827(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2828(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2829(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2830(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2831(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2832(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2833(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2834(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2835(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2836(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2837(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2838(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2839(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2840(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2841(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2842(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2843(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2844(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2845(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2846(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2847(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2848(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2849(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2850(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2851(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2852(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2853(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2854(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2855(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2856(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2857(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2858(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2859(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2860(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2861(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2862(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2863(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2864(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2865(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2866(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2867(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2868(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2869(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2870(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2871(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2872(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2873(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2874(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2875(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2876(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2877(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2878(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2879(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2880(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2881(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2882(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2883(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2884(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2885(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2886(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2887(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2888(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2889(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2890(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2891(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2892(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2893(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2894(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2895(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2896(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2897(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2898(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2899(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2900(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2901(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2902(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2903(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2904(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2905(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2906(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2907(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2908(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2909(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2910(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2911(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2912(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2913(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2914(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2915(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2916(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2917(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2918(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2919(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2920(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2921(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2922(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2923(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2924(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2925(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2926(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2927(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2928(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2929(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2930(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2931(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2932(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2933(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2934(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2935(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2936(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration2937(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration2938(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration2939(clk,q);
input clk;
output q;
    specparam [ 2 : 1?2:3 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration2940(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration2941(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2942(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2943(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2944(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2945(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2946(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2947(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2948(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2949(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2950(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2951(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2952(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2953(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2954(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2955(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2956(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2957(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2958(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2959(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2960(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2961(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2962(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2963(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2964(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2965(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2966(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2967(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2968(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2969(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2970(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2971(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2972(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2973(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2974(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2975(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2976(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2977(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2978(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2979(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2980(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2981(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2982(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2983(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2984(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2985(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2986(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2987(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2988(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2989(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2990(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2991(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration2992(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration2993(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration2994(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration2995(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration2996(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration2997(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration2998(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration2999(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3000(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3001(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3002(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3003(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3004(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3005(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3006(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3007(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3008(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3009(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3010(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3011(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3012(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3013(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration3014(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3015(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3016(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3017(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3018(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3019(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3020(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3021(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3022(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3023(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3024(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3025(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3026(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3027(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3028(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3029(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3030(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3031(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3032(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3033(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3034(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3035(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3036(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3037(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3038(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3039(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3040(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3041(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3042(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3043(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3044(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3045(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3046(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3047(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3048(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3049(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3050(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3051(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3052(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3053(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3054(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3055(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3056(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3057(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3058(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3059(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3060(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3061(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3062(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3063(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3064(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3065(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3066(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3067(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3068(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3069(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3070(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3071(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3072(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3073(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3074(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3075(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3076(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3077(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3078(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3079(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3080(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3081(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3082(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3083(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3084(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3085(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3086(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration3087(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3088(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3089(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3090(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3091(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3092(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3093(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3094(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3095(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3096(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3097(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3098(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3099(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3100(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3101(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3102(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3103(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3104(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3105(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3106(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3107(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3108(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3109(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3110(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3111(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3112(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3113(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3114(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3115(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3116(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3117(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3118(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3119(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3120(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3121(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3122(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3123(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3124(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3125(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3126(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3127(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3128(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3129(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3130(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3131(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3132(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3133(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3134(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3135(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3136(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3137(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3138(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3139(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3140(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3141(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3142(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3143(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3144(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3145(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3146(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3147(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3148(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3149(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3150(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3151(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3152(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3153(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3154(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3155(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3156(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3157(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3158(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3159(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3160(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3161(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3162(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3163(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3164(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3165(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3166(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3167(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3168(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3169(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3170(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3171(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3172(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3173(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3174(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3175(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3176(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3177(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3178(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3179(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3180(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3181(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3182(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3183(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3184(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3185(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3186(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3187(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3188(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3189(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3190(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3191(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3192(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3193(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3194(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3195(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3196(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3197(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3198(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3199(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3200(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3201(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3202(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3203(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3204(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3205(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3206(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3207(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3208(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3209(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3210(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3211(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3212(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3213(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3214(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3215(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3216(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3217(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3218(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3219(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3220(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3221(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3222(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3223(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3224(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3225(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3226(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3227(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3228(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3229(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3230(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3231(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3232(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration3233(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3234(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3235(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3236(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3237(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3238(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3239(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3240(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3241(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3242(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3243(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3244(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3245(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3246(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3247(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3248(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3249(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3250(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3251(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3252(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3253(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3254(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3255(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3256(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3257(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3258(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3259(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3260(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3261(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3262(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3263(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3264(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3265(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3266(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3267(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3268(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3269(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3270(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3271(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3272(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3273(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3274(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3275(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3276(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3277(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3278(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3279(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3280(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3281(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3282(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3283(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3284(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3285(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3286(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3287(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3288(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3289(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3290(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3291(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3292(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3293(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3294(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3295(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3296(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3297(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3298(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3299(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3300(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3301(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3302(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3303(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3304(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3305(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3306(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3307(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3308(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3309(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3310(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3311(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3312(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3313(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3314(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3315(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3316(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3317(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3318(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3319(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3320(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3321(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3322(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3323(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3324(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3325(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3326(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3327(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3328(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3329(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3330(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3331(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3332(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3333(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3334(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3335(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3336(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3337(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3338(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3339(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3340(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3341(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3342(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3343(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3344(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3345(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3346(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3347(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3348(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3349(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3350(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3351(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3352(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3353(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3354(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3355(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3356(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3357(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3358(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3359(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3360(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3361(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3362(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3363(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3364(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3365(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3366(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3367(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3368(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3369(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3370(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3371(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3372(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3373(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3374(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3375(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3376(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3377(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3378(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3379(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3380(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3381(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3382(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3383(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3384(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3385(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3386(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3387(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3388(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3389(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3390(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3391(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3392(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3393(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3394(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3395(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3396(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3397(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3398(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3399(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3400(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3401(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3402(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3403(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3404(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3405(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3406(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3407(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3408(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3409(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3410(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3411(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3412(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3413(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3414(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3415(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3416(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3417(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3418(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3419(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3420(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3421(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3422(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3423(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3424(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3425(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3426(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3427(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3428(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3429(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3430(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3431(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3432(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3433(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3434(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3435(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3436(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3437(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3438(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3439(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3440(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3441(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3442(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3443(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3444(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3445(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3446(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3447(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3448(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3449(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3450(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3451(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3452(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3453(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3454(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3455(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3456(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3457(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3458(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3459(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3460(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3461(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3462(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3463(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3464(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3465(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3466(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3467(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3468(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3469(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3470(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3471(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3472(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3473(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3474(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3475(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3476(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3477(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3478(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3479(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3480(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3481(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3482(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3483(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3484(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3485(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3486(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3487(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3488(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3489(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3490(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3491(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3492(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3493(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3494(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3495(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3496(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3497(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3498(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3499(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3500(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3501(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3502(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3503(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3504(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3505(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3506(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3507(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3508(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3509(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3510(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3511(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3512(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3513(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3514(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3515(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3516(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3517(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3518(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3519(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3520(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3521(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3522(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3523(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3524(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration3525(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration3526(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration3527(clk,q);
input clk;
output q;
    specparam [ 2 : "str" ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration3528(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration3529(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3530(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3531(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3532(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3533(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3534(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3535(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3536(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3537(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3538(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3539(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3540(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3541(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3542(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3543(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3544(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3545(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3546(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3547(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3548(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3549(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3550(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3551(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3552(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3553(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3554(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3555(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3556(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3557(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3558(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3559(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3560(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3561(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3562(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3563(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3564(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3565(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3566(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3567(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3568(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3569(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3570(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3571(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3572(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3573(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3574(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3575(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3576(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3577(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3578(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3579(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3580(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3581(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3582(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3583(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3584(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3585(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3586(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3587(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3588(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3589(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3590(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3591(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3592(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3593(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3594(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3595(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3596(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3597(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3598(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3599(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3600(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3601(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration3602(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3603(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3604(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3605(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3606(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3607(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3608(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3609(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3610(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3611(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3612(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3613(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3614(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3615(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3616(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3617(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3618(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3619(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3620(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3621(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3622(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3623(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3624(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3625(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3626(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3627(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3628(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3629(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3630(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3631(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3632(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3633(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3634(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3635(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3636(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3637(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3638(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3639(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3640(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3641(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3642(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3643(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3644(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3645(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3646(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3647(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3648(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3649(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3650(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3651(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3652(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3653(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3654(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3655(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3656(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3657(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3658(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3659(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3660(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3661(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3662(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3663(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3664(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3665(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3666(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3667(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3668(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3669(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3670(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3671(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3672(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3673(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3674(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration3675(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3676(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3677(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3678(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3679(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3680(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3681(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3682(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3683(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3684(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3685(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3686(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3687(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3688(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3689(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3690(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3691(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3692(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3693(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3694(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3695(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3696(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3697(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3698(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3699(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3700(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3701(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3702(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3703(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3704(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3705(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3706(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3707(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3708(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3709(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3710(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3711(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3712(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3713(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3714(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3715(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3716(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3717(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3718(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3719(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3720(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3721(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3722(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3723(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3724(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3725(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3726(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3727(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3728(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3729(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3730(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3731(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3732(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3733(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3734(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3735(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3736(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3737(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3738(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3739(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3740(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3741(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3742(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3743(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3744(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3745(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3746(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3747(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3748(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3749(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3750(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3751(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3752(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3753(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3754(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3755(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3756(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3757(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3758(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3759(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3760(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3761(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3762(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3763(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3764(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3765(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3766(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3767(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3768(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3769(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3770(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3771(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3772(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3773(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3774(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3775(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3776(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3777(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3778(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3779(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3780(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3781(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3782(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3783(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3784(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3785(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3786(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3787(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3788(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3789(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3790(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3791(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3792(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3793(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3794(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3795(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3796(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3797(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3798(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3799(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3800(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3801(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3802(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3803(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3804(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3805(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3806(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3807(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3808(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3809(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3810(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3811(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3812(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3813(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3814(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3815(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3816(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3817(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3818(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3819(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3820(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration3821(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3822(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3823(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3824(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3825(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3826(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3827(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3828(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3829(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3830(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3831(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3832(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3833(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3834(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3835(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3836(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3837(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3838(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3839(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3840(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3841(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3842(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3843(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3844(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3845(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3846(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3847(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3848(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3849(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3850(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3851(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3852(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3853(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3854(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3855(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3856(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3857(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3858(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3859(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3860(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3861(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3862(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3863(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3864(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3865(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3866(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3867(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3868(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3869(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3870(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3871(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3872(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3873(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3874(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3875(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3876(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3877(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3878(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3879(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3880(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3881(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3882(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3883(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3884(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3885(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3886(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3887(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3888(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3889(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3890(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3891(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3892(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3893(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3894(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3895(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3896(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3897(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3898(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3899(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3900(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3901(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3902(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3903(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3904(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3905(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3906(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3907(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3908(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3909(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3910(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3911(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3912(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3913(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3914(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3915(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3916(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3917(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3918(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3919(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3920(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3921(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3922(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3923(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3924(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3925(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3926(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3927(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3928(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3929(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3930(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3931(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3932(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3933(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3934(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3935(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3936(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3937(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3938(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3939(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3940(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3941(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3942(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3943(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3944(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3945(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3946(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3947(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3948(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3949(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3950(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3951(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3952(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3953(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3954(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3955(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3956(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3957(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3958(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3959(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3960(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3961(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3962(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3963(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3964(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3965(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3966(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3967(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3968(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3969(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3970(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3971(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3972(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3973(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3974(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3975(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3976(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3977(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3978(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3979(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3980(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3981(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3982(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3983(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3984(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3985(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3986(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3987(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3988(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3989(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3990(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3991(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration3992(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration3993(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration3994(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration3995(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration3996(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration3997(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration3998(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration3999(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4000(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4001(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4002(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4003(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4004(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4005(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4006(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4007(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4008(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4009(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4010(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4011(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4012(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4013(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4014(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4015(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4016(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4017(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4018(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4019(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4020(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4021(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4022(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4023(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4024(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4025(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4026(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4027(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4028(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4029(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4030(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4031(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4032(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4033(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4034(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4035(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4036(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4037(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4038(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4039(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4040(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4041(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4042(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4043(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4044(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4045(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4046(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4047(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4048(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4049(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4050(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4051(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4052(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4053(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4054(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4055(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4056(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4057(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4058(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4059(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4060(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4061(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4062(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4063(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4064(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4065(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4066(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4067(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4068(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4069(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4070(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4071(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4072(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4073(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4074(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4075(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4076(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4077(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4078(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4079(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4080(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4081(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4082(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4083(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4084(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4085(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4086(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4087(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4088(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4089(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4090(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4091(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4092(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4093(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4094(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4095(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4096(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4097(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4098(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4099(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4100(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4101(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4102(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4103(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4104(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4105(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4106(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4107(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4108(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4109(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4110(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4111(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4112(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration4113(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration4114(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration4115(clk,q);
input clk;
output q;
    specparam [ +3 : 1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration4116(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration4117(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4118(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4119(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4120(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4121(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4122(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4123(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4124(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4125(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4126(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4127(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4128(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4129(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4130(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4131(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4132(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4133(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4134(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4135(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4136(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4137(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4138(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4139(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4140(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4141(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4142(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4143(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4144(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4145(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4146(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4147(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4148(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4149(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4150(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4151(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4152(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4153(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4154(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4155(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4156(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4157(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4158(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4159(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4160(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4161(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4162(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4163(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4164(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4165(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4166(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4167(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4168(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4169(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4170(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4171(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4172(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4173(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4174(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4175(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4176(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4177(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4178(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4179(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4180(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4181(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4182(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4183(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4184(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4185(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4186(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4187(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4188(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4189(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration4190(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4191(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4192(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4193(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4194(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4195(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4196(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4197(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4198(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4199(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4200(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4201(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4202(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4203(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4204(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4205(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4206(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4207(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4208(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4209(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4210(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4211(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4212(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4213(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4214(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4215(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4216(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4217(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4218(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4219(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4220(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4221(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4222(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4223(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4224(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4225(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4226(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4227(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4228(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4229(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4230(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4231(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4232(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4233(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4234(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4235(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4236(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4237(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4238(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4239(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4240(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4241(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4242(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4243(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4244(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4245(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4246(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4247(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4248(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4249(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4250(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4251(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4252(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4253(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4254(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4255(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4256(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4257(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4258(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4259(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4260(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4261(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4262(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration4263(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4264(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4265(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4266(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4267(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4268(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4269(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4270(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4271(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4272(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4273(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4274(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4275(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4276(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4277(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4278(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4279(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4280(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4281(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4282(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4283(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4284(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4285(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4286(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4287(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4288(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4289(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4290(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4291(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4292(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4293(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4294(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4295(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4296(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4297(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4298(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4299(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4300(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4301(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4302(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4303(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4304(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4305(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4306(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4307(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4308(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4309(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4310(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4311(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4312(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4313(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4314(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4315(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4316(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4317(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4318(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4319(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4320(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4321(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4322(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4323(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4324(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4325(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4326(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4327(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4328(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4329(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4330(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4331(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4332(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4333(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4334(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4335(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4336(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4337(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4338(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4339(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4340(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4341(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4342(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4343(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4344(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4345(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4346(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4347(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4348(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4349(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4350(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4351(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4352(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4353(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4354(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4355(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4356(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4357(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4358(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4359(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4360(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4361(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4362(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4363(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4364(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4365(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4366(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4367(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4368(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4369(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4370(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4371(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4372(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4373(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4374(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4375(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4376(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4377(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4378(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4379(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4380(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4381(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4382(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4383(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4384(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4385(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4386(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4387(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4388(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4389(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4390(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4391(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4392(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4393(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4394(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4395(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4396(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4397(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4398(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4399(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4400(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4401(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4402(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4403(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4404(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4405(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4406(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4407(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4408(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration4409(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4410(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4411(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4412(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4413(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4414(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4415(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4416(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4417(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4418(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4419(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4420(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4421(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4422(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4423(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4424(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4425(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4426(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4427(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4428(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4429(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4430(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4431(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4432(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4433(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4434(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4435(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4436(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4437(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4438(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4439(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4440(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4441(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4442(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4443(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4444(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4445(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4446(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4447(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4448(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4449(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4450(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4451(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4452(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4453(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4454(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4455(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4456(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4457(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4458(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4459(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4460(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4461(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4462(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4463(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4464(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4465(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4466(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4467(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4468(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4469(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4470(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4471(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4472(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4473(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4474(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4475(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4476(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4477(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4478(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4479(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4480(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4481(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4482(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4483(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4484(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4485(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4486(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4487(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4488(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4489(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4490(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4491(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4492(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4493(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4494(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4495(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4496(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4497(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4498(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4499(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4500(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4501(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4502(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4503(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4504(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4505(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4506(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4507(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4508(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4509(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4510(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4511(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4512(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4513(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4514(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4515(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4516(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4517(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4518(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4519(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4520(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4521(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4522(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4523(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4524(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4525(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4526(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4527(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4528(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4529(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4530(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4531(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4532(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4533(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4534(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4535(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4536(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4537(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4538(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4539(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4540(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4541(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4542(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4543(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4544(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4545(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4546(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4547(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4548(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4549(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4550(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4551(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4552(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4553(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4554(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4555(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4556(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4557(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4558(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4559(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4560(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4561(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4562(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4563(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4564(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4565(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4566(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4567(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4568(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4569(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4570(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4571(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4572(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4573(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4574(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4575(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4576(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4577(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4578(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4579(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4580(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4581(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4582(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4583(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4584(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4585(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4586(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4587(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4588(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4589(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4590(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4591(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4592(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4593(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4594(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4595(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4596(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4597(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4598(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4599(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4600(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4601(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4602(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4603(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4604(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4605(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4606(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4607(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4608(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4609(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4610(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4611(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4612(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4613(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4614(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4615(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4616(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4617(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4618(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4619(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4620(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4621(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4622(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4623(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4624(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4625(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4626(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4627(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4628(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4629(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4630(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4631(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4632(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4633(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4634(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4635(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4636(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4637(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4638(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4639(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4640(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4641(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4642(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4643(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4644(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4645(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4646(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4647(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4648(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4649(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4650(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4651(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4652(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4653(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4654(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4655(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4656(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4657(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4658(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4659(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4660(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4661(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4662(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4663(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4664(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4665(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4666(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4667(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4668(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4669(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4670(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4671(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4672(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4673(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4674(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4675(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4676(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4677(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4678(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4679(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4680(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4681(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4682(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4683(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4684(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4685(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4686(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4687(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4688(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4689(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4690(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4691(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4692(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4693(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4694(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4695(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4696(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4697(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4698(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4699(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4700(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration4701(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration4702(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration4703(clk,q);
input clk;
output q;
    specparam [ +3 : +1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration4704(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration4705(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4706(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4707(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4708(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4709(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4710(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4711(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4712(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4713(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4714(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4715(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4716(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4717(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4718(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4719(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4720(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4721(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4722(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4723(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4724(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4725(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4726(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4727(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4728(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4729(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4730(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4731(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4732(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4733(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4734(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4735(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4736(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4737(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4738(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4739(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4740(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4741(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4742(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4743(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4744(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4745(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4746(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4747(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4748(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4749(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4750(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4751(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4752(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4753(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4754(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4755(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4756(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4757(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4758(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4759(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4760(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4761(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4762(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4763(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4764(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4765(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4766(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4767(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4768(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4769(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4770(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4771(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4772(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4773(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4774(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4775(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4776(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4777(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration4778(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4779(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4780(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4781(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4782(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4783(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4784(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4785(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4786(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4787(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4788(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4789(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4790(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4791(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4792(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4793(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4794(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4795(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4796(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4797(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4798(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4799(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4800(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4801(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4802(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4803(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4804(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4805(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4806(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4807(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4808(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4809(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4810(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4811(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4812(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4813(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4814(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4815(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4816(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4817(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4818(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4819(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4820(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4821(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4822(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4823(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4824(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4825(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4826(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4827(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4828(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4829(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4830(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4831(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4832(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4833(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4834(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4835(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4836(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4837(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4838(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4839(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4840(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4841(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4842(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4843(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4844(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4845(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4846(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4847(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4848(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4849(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4850(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration4851(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4852(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4853(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4854(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4855(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4856(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4857(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4858(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4859(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4860(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4861(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4862(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4863(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4864(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4865(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4866(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4867(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4868(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4869(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4870(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4871(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4872(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4873(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4874(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4875(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4876(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4877(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4878(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4879(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4880(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4881(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4882(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4883(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4884(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4885(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4886(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4887(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4888(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4889(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4890(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4891(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4892(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4893(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4894(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4895(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4896(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4897(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4898(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4899(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4900(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4901(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4902(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4903(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4904(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4905(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4906(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4907(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4908(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4909(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4910(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4911(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4912(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4913(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4914(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4915(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4916(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4917(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4918(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4919(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4920(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4921(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4922(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4923(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4924(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4925(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4926(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4927(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4928(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4929(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4930(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4931(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4932(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4933(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4934(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4935(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4936(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4937(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4938(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4939(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4940(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4941(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4942(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4943(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4944(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4945(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4946(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4947(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4948(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4949(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4950(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4951(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4952(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4953(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4954(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4955(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4956(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4957(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4958(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4959(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4960(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4961(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4962(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4963(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4964(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4965(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4966(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4967(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4968(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4969(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4970(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4971(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4972(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4973(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4974(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4975(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4976(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4977(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4978(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4979(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4980(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4981(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4982(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4983(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4984(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4985(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4986(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4987(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4988(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4989(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4990(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration4991(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration4992(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration4993(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration4994(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration4995(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration4996(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration4997(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration4998(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration4999(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5000(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5001(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5002(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5003(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5004(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5005(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5006(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5007(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5008(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5009(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5010(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5011(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5012(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5013(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5014(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5015(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5016(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5017(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5018(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5019(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5020(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5021(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5022(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5023(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5024(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5025(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5026(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5027(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5028(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5029(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5030(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5031(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5032(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5033(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5034(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5035(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5036(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5037(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5038(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5039(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5040(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5041(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5042(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5043(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5044(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5045(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5046(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5047(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5048(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5049(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5050(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5051(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5052(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5053(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5054(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5055(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5056(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5057(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5058(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5059(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5060(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5061(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5062(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5063(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5064(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5065(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5066(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5067(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5068(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5069(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5070(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5071(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5072(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5073(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5074(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5075(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5076(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5077(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5078(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5079(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5080(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5081(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5082(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5083(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5084(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5085(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5086(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5087(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5088(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5089(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5090(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5091(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5092(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5093(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5094(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5095(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5096(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5097(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5098(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5099(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5100(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5101(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5102(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5103(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5104(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5105(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5106(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5107(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5108(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5109(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5110(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5111(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5112(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5113(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5114(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5115(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5116(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5117(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5118(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5119(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5120(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5121(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5122(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5123(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5124(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5125(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5126(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5127(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5128(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5129(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5130(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5131(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5132(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5133(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5134(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5135(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5136(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5137(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5138(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5139(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5140(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5141(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5142(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5143(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5144(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5145(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5146(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5147(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5148(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5149(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5150(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5151(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5152(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5153(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5154(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5155(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5156(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5157(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5158(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5159(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5160(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5161(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5162(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5163(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5164(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5165(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5166(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5167(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5168(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5169(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5170(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5171(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5172(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5173(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5174(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5175(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5176(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5177(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5178(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5179(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5180(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5181(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5182(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5183(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5184(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5185(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5186(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5187(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5188(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5189(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5190(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5191(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5192(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5193(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5194(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5195(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5196(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5197(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5198(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5199(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5200(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5201(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5202(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5203(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5204(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5205(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5206(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5207(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5208(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5209(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5210(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5211(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5212(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5213(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5214(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5215(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5216(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5217(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5218(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5219(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5220(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5221(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5222(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5223(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5224(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5225(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5226(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5227(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5228(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5229(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5230(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5231(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5232(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5233(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5234(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5235(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5236(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5237(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5238(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5239(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5240(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5241(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5242(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5243(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5244(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5245(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5246(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5247(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5248(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5249(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5250(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5251(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5252(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5253(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5254(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5255(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5256(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5257(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5258(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5259(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5260(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5261(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5262(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5263(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5264(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5265(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5266(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5267(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5268(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5269(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5270(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5271(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5272(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5273(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5274(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5275(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5276(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5277(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5278(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5279(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5280(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5281(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5282(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5283(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5284(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5285(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5286(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5287(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5288(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration5289(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration5290(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration5291(clk,q);
input clk;
output q;
    specparam [ +3 : 2-1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration5292(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration5293(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5294(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5295(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5296(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5297(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5298(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5299(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5300(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5301(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5302(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5303(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5304(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5305(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5306(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5307(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5308(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5309(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5310(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5311(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5312(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5313(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5314(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5315(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5316(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5317(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5318(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5319(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5320(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5321(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5322(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5323(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5324(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5325(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5326(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5327(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5328(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5329(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5330(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5331(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5332(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5333(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5334(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5335(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5336(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5337(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5338(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5339(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5340(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5341(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5342(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5343(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5344(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5345(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5346(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5347(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5348(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5349(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5350(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5351(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5352(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5353(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5354(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5355(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5356(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5357(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5358(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5359(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5360(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5361(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5362(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5363(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5364(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5365(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration5366(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5367(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5368(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5369(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5370(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5371(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5372(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5373(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5374(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5375(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5376(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5377(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5378(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5379(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5380(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5381(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5382(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5383(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5384(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5385(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5386(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5387(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5388(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5389(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5390(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5391(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5392(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5393(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5394(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5395(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5396(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5397(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5398(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5399(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5400(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5401(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5402(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5403(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5404(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5405(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5406(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5407(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5408(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5409(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5410(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5411(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5412(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5413(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5414(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5415(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5416(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5417(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5418(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5419(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5420(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5421(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5422(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5423(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5424(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5425(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5426(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5427(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5428(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5429(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5430(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5431(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5432(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5433(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5434(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5435(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5436(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5437(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5438(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration5439(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5440(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5441(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5442(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5443(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5444(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5445(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5446(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5447(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5448(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5449(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5450(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5451(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5452(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5453(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5454(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5455(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5456(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5457(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5458(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5459(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5460(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5461(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5462(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5463(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5464(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5465(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5466(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5467(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5468(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5469(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5470(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5471(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5472(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5473(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5474(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5475(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5476(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5477(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5478(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5479(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5480(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5481(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5482(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5483(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5484(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5485(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5486(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5487(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5488(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5489(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5490(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5491(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5492(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5493(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5494(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5495(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5496(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5497(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5498(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5499(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5500(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5501(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5502(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5503(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5504(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5505(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5506(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5507(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5508(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5509(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5510(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5511(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5512(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5513(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5514(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5515(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5516(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5517(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5518(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5519(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5520(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5521(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5522(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5523(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5524(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5525(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5526(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5527(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5528(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5529(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5530(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5531(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5532(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5533(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5534(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5535(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5536(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5537(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5538(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5539(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5540(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5541(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5542(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5543(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5544(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5545(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5546(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5547(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5548(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5549(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5550(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5551(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5552(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5553(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5554(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5555(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5556(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5557(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5558(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5559(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5560(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5561(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5562(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5563(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5564(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5565(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5566(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5567(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5568(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5569(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5570(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5571(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5572(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5573(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5574(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5575(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5576(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5577(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5578(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5579(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5580(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5581(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5582(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5583(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5584(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration5585(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5586(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5587(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5588(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5589(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5590(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5591(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5592(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5593(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5594(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5595(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5596(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5597(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5598(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5599(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5600(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5601(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5602(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5603(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5604(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5605(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5606(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5607(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5608(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5609(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5610(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5611(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5612(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5613(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5614(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5615(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5616(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5617(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5618(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5619(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5620(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5621(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5622(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5623(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5624(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5625(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5626(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5627(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5628(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5629(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5630(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5631(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5632(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5633(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5634(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5635(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5636(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5637(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5638(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5639(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5640(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5641(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5642(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5643(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5644(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5645(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5646(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5647(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5648(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5649(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5650(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5651(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5652(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5653(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5654(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5655(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5656(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5657(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5658(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5659(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5660(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5661(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5662(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5663(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5664(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5665(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5666(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5667(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5668(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5669(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5670(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5671(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5672(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5673(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5674(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5675(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5676(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5677(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5678(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5679(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5680(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5681(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5682(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5683(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5684(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5685(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5686(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5687(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5688(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5689(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5690(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5691(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5692(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5693(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5694(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5695(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5696(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5697(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5698(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5699(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5700(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5701(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5702(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5703(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5704(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5705(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5706(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5707(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5708(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5709(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5710(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5711(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5712(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5713(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5714(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5715(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5716(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5717(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5718(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5719(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5720(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5721(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5722(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5723(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5724(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5725(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5726(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5727(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5728(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5729(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5730(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5731(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5732(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5733(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5734(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5735(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5736(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5737(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5738(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5739(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5740(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5741(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5742(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5743(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5744(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5745(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5746(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5747(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5748(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5749(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5750(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5751(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5752(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5753(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5754(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5755(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5756(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5757(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5758(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5759(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5760(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5761(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5762(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5763(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5764(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5765(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5766(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5767(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5768(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5769(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5770(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5771(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5772(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5773(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5774(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5775(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5776(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5777(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5778(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5779(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5780(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5781(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5782(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5783(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5784(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5785(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5786(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5787(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5788(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5789(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5790(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5791(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5792(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5793(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5794(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5795(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5796(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5797(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5798(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5799(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5800(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5801(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5802(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5803(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5804(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5805(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5806(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5807(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5808(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5809(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5810(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5811(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5812(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5813(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5814(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5815(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5816(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5817(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5818(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5819(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5820(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5821(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5822(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5823(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5824(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5825(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5826(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5827(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5828(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5829(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5830(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5831(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5832(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5833(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5834(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5835(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5836(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5837(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5838(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5839(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5840(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5841(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5842(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5843(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5844(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5845(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5846(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5847(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5848(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5849(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5850(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5851(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5852(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5853(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5854(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5855(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5856(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5857(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5858(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5859(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5860(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5861(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5862(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5863(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5864(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5865(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5866(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5867(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5868(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5869(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5870(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5871(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5872(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5873(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5874(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5875(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5876(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration5877(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration5878(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration5879(clk,q);
input clk;
output q;
    specparam [ +3 : 1?2:3 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration5880(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration5881(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5882(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5883(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5884(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5885(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5886(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5887(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5888(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5889(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5890(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5891(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5892(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5893(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5894(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5895(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5896(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5897(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5898(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5899(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5900(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5901(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5902(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5903(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5904(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5905(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5906(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5907(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5908(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5909(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5910(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5911(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5912(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5913(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5914(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5915(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5916(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5917(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5918(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5919(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5920(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5921(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5922(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5923(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5924(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5925(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5926(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5927(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5928(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5929(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5930(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5931(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5932(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5933(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5934(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5935(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5936(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5937(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5938(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5939(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5940(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5941(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5942(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5943(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5944(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5945(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5946(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5947(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5948(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5949(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5950(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5951(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5952(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5953(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration5954(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5955(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5956(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5957(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5958(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5959(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5960(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5961(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5962(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5963(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5964(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5965(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5966(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5967(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5968(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5969(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5970(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5971(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5972(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5973(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5974(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5975(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5976(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5977(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5978(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5979(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5980(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5981(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5982(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5983(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5984(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5985(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5986(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5987(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5988(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5989(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5990(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5991(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration5992(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration5993(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration5994(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration5995(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration5996(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration5997(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration5998(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration5999(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6000(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6001(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6002(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6003(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6004(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6005(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6006(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6007(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6008(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6009(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6010(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6011(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6012(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6013(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6014(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6015(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6016(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6017(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6018(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6019(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6020(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6021(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6022(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6023(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6024(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6025(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6026(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration6027(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6028(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6029(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6030(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6031(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6032(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6033(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6034(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6035(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6036(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6037(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6038(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6039(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6040(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6041(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6042(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6043(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6044(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6045(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6046(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6047(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6048(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6049(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6050(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6051(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6052(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6053(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6054(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6055(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6056(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6057(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6058(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6059(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6060(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6061(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6062(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6063(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6064(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6065(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6066(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6067(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6068(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6069(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6070(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6071(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6072(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6073(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6074(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6075(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6076(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6077(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6078(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6079(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6080(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6081(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6082(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6083(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6084(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6085(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6086(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6087(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6088(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6089(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6090(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6091(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6092(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6093(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6094(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6095(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6096(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6097(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6098(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6099(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6100(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6101(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6102(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6103(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6104(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6105(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6106(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6107(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6108(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6109(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6110(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6111(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6112(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6113(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6114(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6115(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6116(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6117(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6118(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6119(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6120(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6121(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6122(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6123(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6124(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6125(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6126(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6127(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6128(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6129(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6130(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6131(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6132(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6133(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6134(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6135(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6136(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6137(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6138(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6139(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6140(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6141(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6142(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6143(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6144(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6145(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6146(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6147(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6148(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6149(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6150(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6151(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6152(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6153(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6154(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6155(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6156(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6157(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6158(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6159(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6160(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6161(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6162(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6163(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6164(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6165(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6166(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6167(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6168(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6169(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6170(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6171(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6172(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration6173(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6174(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6175(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6176(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6177(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6178(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6179(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6180(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6181(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6182(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6183(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6184(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6185(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6186(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6187(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6188(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6189(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6190(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6191(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6192(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6193(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6194(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6195(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6196(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6197(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6198(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6199(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6200(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6201(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6202(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6203(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6204(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6205(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6206(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6207(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6208(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6209(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6210(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6211(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6212(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6213(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6214(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6215(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6216(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6217(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6218(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6219(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6220(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6221(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6222(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6223(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6224(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6225(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6226(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6227(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6228(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6229(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6230(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6231(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6232(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6233(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6234(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6235(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6236(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6237(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6238(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6239(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6240(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6241(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6242(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6243(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6244(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6245(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6246(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6247(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6248(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6249(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6250(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6251(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6252(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6253(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6254(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6255(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6256(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6257(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6258(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6259(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6260(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6261(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6262(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6263(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6264(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6265(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6266(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6267(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6268(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6269(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6270(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6271(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6272(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6273(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6274(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6275(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6276(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6277(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6278(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6279(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6280(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6281(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6282(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6283(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6284(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6285(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6286(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6287(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6288(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6289(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6290(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6291(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6292(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6293(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6294(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6295(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6296(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6297(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6298(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6299(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6300(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6301(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6302(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6303(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6304(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6305(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6306(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6307(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6308(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6309(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6310(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6311(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6312(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6313(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6314(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6315(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6316(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6317(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6318(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6319(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6320(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6321(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6322(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6323(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6324(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6325(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6326(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6327(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6328(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6329(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6330(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6331(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6332(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6333(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6334(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6335(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6336(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6337(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6338(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6339(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6340(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6341(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6342(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6343(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6344(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6345(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6346(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6347(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6348(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6349(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6350(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6351(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6352(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6353(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6354(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6355(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6356(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6357(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6358(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6359(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6360(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6361(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6362(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6363(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6364(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6365(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6366(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6367(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6368(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6369(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6370(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6371(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6372(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6373(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6374(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6375(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6376(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6377(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6378(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6379(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6380(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6381(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6382(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6383(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6384(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6385(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6386(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6387(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6388(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6389(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6390(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6391(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6392(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6393(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6394(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6395(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6396(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6397(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6398(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6399(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6400(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6401(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6402(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6403(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6404(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6405(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6406(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6407(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6408(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6409(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6410(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6411(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6412(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6413(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6414(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6415(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6416(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6417(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6418(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6419(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6420(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6421(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6422(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6423(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6424(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6425(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6426(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6427(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6428(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6429(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6430(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6431(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6432(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6433(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6434(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6435(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6436(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6437(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6438(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6439(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6440(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6441(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6442(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6443(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6444(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6445(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6446(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6447(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6448(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6449(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6450(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6451(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6452(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6453(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6454(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6455(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6456(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6457(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6458(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6459(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6460(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6461(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6462(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6463(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6464(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration6465(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration6466(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration6467(clk,q);
input clk;
output q;
    specparam [ +3 : "str" ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration6468(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration6469(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6470(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6471(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6472(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6473(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6474(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6475(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6476(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6477(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6478(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6479(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6480(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6481(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6482(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6483(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6484(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6485(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6486(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6487(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6488(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6489(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6490(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6491(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6492(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6493(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6494(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6495(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6496(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6497(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6498(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6499(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6500(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6501(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6502(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6503(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6504(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6505(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6506(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6507(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6508(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6509(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6510(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6511(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6512(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6513(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6514(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6515(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6516(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6517(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6518(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6519(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6520(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6521(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6522(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6523(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6524(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6525(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6526(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6527(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6528(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6529(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6530(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6531(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6532(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6533(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6534(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6535(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6536(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6537(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6538(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6539(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6540(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6541(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration6542(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6543(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6544(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6545(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6546(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6547(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6548(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6549(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6550(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6551(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6552(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6553(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6554(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6555(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6556(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6557(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6558(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6559(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6560(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6561(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6562(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6563(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6564(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6565(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6566(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6567(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6568(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6569(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6570(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6571(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6572(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6573(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6574(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6575(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6576(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6577(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6578(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6579(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6580(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6581(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6582(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6583(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6584(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6585(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6586(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6587(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6588(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6589(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6590(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6591(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6592(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6593(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6594(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6595(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6596(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6597(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6598(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6599(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6600(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6601(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6602(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6603(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6604(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6605(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6606(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6607(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6608(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6609(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6610(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6611(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6612(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6613(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6614(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration6615(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6616(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6617(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6618(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6619(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6620(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6621(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6622(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6623(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6624(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6625(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6626(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6627(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6628(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6629(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6630(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6631(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6632(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6633(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6634(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6635(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6636(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6637(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6638(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6639(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6640(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6641(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6642(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6643(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6644(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6645(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6646(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6647(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6648(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6649(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6650(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6651(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6652(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6653(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6654(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6655(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6656(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6657(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6658(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6659(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6660(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6661(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6662(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6663(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6664(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6665(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6666(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6667(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6668(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6669(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6670(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6671(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6672(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6673(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6674(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6675(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6676(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6677(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6678(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6679(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6680(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6681(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6682(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6683(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6684(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6685(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6686(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6687(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6688(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6689(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6690(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6691(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6692(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6693(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6694(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6695(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6696(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6697(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6698(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6699(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6700(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6701(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6702(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6703(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6704(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6705(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6706(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6707(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6708(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6709(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6710(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6711(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6712(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6713(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6714(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6715(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6716(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6717(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6718(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6719(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6720(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6721(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6722(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6723(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6724(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6725(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6726(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6727(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6728(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6729(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6730(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6731(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6732(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6733(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6734(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6735(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6736(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6737(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6738(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6739(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6740(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6741(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6742(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6743(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6744(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6745(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6746(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6747(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6748(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6749(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6750(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6751(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6752(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6753(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6754(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6755(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6756(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6757(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6758(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6759(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6760(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration6761(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6762(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6763(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6764(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6765(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6766(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6767(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6768(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6769(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6770(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6771(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6772(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6773(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6774(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6775(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6776(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6777(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6778(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6779(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6780(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6781(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6782(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6783(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6784(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6785(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6786(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6787(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6788(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6789(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6790(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6791(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6792(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6793(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6794(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6795(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6796(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6797(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6798(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6799(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6800(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6801(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6802(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6803(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6804(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6805(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6806(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6807(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6808(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6809(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6810(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6811(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6812(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6813(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6814(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6815(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6816(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6817(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6818(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6819(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6820(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6821(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6822(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6823(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6824(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6825(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6826(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6827(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6828(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6829(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6830(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6831(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6832(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6833(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6834(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6835(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6836(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6837(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6838(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6839(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6840(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6841(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6842(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6843(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6844(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6845(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6846(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6847(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6848(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6849(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6850(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6851(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6852(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6853(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6854(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6855(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6856(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6857(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6858(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6859(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6860(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6861(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6862(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6863(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6864(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6865(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6866(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6867(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6868(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6869(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6870(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6871(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6872(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6873(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6874(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6875(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6876(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6877(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6878(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6879(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6880(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6881(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6882(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6883(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6884(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6885(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6886(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6887(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6888(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6889(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6890(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6891(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6892(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6893(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6894(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6895(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6896(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6897(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6898(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6899(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6900(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6901(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6902(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6903(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6904(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6905(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6906(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6907(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6908(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6909(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6910(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6911(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6912(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6913(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6914(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6915(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6916(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6917(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6918(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6919(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6920(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6921(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6922(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6923(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6924(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6925(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6926(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6927(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6928(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6929(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6930(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6931(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6932(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6933(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6934(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6935(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6936(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6937(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6938(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6939(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6940(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6941(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6942(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6943(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6944(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6945(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6946(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6947(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6948(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6949(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6950(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6951(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6952(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6953(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6954(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6955(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6956(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6957(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6958(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6959(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6960(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6961(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6962(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6963(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6964(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6965(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6966(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6967(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6968(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6969(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6970(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6971(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6972(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6973(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6974(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6975(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6976(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6977(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6978(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6979(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6980(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6981(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6982(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6983(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6984(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6985(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6986(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6987(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6988(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6989(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6990(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6991(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration6992(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration6993(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration6994(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration6995(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration6996(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration6997(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration6998(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration6999(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7000(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7001(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7002(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7003(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7004(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7005(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7006(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7007(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7008(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7009(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7010(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7011(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7012(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7013(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7014(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7015(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7016(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7017(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7018(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7019(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7020(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7021(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7022(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7023(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7024(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7025(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7026(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7027(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7028(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7029(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7030(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7031(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7032(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7033(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7034(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7035(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7036(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7037(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7038(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7039(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7040(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7041(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7042(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7043(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7044(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7045(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7046(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7047(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7048(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7049(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7050(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7051(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7052(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration7053(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration7054(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration7055(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration7056(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration7057(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7058(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7059(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7060(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7061(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7062(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7063(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7064(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7065(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7066(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7067(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7068(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7069(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7070(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7071(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7072(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7073(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7074(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7075(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7076(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7077(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7078(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7079(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7080(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7081(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7082(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7083(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7084(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7085(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7086(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7087(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7088(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7089(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7090(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7091(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7092(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7093(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7094(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7095(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7096(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7097(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7098(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7099(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7100(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7101(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7102(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7103(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7104(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7105(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7106(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7107(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7108(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7109(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7110(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7111(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7112(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7113(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7114(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7115(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7116(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7117(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7118(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7119(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7120(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7121(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7122(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7123(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7124(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7125(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7126(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7127(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7128(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7129(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration7130(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7131(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7132(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7133(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7134(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7135(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7136(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7137(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7138(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7139(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7140(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7141(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7142(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7143(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7144(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7145(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7146(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7147(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7148(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7149(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7150(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7151(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7152(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7153(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7154(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7155(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7156(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7157(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7158(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7159(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7160(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7161(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7162(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7163(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7164(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7165(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7166(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7167(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7168(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7169(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7170(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7171(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7172(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7173(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7174(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7175(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7176(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7177(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7178(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7179(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7180(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7181(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7182(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7183(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7184(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7185(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7186(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7187(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7188(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7189(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7190(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7191(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7192(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7193(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7194(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7195(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7196(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7197(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7198(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7199(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7200(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7201(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7202(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration7203(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7204(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7205(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7206(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7207(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7208(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7209(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7210(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7211(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7212(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7213(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7214(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7215(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7216(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7217(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7218(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7219(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7220(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7221(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7222(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7223(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7224(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7225(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7226(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7227(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7228(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7229(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7230(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7231(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7232(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7233(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7234(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7235(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7236(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7237(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7238(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7239(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7240(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7241(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7242(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7243(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7244(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7245(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7246(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7247(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7248(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7249(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7250(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7251(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7252(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7253(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7254(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7255(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7256(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7257(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7258(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7259(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7260(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7261(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7262(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7263(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7264(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7265(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7266(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7267(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7268(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7269(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7270(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7271(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7272(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7273(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7274(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7275(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7276(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7277(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7278(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7279(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7280(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7281(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7282(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7283(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7284(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7285(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7286(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7287(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7288(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7289(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7290(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7291(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7292(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7293(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7294(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7295(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7296(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7297(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7298(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7299(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7300(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7301(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7302(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7303(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7304(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7305(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7306(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7307(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7308(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7309(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7310(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7311(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7312(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7313(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7314(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7315(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7316(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7317(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7318(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7319(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7320(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7321(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7322(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7323(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7324(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7325(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7326(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7327(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7328(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7329(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7330(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7331(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7332(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7333(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7334(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7335(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7336(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7337(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7338(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7339(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7340(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7341(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7342(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7343(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7344(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7345(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7346(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7347(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7348(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration7349(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7350(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7351(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7352(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7353(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7354(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7355(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7356(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7357(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7358(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7359(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7360(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7361(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7362(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7363(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7364(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7365(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7366(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7367(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7368(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7369(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7370(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7371(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7372(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7373(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7374(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7375(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7376(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7377(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7378(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7379(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7380(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7381(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7382(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7383(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7384(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7385(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7386(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7387(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7388(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7389(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7390(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7391(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7392(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7393(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7394(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7395(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7396(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7397(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7398(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7399(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7400(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7401(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7402(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7403(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7404(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7405(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7406(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7407(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7408(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7409(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7410(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7411(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7412(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7413(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7414(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7415(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7416(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7417(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7418(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7419(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7420(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7421(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7422(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7423(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7424(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7425(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7426(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7427(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7428(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7429(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7430(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7431(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7432(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7433(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7434(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7435(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7436(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7437(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7438(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7439(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7440(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7441(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7442(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7443(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7444(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7445(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7446(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7447(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7448(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7449(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7450(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7451(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7452(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7453(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7454(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7455(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7456(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7457(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7458(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7459(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7460(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7461(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7462(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7463(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7464(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7465(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7466(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7467(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7468(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7469(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7470(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7471(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7472(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7473(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7474(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7475(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7476(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7477(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7478(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7479(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7480(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7481(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7482(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7483(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7484(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7485(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7486(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7487(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7488(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7489(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7490(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7491(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7492(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7493(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7494(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7495(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7496(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7497(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7498(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7499(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7500(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7501(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7502(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7503(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7504(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7505(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7506(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7507(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7508(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7509(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7510(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7511(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7512(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7513(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7514(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7515(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7516(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7517(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7518(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7519(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7520(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7521(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7522(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7523(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7524(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7525(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7526(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7527(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7528(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7529(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7530(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7531(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7532(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7533(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7534(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7535(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7536(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7537(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7538(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7539(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7540(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7541(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7542(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7543(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7544(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7545(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7546(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7547(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7548(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7549(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7550(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7551(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7552(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7553(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7554(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7555(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7556(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7557(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7558(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7559(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7560(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7561(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7562(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7563(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7564(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7565(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7566(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7567(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7568(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7569(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7570(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7571(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7572(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7573(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7574(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7575(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7576(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7577(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7578(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7579(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7580(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7581(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7582(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7583(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7584(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7585(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7586(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7587(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7588(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7589(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7590(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7591(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7592(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7593(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7594(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7595(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7596(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7597(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7598(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7599(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7600(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7601(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7602(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7603(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7604(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7605(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7606(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7607(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7608(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7609(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7610(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7611(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7612(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7613(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7614(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7615(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7616(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7617(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7618(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7619(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7620(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7621(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7622(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7623(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7624(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7625(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7626(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7627(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7628(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7629(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7630(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7631(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7632(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7633(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7634(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7635(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7636(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7637(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7638(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7639(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7640(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration7641(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration7642(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration7643(clk,q);
input clk;
output q;
    specparam [ 2-1 : +1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration7644(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration7645(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7646(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7647(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7648(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7649(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7650(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7651(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7652(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7653(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7654(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7655(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7656(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7657(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7658(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7659(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7660(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7661(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7662(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7663(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7664(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7665(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7666(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7667(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7668(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7669(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7670(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7671(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7672(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7673(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7674(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7675(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7676(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7677(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7678(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7679(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7680(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7681(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7682(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7683(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7684(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7685(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7686(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7687(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7688(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7689(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7690(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7691(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7692(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7693(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7694(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7695(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7696(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7697(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7698(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7699(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7700(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7701(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7702(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7703(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7704(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7705(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7706(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7707(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7708(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7709(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7710(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7711(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7712(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7713(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7714(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7715(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7716(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7717(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration7718(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7719(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7720(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7721(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7722(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7723(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7724(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7725(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7726(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7727(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7728(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7729(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7730(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7731(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7732(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7733(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7734(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7735(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7736(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7737(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7738(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7739(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7740(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7741(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7742(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7743(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7744(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7745(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7746(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7747(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7748(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7749(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7750(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7751(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7752(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7753(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7754(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7755(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7756(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7757(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7758(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7759(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7760(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7761(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7762(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7763(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7764(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7765(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7766(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7767(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7768(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7769(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7770(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7771(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7772(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7773(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7774(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7775(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7776(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7777(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7778(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7779(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7780(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7781(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7782(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7783(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7784(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7785(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7786(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7787(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7788(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7789(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7790(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration7791(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7792(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7793(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7794(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7795(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7796(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7797(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7798(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7799(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7800(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7801(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7802(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7803(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7804(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7805(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7806(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7807(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7808(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7809(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7810(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7811(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7812(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7813(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7814(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7815(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7816(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7817(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7818(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7819(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7820(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7821(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7822(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7823(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7824(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7825(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7826(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7827(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7828(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7829(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7830(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7831(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7832(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7833(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7834(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7835(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7836(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7837(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7838(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7839(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7840(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7841(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7842(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7843(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7844(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7845(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7846(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7847(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7848(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7849(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7850(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7851(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7852(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7853(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7854(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7855(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7856(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7857(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7858(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7859(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7860(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7861(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7862(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7863(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7864(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7865(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7866(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7867(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7868(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7869(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7870(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7871(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7872(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7873(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7874(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7875(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7876(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7877(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7878(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7879(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7880(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7881(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7882(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7883(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7884(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7885(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7886(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7887(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7888(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7889(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7890(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7891(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7892(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7893(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7894(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7895(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7896(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7897(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7898(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7899(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7900(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7901(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7902(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7903(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7904(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7905(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7906(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7907(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7908(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7909(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7910(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7911(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7912(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7913(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7914(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7915(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7916(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7917(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7918(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7919(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7920(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7921(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7922(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7923(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7924(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7925(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7926(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7927(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7928(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7929(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7930(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7931(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7932(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7933(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7934(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7935(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7936(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration7937(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7938(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7939(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7940(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7941(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7942(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7943(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7944(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7945(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7946(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7947(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7948(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7949(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7950(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7951(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7952(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7953(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7954(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7955(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7956(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7957(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7958(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7959(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7960(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7961(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7962(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7963(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7964(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7965(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7966(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7967(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7968(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7969(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7970(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7971(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7972(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7973(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7974(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7975(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7976(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7977(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7978(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7979(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7980(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7981(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7982(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7983(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7984(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7985(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7986(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7987(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7988(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7989(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7990(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7991(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration7992(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration7993(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration7994(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration7995(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration7996(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration7997(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration7998(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration7999(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8000(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8001(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8002(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8003(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8004(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8005(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8006(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8007(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8008(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8009(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8010(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8011(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8012(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8013(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8014(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8015(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8016(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8017(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8018(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8019(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8020(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8021(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8022(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8023(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8024(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8025(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8026(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8027(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8028(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8029(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8030(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8031(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8032(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8033(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8034(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8035(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8036(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8037(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8038(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8039(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8040(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8041(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8042(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8043(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8044(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8045(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8046(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8047(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8048(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8049(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8050(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8051(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8052(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8053(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8054(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8055(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8056(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8057(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8058(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8059(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8060(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8061(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8062(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8063(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8064(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8065(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8066(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8067(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8068(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8069(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8070(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8071(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8072(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8073(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8074(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8075(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8076(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8077(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8078(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8079(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8080(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8081(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8082(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8083(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8084(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8085(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8086(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8087(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8088(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8089(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8090(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8091(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8092(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8093(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8094(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8095(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8096(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8097(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8098(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8099(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8100(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8101(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8102(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8103(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8104(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8105(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8106(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8107(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8108(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8109(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8110(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8111(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8112(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8113(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8114(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8115(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8116(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8117(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8118(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8119(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8120(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8121(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8122(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8123(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8124(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8125(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8126(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8127(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8128(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8129(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8130(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8131(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8132(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8133(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8134(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8135(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8136(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8137(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8138(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8139(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8140(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8141(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8142(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8143(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8144(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8145(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8146(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8147(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8148(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8149(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8150(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8151(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8152(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8153(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8154(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8155(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8156(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8157(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8158(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8159(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8160(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8161(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8162(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8163(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8164(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8165(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8166(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8167(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8168(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8169(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8170(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8171(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8172(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8173(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8174(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8175(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8176(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8177(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8178(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8179(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8180(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8181(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8182(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8183(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8184(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8185(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8186(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8187(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8188(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8189(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8190(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8191(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8192(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8193(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8194(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8195(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8196(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8197(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8198(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8199(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8200(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8201(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8202(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8203(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8204(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8205(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8206(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8207(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8208(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8209(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8210(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8211(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8212(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8213(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8214(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8215(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8216(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8217(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8218(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8219(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8220(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8221(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8222(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8223(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8224(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8225(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8226(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8227(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8228(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration8229(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration8230(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration8231(clk,q);
input clk;
output q;
    specparam [ 2-1 : 2-1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration8232(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration8233(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8234(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8235(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8236(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8237(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8238(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8239(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8240(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8241(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8242(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8243(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8244(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8245(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8246(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8247(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8248(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8249(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8250(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8251(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8252(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8253(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8254(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8255(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8256(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8257(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8258(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8259(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8260(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8261(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8262(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8263(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8264(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8265(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8266(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8267(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8268(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8269(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8270(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8271(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8272(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8273(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8274(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8275(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8276(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8277(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8278(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8279(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8280(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8281(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8282(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8283(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8284(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8285(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8286(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8287(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8288(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8289(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8290(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8291(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8292(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8293(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8294(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8295(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8296(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8297(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8298(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8299(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8300(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8301(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8302(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8303(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8304(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8305(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration8306(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8307(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8308(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8309(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8310(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8311(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8312(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8313(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8314(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8315(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8316(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8317(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8318(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8319(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8320(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8321(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8322(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8323(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8324(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8325(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8326(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8327(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8328(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8329(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8330(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8331(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8332(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8333(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8334(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8335(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8336(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8337(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8338(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8339(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8340(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8341(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8342(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8343(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8344(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8345(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8346(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8347(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8348(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8349(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8350(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8351(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8352(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8353(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8354(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8355(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8356(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8357(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8358(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8359(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8360(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8361(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8362(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8363(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8364(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8365(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8366(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8367(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8368(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8369(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8370(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8371(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8372(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8373(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8374(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8375(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8376(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8377(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8378(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration8379(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8380(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8381(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8382(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8383(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8384(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8385(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8386(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8387(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8388(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8389(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8390(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8391(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8392(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8393(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8394(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8395(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8396(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8397(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8398(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8399(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8400(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8401(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8402(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8403(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8404(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8405(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8406(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8407(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8408(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8409(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8410(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8411(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8412(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8413(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8414(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8415(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8416(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8417(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8418(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8419(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8420(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8421(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8422(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8423(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8424(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8425(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8426(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8427(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8428(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8429(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8430(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8431(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8432(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8433(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8434(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8435(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8436(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8437(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8438(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8439(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8440(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8441(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8442(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8443(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8444(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8445(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8446(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8447(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8448(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8449(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8450(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8451(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8452(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8453(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8454(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8455(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8456(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8457(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8458(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8459(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8460(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8461(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8462(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8463(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8464(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8465(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8466(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8467(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8468(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8469(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8470(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8471(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8472(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8473(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8474(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8475(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8476(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8477(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8478(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8479(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8480(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8481(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8482(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8483(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8484(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8485(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8486(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8487(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8488(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8489(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8490(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8491(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8492(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8493(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8494(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8495(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8496(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8497(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8498(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8499(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8500(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8501(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8502(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8503(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8504(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8505(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8506(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8507(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8508(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8509(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8510(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8511(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8512(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8513(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8514(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8515(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8516(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8517(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8518(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8519(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8520(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8521(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8522(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8523(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8524(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration8525(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8526(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8527(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8528(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8529(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8530(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8531(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8532(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8533(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8534(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8535(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8536(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8537(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8538(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8539(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8540(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8541(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8542(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8543(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8544(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8545(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8546(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8547(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8548(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8549(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8550(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8551(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8552(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8553(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8554(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8555(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8556(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8557(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8558(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8559(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8560(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8561(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8562(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8563(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8564(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8565(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8566(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8567(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8568(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8569(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8570(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8571(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8572(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8573(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8574(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8575(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8576(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8577(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8578(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8579(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8580(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8581(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8582(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8583(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8584(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8585(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8586(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8587(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8588(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8589(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8590(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8591(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8592(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8593(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8594(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8595(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8596(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8597(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8598(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8599(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8600(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8601(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8602(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8603(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8604(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8605(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8606(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8607(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8608(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8609(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8610(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8611(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8612(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8613(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8614(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8615(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8616(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8617(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8618(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8619(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8620(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8621(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8622(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8623(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8624(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8625(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8626(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8627(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8628(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8629(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8630(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8631(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8632(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8633(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8634(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8635(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8636(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8637(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8638(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8639(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8640(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8641(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8642(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8643(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8644(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8645(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8646(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8647(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8648(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8649(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8650(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8651(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8652(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8653(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8654(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8655(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8656(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8657(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8658(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8659(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8660(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8661(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8662(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8663(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8664(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8665(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8666(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8667(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8668(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8669(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8670(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8671(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8672(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8673(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8674(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8675(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8676(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8677(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8678(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8679(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8680(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8681(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8682(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8683(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8684(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8685(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8686(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8687(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8688(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8689(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8690(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8691(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8692(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8693(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8694(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8695(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8696(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8697(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8698(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8699(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8700(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8701(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8702(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8703(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8704(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8705(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8706(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8707(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8708(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8709(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8710(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8711(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8712(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8713(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8714(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8715(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8716(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8717(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8718(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8719(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8720(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8721(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8722(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8723(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8724(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8725(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8726(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8727(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8728(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8729(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8730(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8731(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8732(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8733(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8734(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8735(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8736(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8737(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8738(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8739(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8740(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8741(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8742(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8743(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8744(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8745(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8746(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8747(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8748(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8749(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8750(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8751(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8752(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8753(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8754(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8755(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8756(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8757(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8758(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8759(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8760(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8761(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8762(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8763(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8764(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8765(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8766(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8767(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8768(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8769(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8770(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8771(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8772(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8773(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8774(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8775(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8776(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8777(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8778(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8779(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8780(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8781(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8782(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8783(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8784(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8785(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8786(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8787(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8788(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8789(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8790(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8791(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8792(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8793(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8794(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8795(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8796(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8797(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8798(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8799(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8800(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8801(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8802(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8803(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8804(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8805(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8806(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8807(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8808(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8809(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8810(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8811(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8812(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8813(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8814(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8815(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8816(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration8817(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration8818(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration8819(clk,q);
input clk;
output q;
    specparam [ 2-1 : 1?2:3 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration8820(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration8821(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8822(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8823(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8824(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8825(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8826(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8827(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8828(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8829(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8830(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8831(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8832(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8833(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8834(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8835(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8836(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8837(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8838(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8839(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8840(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8841(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8842(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8843(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8844(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8845(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8846(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8847(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8848(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8849(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8850(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8851(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8852(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8853(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8854(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8855(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8856(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8857(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8858(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8859(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8860(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8861(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8862(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8863(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8864(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8865(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8866(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8867(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8868(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8869(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8870(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8871(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8872(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8873(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8874(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8875(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8876(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8877(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8878(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8879(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8880(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8881(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8882(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8883(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8884(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8885(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8886(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8887(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8888(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8889(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8890(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8891(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8892(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8893(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration8894(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8895(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8896(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8897(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8898(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8899(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8900(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8901(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8902(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8903(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8904(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8905(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8906(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8907(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8908(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8909(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8910(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8911(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8912(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8913(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8914(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8915(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8916(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8917(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8918(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8919(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8920(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8921(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8922(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8923(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8924(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8925(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8926(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8927(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8928(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8929(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8930(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8931(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8932(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8933(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8934(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8935(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8936(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8937(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8938(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8939(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8940(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8941(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8942(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8943(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8944(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8945(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8946(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8947(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8948(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8949(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8950(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8951(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8952(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8953(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8954(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8955(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8956(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8957(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8958(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8959(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8960(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8961(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8962(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8963(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8964(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8965(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8966(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration8967(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8968(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8969(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8970(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8971(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8972(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8973(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8974(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8975(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8976(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8977(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8978(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8979(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8980(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8981(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8982(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8983(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8984(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8985(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8986(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8987(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8988(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8989(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8990(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8991(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration8992(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration8993(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration8994(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration8995(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration8996(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration8997(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration8998(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration8999(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9000(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9001(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9002(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9003(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9004(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9005(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9006(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9007(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9008(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9009(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9010(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9011(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9012(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9013(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9014(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9015(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9016(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9017(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9018(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9019(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9020(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9021(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9022(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9023(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9024(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9025(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9026(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9027(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9028(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9029(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9030(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9031(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9032(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9033(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9034(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9035(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9036(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9037(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9038(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9039(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9040(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9041(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9042(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9043(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9044(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9045(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9046(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9047(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9048(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9049(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9050(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9051(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9052(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9053(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9054(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9055(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9056(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9057(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9058(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9059(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9060(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9061(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9062(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9063(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9064(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9065(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9066(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9067(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9068(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9069(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9070(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9071(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9072(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9073(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9074(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9075(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9076(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9077(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9078(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9079(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9080(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9081(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9082(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9083(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9084(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9085(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9086(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9087(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9088(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9089(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9090(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9091(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9092(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9093(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9094(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9095(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9096(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9097(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9098(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9099(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9100(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9101(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9102(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9103(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9104(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9105(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9106(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9107(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9108(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9109(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9110(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9111(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9112(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration9113(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9114(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9115(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9116(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9117(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9118(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9119(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9120(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9121(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9122(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9123(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9124(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9125(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9126(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9127(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9128(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9129(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9130(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9131(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9132(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9133(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9134(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9135(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9136(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9137(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9138(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9139(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9140(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9141(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9142(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9143(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9144(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9145(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9146(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9147(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9148(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9149(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9150(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9151(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9152(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9153(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9154(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9155(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9156(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9157(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9158(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9159(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9160(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9161(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9162(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9163(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9164(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9165(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9166(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9167(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9168(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9169(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9170(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9171(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9172(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9173(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9174(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9175(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9176(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9177(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9178(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9179(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9180(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9181(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9182(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9183(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9184(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9185(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9186(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9187(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9188(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9189(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9190(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9191(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9192(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9193(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9194(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9195(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9196(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9197(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9198(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9199(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9200(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9201(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9202(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9203(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9204(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9205(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9206(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9207(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9208(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9209(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9210(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9211(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9212(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9213(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9214(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9215(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9216(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9217(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9218(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9219(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9220(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9221(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9222(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9223(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9224(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9225(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9226(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9227(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9228(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9229(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9230(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9231(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9232(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9233(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9234(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9235(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9236(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9237(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9238(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9239(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9240(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9241(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9242(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9243(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9244(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9245(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9246(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9247(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9248(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9249(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9250(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9251(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9252(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9253(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9254(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9255(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9256(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9257(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9258(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9259(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9260(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9261(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9262(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9263(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9264(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9265(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9266(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9267(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9268(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9269(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9270(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9271(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9272(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9273(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9274(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9275(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9276(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9277(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9278(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9279(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9280(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9281(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9282(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9283(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9284(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9285(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9286(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9287(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9288(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9289(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9290(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9291(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9292(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9293(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9294(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9295(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9296(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9297(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9298(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9299(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9300(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9301(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9302(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9303(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9304(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9305(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9306(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9307(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9308(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9309(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9310(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9311(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9312(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9313(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9314(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9315(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9316(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9317(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9318(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9319(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9320(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9321(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9322(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9323(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9324(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9325(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9326(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9327(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9328(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9329(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9330(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9331(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9332(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9333(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9334(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9335(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9336(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9337(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9338(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9339(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9340(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9341(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9342(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9343(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9344(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9345(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9346(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9347(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9348(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9349(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9350(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9351(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9352(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9353(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9354(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9355(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9356(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9357(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9358(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9359(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9360(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9361(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9362(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9363(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9364(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9365(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9366(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9367(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9368(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9369(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9370(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9371(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9372(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9373(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9374(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9375(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9376(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9377(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9378(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9379(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9380(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9381(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9382(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9383(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9384(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9385(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9386(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9387(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9388(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9389(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9390(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9391(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9392(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9393(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9394(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9395(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9396(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9397(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9398(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9399(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9400(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9401(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9402(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9403(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9404(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration9405(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration9406(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration9407(clk,q);
input clk;
output q;
    specparam [ 2-1 : "str" ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration9408(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration9409(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9410(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9411(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9412(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9413(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9414(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9415(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9416(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9417(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9418(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9419(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9420(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9421(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9422(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9423(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9424(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9425(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9426(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9427(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9428(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9429(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9430(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9431(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9432(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9433(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9434(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9435(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9436(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9437(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9438(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9439(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9440(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9441(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9442(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9443(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9444(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9445(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9446(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9447(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9448(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9449(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9450(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9451(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9452(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9453(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9454(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9455(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9456(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9457(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9458(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9459(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9460(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9461(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9462(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9463(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9464(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9465(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9466(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9467(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9468(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9469(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9470(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9471(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9472(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9473(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9474(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9475(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9476(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9477(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9478(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9479(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9480(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9481(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration9482(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9483(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9484(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9485(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9486(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9487(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9488(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9489(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9490(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9491(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9492(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9493(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9494(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9495(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9496(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9497(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9498(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9499(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9500(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9501(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9502(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9503(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9504(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9505(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9506(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9507(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9508(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9509(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9510(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9511(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9512(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9513(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9514(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9515(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9516(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9517(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9518(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9519(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9520(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9521(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9522(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9523(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9524(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9525(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9526(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9527(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9528(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9529(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9530(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9531(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9532(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9533(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9534(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9535(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9536(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9537(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9538(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9539(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9540(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9541(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9542(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9543(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9544(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9545(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9546(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9547(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9548(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9549(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9550(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9551(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9552(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9553(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9554(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration9555(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9556(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9557(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9558(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9559(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9560(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9561(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9562(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9563(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9564(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9565(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9566(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9567(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9568(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9569(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9570(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9571(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9572(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9573(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9574(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9575(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9576(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9577(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9578(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9579(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9580(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9581(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9582(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9583(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9584(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9585(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9586(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9587(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9588(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9589(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9590(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9591(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9592(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9593(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9594(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9595(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9596(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9597(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9598(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9599(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9600(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9601(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9602(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9603(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9604(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9605(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9606(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9607(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9608(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9609(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9610(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9611(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9612(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9613(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9614(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9615(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9616(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9617(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9618(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9619(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9620(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9621(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9622(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9623(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9624(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9625(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9626(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9627(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9628(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9629(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9630(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9631(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9632(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9633(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9634(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9635(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9636(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9637(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9638(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9639(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9640(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9641(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9642(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9643(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9644(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9645(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9646(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9647(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9648(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9649(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9650(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9651(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9652(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9653(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9654(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9655(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9656(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9657(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9658(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9659(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9660(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9661(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9662(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9663(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9664(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9665(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9666(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9667(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9668(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9669(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9670(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9671(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9672(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9673(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9674(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9675(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9676(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9677(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9678(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9679(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9680(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9681(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9682(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9683(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9684(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9685(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9686(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9687(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9688(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9689(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9690(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9691(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9692(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9693(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9694(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9695(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9696(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9697(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9698(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9699(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9700(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration9701(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9702(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9703(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9704(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9705(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9706(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9707(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9708(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9709(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9710(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9711(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9712(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9713(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9714(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9715(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9716(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9717(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9718(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9719(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9720(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9721(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9722(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9723(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9724(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9725(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9726(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9727(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9728(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9729(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9730(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9731(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9732(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9733(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9734(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9735(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9736(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9737(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9738(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9739(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9740(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9741(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9742(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9743(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9744(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9745(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9746(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9747(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9748(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9749(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9750(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9751(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9752(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9753(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9754(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9755(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9756(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9757(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9758(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9759(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9760(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9761(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9762(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9763(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9764(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9765(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9766(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9767(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9768(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9769(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9770(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9771(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9772(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9773(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9774(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9775(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9776(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9777(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9778(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9779(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9780(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9781(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9782(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9783(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9784(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9785(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9786(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9787(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9788(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9789(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9790(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9791(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9792(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9793(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9794(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9795(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9796(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9797(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9798(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9799(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9800(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9801(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9802(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9803(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9804(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9805(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9806(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9807(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9808(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9809(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9810(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9811(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9812(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9813(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9814(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9815(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9816(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9817(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9818(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9819(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9820(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9821(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9822(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9823(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9824(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9825(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9826(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9827(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9828(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9829(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9830(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9831(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9832(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9833(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9834(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9835(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9836(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9837(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9838(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9839(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9840(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9841(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9842(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9843(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9844(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9845(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9846(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9847(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9848(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9849(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9850(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9851(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9852(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9853(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9854(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9855(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9856(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9857(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9858(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9859(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9860(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9861(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9862(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9863(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9864(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9865(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9866(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9867(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9868(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9869(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9870(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9871(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9872(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9873(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9874(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9875(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9876(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9877(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9878(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9879(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9880(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9881(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9882(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9883(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9884(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9885(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9886(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9887(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9888(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9889(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9890(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9891(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9892(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9893(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9894(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9895(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9896(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9897(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9898(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9899(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9900(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9901(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9902(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9903(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9904(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9905(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9906(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9907(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9908(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9909(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9910(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9911(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9912(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9913(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9914(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9915(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9916(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9917(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9918(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9919(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9920(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9921(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9922(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9923(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9924(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9925(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9926(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9927(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9928(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9929(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9930(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9931(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9932(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9933(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9934(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9935(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9936(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9937(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9938(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9939(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9940(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9941(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9942(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9943(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9944(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9945(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9946(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9947(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9948(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9949(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9950(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9951(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9952(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9953(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9954(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9955(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9956(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9957(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9958(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9959(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9960(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9961(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9962(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9963(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9964(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9965(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9966(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9967(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9968(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9969(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9970(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9971(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9972(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9973(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9974(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9975(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9976(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9977(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9978(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9979(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9980(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9981(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9982(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9983(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9984(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9985(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9986(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration9987(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration9988(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration9989(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration9990(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration9991(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration9992(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration9993(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration9994(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration9995(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration9996(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration9997(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration9998(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration9999(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10000(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10001(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10002(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10003(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10004(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10005(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10006(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10007(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10008(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10009(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10010(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10011(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10012(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10013(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10014(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10015(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10016(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10017(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10018(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10019(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10020(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10021(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10022(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10023(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10024(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10025(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10026(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10027(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10028(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10029(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10030(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10031(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10032(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10033(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10034(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10035(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10036(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10037(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10038(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10039(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10040(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10041(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10042(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10043(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10044(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10045(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10046(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10047(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10048(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10049(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10050(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10051(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10052(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10053(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10054(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10055(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10056(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10057(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10058(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10059(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10060(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10061(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10062(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10063(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10064(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10065(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10066(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10067(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10068(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10069(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration10070(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10071(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10072(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10073(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10074(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10075(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10076(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10077(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10078(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10079(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10080(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10081(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10082(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10083(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10084(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10085(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10086(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10087(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10088(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10089(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10090(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10091(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10092(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10093(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10094(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10095(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10096(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10097(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10098(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10099(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10100(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10101(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10102(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10103(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10104(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10105(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10106(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10107(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10108(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10109(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10110(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10111(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10112(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10113(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10114(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10115(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10116(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10117(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10118(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10119(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10120(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10121(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10122(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10123(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10124(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10125(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10126(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10127(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10128(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10129(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10130(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10131(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10132(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10133(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10134(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10135(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10136(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10137(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10138(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10139(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10140(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10141(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10142(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration10143(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10144(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10145(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10146(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10147(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10148(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10149(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10150(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10151(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10152(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10153(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10154(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10155(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10156(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10157(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10158(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10159(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10160(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10161(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10162(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10163(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10164(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10165(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10166(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10167(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10168(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10169(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10170(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10171(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10172(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10173(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10174(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10175(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10176(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10177(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10178(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10179(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10180(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10181(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10182(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10183(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10184(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10185(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10186(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10187(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10188(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10189(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10190(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10191(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10192(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10193(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10194(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10195(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10196(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10197(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10198(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10199(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10200(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10201(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10202(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10203(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10204(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10205(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10206(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10207(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10208(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10209(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10210(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10211(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10212(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10213(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10214(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10215(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10216(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10217(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10218(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10219(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10220(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10221(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10222(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10223(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10224(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10225(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10226(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10227(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10228(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10229(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10230(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10231(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10232(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10233(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10234(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10235(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10236(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10237(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10238(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10239(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10240(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10241(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10242(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10243(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10244(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10245(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10246(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10247(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10248(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10249(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10250(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10251(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10252(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10253(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10254(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10255(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10256(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10257(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10258(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10259(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10260(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10261(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10262(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10263(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10264(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10265(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10266(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10267(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10268(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10269(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10270(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10271(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10272(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10273(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10274(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10275(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10276(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10277(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10278(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10279(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10280(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10281(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10282(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10283(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10284(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10285(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10286(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10287(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10288(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration10289(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10290(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10291(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10292(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10293(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10294(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10295(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10296(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10297(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10298(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10299(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10300(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10301(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10302(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10303(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10304(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10305(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10306(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10307(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10308(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10309(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10310(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10311(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10312(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10313(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10314(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10315(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10316(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10317(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10318(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10319(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10320(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10321(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10322(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10323(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10324(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10325(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10326(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10327(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10328(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10329(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10330(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10331(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10332(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10333(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10334(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10335(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10336(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10337(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10338(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10339(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10340(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10341(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10342(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10343(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10344(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10345(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10346(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10347(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10348(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10349(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10350(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10351(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10352(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10353(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10354(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10355(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10356(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10357(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10358(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10359(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10360(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10361(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10362(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10363(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10364(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10365(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10366(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10367(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10368(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10369(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10370(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10371(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10372(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10373(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10374(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10375(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10376(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10377(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10378(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10379(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10380(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10381(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10382(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10383(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10384(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10385(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10386(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10387(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10388(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10389(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10390(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10391(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10392(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10393(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10394(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10395(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10396(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10397(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10398(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10399(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10400(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10401(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10402(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10403(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10404(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10405(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10406(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10407(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10408(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10409(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10410(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10411(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10412(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10413(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10414(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10415(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10416(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10417(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10418(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10419(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10420(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10421(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10422(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10423(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10424(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10425(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10426(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10427(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10428(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10429(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10430(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10431(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10432(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10433(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10434(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10435(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10436(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10437(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10438(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10439(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10440(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10441(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10442(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10443(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10444(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10445(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10446(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10447(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10448(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10449(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10450(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10451(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10452(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10453(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10454(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10455(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10456(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10457(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10458(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10459(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10460(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10461(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10462(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10463(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10464(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10465(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10466(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10467(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10468(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10469(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10470(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10471(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10472(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10473(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10474(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10475(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10476(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10477(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10478(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10479(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10480(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10481(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10482(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10483(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10484(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10485(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10486(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10487(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10488(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10489(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10490(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10491(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10492(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10493(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10494(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10495(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10496(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10497(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10498(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10499(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10500(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10501(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10502(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10503(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10504(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10505(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10506(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10507(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10508(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10509(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10510(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10511(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10512(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10513(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10514(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10515(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10516(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10517(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10518(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10519(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10520(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10521(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10522(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10523(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10524(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10525(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10526(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10527(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10528(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10529(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10530(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10531(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10532(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10533(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10534(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10535(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10536(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10537(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10538(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10539(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10540(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10541(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10542(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10543(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10544(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10545(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10546(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10547(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10548(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10549(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10550(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10551(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10552(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10553(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10554(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10555(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10556(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10557(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10558(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10559(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10560(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10561(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10562(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10563(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10564(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10565(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10566(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10567(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10568(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10569(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10570(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10571(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10572(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10573(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10574(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10575(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10576(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10577(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10578(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10579(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10580(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration10581(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration10582(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration10583(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : +1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration10584(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration10585(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10586(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10587(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10588(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10589(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10590(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10591(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10592(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10593(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10594(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10595(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10596(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10597(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10598(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10599(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10600(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10601(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10602(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10603(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10604(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10605(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10606(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10607(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10608(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10609(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10610(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10611(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10612(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10613(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10614(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10615(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10616(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10617(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10618(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10619(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10620(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10621(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10622(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10623(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10624(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10625(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10626(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10627(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10628(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10629(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10630(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10631(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10632(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10633(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10634(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10635(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10636(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10637(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10638(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10639(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10640(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10641(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10642(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10643(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10644(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10645(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10646(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10647(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10648(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10649(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10650(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10651(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10652(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10653(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10654(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10655(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10656(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10657(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration10658(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10659(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10660(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10661(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10662(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10663(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10664(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10665(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10666(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10667(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10668(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10669(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10670(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10671(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10672(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10673(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10674(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10675(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10676(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10677(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10678(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10679(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10680(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10681(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10682(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10683(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10684(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10685(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10686(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10687(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10688(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10689(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10690(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10691(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10692(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10693(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10694(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10695(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10696(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10697(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10698(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10699(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10700(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10701(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10702(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10703(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10704(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10705(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10706(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10707(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10708(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10709(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10710(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10711(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10712(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10713(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10714(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10715(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10716(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10717(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10718(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10719(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10720(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10721(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10722(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10723(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10724(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10725(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10726(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10727(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10728(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10729(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10730(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration10731(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10732(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10733(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10734(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10735(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10736(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10737(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10738(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10739(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10740(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10741(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10742(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10743(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10744(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10745(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10746(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10747(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10748(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10749(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10750(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10751(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10752(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10753(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10754(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10755(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10756(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10757(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10758(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10759(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10760(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10761(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10762(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10763(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10764(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10765(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10766(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10767(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10768(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10769(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10770(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10771(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10772(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10773(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10774(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10775(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10776(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10777(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10778(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10779(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10780(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10781(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10782(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10783(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10784(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10785(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10786(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10787(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10788(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10789(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10790(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10791(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10792(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10793(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10794(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10795(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10796(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10797(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10798(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10799(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10800(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10801(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10802(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10803(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10804(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10805(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10806(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10807(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10808(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10809(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10810(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10811(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10812(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10813(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10814(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10815(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10816(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10817(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10818(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10819(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10820(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10821(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10822(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10823(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10824(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10825(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10826(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10827(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10828(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10829(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10830(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10831(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10832(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10833(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10834(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10835(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10836(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10837(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10838(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10839(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10840(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10841(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10842(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10843(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10844(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10845(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10846(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10847(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10848(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10849(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10850(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10851(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10852(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10853(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10854(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10855(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10856(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10857(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10858(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10859(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10860(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10861(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10862(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10863(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10864(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10865(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10866(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10867(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10868(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10869(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10870(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10871(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10872(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10873(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10874(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10875(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10876(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration10877(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10878(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10879(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10880(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10881(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10882(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10883(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10884(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10885(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10886(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10887(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10888(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10889(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10890(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10891(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10892(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10893(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10894(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10895(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10896(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10897(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10898(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10899(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10900(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10901(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10902(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10903(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10904(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10905(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10906(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10907(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10908(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10909(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10910(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10911(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10912(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10913(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10914(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10915(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10916(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10917(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10918(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10919(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10920(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10921(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10922(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10923(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10924(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10925(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10926(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10927(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10928(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10929(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10930(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10931(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10932(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10933(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10934(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10935(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10936(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10937(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10938(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10939(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10940(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10941(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10942(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10943(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10944(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10945(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10946(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10947(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10948(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10949(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10950(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10951(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10952(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10953(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10954(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10955(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10956(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10957(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10958(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10959(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10960(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10961(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10962(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10963(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10964(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10965(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10966(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10967(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10968(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10969(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10970(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10971(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10972(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10973(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10974(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10975(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10976(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10977(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10978(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10979(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10980(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10981(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10982(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10983(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10984(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10985(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10986(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10987(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10988(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10989(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10990(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10991(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration10992(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration10993(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration10994(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration10995(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration10996(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration10997(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration10998(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration10999(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11000(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11001(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11002(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11003(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11004(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11005(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11006(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11007(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11008(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11009(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11010(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11011(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11012(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11013(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11014(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11015(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11016(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11017(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11018(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11019(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11020(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11021(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11022(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11023(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11024(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11025(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11026(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11027(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11028(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11029(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11030(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11031(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11032(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11033(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11034(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11035(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11036(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11037(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11038(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11039(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11040(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11041(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11042(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11043(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11044(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11045(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11046(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11047(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11048(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11049(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11050(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11051(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11052(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11053(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11054(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11055(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11056(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11057(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11058(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11059(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11060(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11061(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11062(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11063(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11064(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11065(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11066(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11067(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11068(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11069(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11070(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11071(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11072(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11073(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11074(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11075(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11076(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11077(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11078(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11079(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11080(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11081(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11082(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11083(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11084(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11085(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11086(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11087(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11088(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11089(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11090(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11091(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11092(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11093(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11094(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11095(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11096(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11097(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11098(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11099(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11100(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11101(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11102(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11103(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11104(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11105(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11106(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11107(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11108(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11109(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11110(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11111(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11112(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11113(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11114(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11115(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11116(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11117(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11118(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11119(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11120(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11121(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11122(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11123(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11124(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11125(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11126(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11127(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11128(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11129(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11130(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11131(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11132(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11133(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11134(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11135(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11136(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11137(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11138(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11139(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11140(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11141(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11142(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11143(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11144(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11145(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11146(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11147(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11148(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11149(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11150(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11151(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11152(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11153(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11154(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11155(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11156(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11157(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11158(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11159(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11160(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11161(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11162(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11163(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11164(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11165(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11166(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11167(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11168(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration11169(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration11170(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration11171(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 2-1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration11172(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration11173(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11174(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11175(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11176(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11177(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11178(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11179(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11180(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11181(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11182(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11183(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11184(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11185(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11186(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11187(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11188(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11189(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11190(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11191(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11192(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11193(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11194(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11195(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11196(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11197(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11198(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11199(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11200(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11201(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11202(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11203(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11204(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11205(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11206(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11207(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11208(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11209(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11210(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11211(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11212(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11213(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11214(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11215(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11216(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11217(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11218(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11219(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11220(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11221(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11222(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11223(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11224(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11225(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11226(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11227(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11228(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11229(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11230(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11231(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11232(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11233(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11234(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11235(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11236(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11237(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11238(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11239(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11240(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11241(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11242(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11243(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11244(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11245(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration11246(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11247(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11248(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11249(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11250(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11251(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11252(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11253(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11254(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11255(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11256(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11257(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11258(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11259(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11260(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11261(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11262(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11263(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11264(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11265(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11266(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11267(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11268(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11269(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11270(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11271(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11272(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11273(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11274(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11275(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11276(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11277(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11278(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11279(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11280(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11281(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11282(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11283(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11284(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11285(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11286(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11287(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11288(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11289(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11290(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11291(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11292(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11293(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11294(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11295(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11296(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11297(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11298(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11299(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11300(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11301(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11302(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11303(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11304(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11305(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11306(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11307(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11308(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11309(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11310(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11311(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11312(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11313(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11314(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11315(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11316(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11317(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11318(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration11319(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11320(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11321(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11322(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11323(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11324(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11325(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11326(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11327(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11328(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11329(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11330(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11331(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11332(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11333(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11334(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11335(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11336(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11337(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11338(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11339(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11340(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11341(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11342(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11343(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11344(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11345(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11346(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11347(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11348(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11349(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11350(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11351(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11352(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11353(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11354(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11355(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11356(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11357(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11358(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11359(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11360(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11361(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11362(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11363(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11364(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11365(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11366(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11367(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11368(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11369(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11370(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11371(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11372(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11373(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11374(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11375(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11376(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11377(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11378(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11379(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11380(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11381(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11382(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11383(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11384(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11385(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11386(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11387(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11388(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11389(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11390(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11391(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11392(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11393(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11394(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11395(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11396(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11397(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11398(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11399(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11400(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11401(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11402(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11403(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11404(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11405(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11406(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11407(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11408(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11409(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11410(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11411(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11412(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11413(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11414(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11415(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11416(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11417(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11418(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11419(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11420(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11421(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11422(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11423(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11424(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11425(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11426(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11427(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11428(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11429(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11430(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11431(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11432(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11433(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11434(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11435(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11436(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11437(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11438(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11439(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11440(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11441(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11442(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11443(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11444(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11445(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11446(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11447(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11448(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11449(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11450(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11451(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11452(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11453(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11454(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11455(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11456(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11457(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11458(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11459(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11460(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11461(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11462(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11463(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11464(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration11465(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11466(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11467(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11468(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11469(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11470(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11471(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11472(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11473(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11474(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11475(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11476(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11477(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11478(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11479(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11480(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11481(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11482(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11483(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11484(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11485(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11486(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11487(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11488(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11489(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11490(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11491(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11492(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11493(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11494(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11495(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11496(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11497(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11498(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11499(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11500(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11501(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11502(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11503(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11504(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11505(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11506(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11507(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11508(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11509(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11510(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11511(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11512(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11513(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11514(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11515(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11516(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11517(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11518(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11519(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11520(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11521(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11522(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11523(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11524(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11525(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11526(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11527(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11528(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11529(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11530(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11531(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11532(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11533(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11534(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11535(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11536(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11537(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11538(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11539(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11540(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11541(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11542(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11543(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11544(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11545(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11546(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11547(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11548(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11549(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11550(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11551(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11552(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11553(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11554(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11555(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11556(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11557(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11558(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11559(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11560(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11561(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11562(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11563(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11564(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11565(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11566(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11567(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11568(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11569(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11570(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11571(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11572(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11573(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11574(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11575(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11576(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11577(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11578(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11579(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11580(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11581(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11582(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11583(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11584(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11585(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11586(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11587(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11588(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11589(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11590(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11591(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11592(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11593(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11594(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11595(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11596(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11597(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11598(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11599(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11600(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11601(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11602(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11603(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11604(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11605(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11606(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11607(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11608(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11609(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11610(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11611(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11612(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11613(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11614(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11615(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11616(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11617(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11618(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11619(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11620(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11621(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11622(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11623(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11624(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11625(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11626(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11627(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11628(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11629(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11630(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11631(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11632(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11633(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11634(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11635(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11636(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11637(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11638(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11639(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11640(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11641(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11642(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11643(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11644(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11645(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11646(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11647(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11648(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11649(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11650(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11651(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11652(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11653(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11654(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11655(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11656(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11657(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11658(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11659(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11660(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11661(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11662(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11663(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11664(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11665(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11666(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11667(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11668(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11669(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11670(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11671(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11672(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11673(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11674(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11675(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11676(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11677(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11678(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11679(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11680(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11681(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11682(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11683(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11684(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11685(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11686(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11687(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11688(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11689(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11690(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11691(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11692(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11693(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11694(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11695(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11696(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11697(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11698(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11699(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11700(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11701(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11702(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11703(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11704(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11705(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11706(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11707(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11708(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11709(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11710(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11711(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11712(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11713(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11714(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11715(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11716(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11717(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11718(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11719(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11720(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11721(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11722(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11723(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11724(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11725(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11726(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11727(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11728(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11729(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11730(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11731(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11732(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11733(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11734(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11735(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11736(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11737(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11738(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11739(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11740(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11741(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11742(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11743(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11744(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11745(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11746(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11747(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11748(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11749(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11750(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11751(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11752(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11753(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11754(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11755(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11756(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration11757(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration11758(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration11759(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : 1?2:3 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration11760(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration11761(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11762(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11763(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11764(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11765(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11766(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11767(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11768(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11769(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11770(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11771(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11772(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11773(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11774(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11775(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11776(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11777(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11778(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11779(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11780(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11781(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11782(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11783(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11784(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11785(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11786(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11787(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11788(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11789(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11790(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11791(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11792(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11793(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11794(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11795(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11796(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11797(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11798(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11799(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11800(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11801(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11802(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11803(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11804(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11805(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11806(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11807(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11808(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11809(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11810(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11811(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11812(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11813(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11814(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11815(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11816(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11817(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11818(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11819(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11820(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11821(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11822(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11823(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11824(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11825(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11826(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11827(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11828(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11829(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11830(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11831(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11832(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11833(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration11834(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11835(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11836(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11837(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11838(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11839(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11840(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11841(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11842(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11843(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11844(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11845(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11846(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11847(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11848(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11849(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11850(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11851(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11852(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11853(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11854(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11855(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11856(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11857(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11858(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11859(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11860(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11861(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11862(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11863(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11864(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11865(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11866(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11867(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11868(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11869(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11870(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11871(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11872(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11873(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11874(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11875(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11876(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11877(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11878(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11879(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11880(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11881(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11882(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11883(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11884(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11885(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11886(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11887(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11888(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11889(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11890(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11891(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11892(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11893(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11894(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11895(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11896(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11897(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11898(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11899(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11900(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11901(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11902(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11903(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11904(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11905(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11906(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration11907(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11908(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11909(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11910(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11911(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11912(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11913(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11914(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11915(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11916(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11917(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11918(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11919(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11920(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11921(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11922(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11923(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11924(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11925(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11926(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11927(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11928(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11929(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11930(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11931(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11932(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11933(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11934(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11935(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11936(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11937(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11938(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11939(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11940(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11941(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11942(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11943(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11944(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11945(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11946(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11947(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11948(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11949(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11950(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11951(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11952(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11953(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11954(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11955(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11956(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11957(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11958(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11959(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11960(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11961(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11962(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11963(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11964(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11965(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11966(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11967(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11968(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11969(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11970(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11971(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11972(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11973(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11974(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11975(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11976(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11977(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11978(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11979(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11980(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11981(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11982(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11983(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11984(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11985(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11986(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11987(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11988(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11989(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11990(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11991(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration11992(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration11993(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration11994(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration11995(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration11996(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration11997(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration11998(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration11999(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12000(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12001(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12002(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12003(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12004(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12005(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12006(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12007(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12008(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12009(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12010(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12011(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12012(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12013(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12014(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12015(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12016(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12017(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12018(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12019(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12020(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12021(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12022(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12023(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12024(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12025(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12026(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12027(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12028(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12029(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12030(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12031(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12032(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12033(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12034(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12035(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12036(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12037(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12038(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12039(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12040(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12041(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12042(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12043(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12044(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12045(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12046(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12047(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12048(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12049(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12050(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12051(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12052(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration12053(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12054(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12055(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12056(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12057(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12058(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12059(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12060(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12061(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12062(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12063(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12064(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12065(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12066(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12067(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12068(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12069(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12070(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12071(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12072(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12073(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12074(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12075(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12076(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12077(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12078(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12079(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12080(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12081(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12082(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12083(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12084(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12085(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12086(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12087(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12088(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12089(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12090(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12091(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12092(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12093(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12094(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12095(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12096(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12097(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12098(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12099(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12100(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12101(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12102(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12103(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12104(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12105(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12106(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12107(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12108(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12109(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12110(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12111(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12112(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12113(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12114(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12115(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12116(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12117(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12118(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12119(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12120(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12121(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12122(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12123(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12124(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12125(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12126(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12127(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12128(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12129(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12130(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12131(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12132(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12133(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12134(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12135(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12136(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12137(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12138(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12139(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12140(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12141(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12142(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12143(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12144(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12145(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12146(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12147(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12148(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12149(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12150(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12151(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12152(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12153(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12154(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12155(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12156(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12157(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12158(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12159(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12160(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12161(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12162(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12163(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12164(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12165(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12166(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12167(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12168(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12169(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12170(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12171(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12172(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12173(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12174(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12175(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12176(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12177(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12178(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12179(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12180(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12181(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12182(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12183(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12184(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12185(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12186(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12187(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12188(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12189(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12190(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12191(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12192(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12193(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12194(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12195(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12196(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12197(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12198(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12199(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12200(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12201(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12202(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12203(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12204(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12205(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12206(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12207(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12208(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12209(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12210(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12211(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12212(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12213(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12214(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12215(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12216(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12217(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12218(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12219(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12220(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12221(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12222(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12223(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12224(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12225(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12226(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12227(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12228(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12229(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12230(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12231(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12232(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12233(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12234(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12235(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12236(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12237(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12238(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12239(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12240(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12241(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12242(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12243(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12244(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12245(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12246(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12247(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12248(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12249(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12250(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12251(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12252(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12253(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12254(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12255(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12256(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12257(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12258(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12259(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12260(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12261(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12262(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12263(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12264(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12265(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12266(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12267(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12268(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12269(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12270(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12271(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12272(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12273(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12274(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12275(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12276(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12277(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12278(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12279(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12280(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12281(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12282(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12283(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12284(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12285(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12286(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12287(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12288(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12289(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12290(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12291(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12292(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12293(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12294(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12295(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12296(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12297(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12298(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12299(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12300(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12301(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12302(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12303(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12304(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12305(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12306(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12307(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12308(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12309(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12310(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12311(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12312(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12313(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12314(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12315(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12316(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12317(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12318(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12319(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12320(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12321(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12322(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12323(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12324(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12325(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12326(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12327(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12328(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12329(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12330(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12331(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12332(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12333(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12334(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12335(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12336(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12337(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12338(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12339(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12340(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12341(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12342(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12343(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12344(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration12345(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration12346(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration12347(clk,q);
input clk;
output q;
    specparam [ 1?2:3 : "str" ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration12348(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration12349(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12350(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12351(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12352(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12353(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12354(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12355(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12356(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12357(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12358(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12359(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12360(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12361(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12362(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12363(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12364(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12365(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12366(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12367(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12368(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12369(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12370(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12371(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12372(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12373(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12374(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12375(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12376(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12377(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12378(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12379(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12380(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12381(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12382(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12383(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12384(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12385(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12386(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12387(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12388(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12389(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12390(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12391(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12392(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12393(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12394(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12395(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12396(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12397(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12398(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12399(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12400(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12401(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12402(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12403(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12404(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12405(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12406(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12407(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12408(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12409(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12410(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12411(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12412(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12413(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12414(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12415(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12416(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12417(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12418(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12419(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12420(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12421(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration12422(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12423(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12424(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12425(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12426(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12427(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12428(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12429(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12430(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12431(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12432(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12433(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12434(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12435(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12436(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12437(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12438(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12439(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12440(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12441(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12442(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12443(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12444(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12445(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12446(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12447(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12448(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12449(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12450(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12451(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12452(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12453(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12454(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12455(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12456(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12457(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12458(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12459(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12460(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12461(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12462(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12463(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12464(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12465(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12466(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12467(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12468(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12469(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12470(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12471(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12472(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12473(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12474(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12475(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12476(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12477(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12478(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12479(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12480(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12481(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12482(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12483(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12484(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12485(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12486(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12487(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12488(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12489(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12490(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12491(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12492(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12493(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12494(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration12495(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12496(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12497(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12498(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12499(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12500(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12501(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12502(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12503(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12504(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12505(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12506(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12507(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12508(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12509(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12510(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12511(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12512(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12513(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12514(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12515(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12516(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12517(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12518(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12519(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12520(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12521(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12522(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12523(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12524(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12525(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12526(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12527(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12528(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12529(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12530(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12531(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12532(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12533(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12534(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12535(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12536(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12537(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12538(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12539(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12540(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12541(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12542(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12543(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12544(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12545(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12546(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12547(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12548(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12549(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12550(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12551(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12552(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12553(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12554(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12555(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12556(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12557(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12558(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12559(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12560(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12561(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12562(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12563(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12564(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12565(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12566(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12567(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12568(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12569(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12570(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12571(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12572(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12573(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12574(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12575(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12576(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12577(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12578(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12579(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12580(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12581(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12582(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12583(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12584(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12585(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12586(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12587(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12588(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12589(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12590(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12591(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12592(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12593(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12594(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12595(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12596(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12597(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12598(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12599(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12600(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12601(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12602(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12603(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12604(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12605(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12606(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12607(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12608(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12609(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12610(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12611(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12612(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12613(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12614(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12615(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12616(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12617(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12618(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12619(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12620(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12621(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12622(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12623(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12624(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12625(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12626(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12627(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12628(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12629(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12630(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12631(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12632(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12633(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12634(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12635(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12636(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12637(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12638(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12639(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12640(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration12641(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12642(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12643(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12644(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12645(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12646(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12647(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12648(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12649(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12650(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12651(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12652(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12653(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12654(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12655(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12656(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12657(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12658(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12659(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12660(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12661(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12662(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12663(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12664(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12665(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12666(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12667(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12668(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12669(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12670(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12671(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12672(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12673(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12674(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12675(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12676(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12677(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12678(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12679(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12680(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12681(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12682(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12683(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12684(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12685(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12686(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12687(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12688(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12689(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12690(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12691(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12692(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12693(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12694(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12695(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12696(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12697(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12698(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12699(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12700(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12701(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12702(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12703(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12704(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12705(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12706(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12707(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12708(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12709(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12710(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12711(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12712(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12713(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12714(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12715(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12716(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12717(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12718(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12719(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12720(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12721(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12722(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12723(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12724(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12725(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12726(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12727(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12728(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12729(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12730(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12731(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12732(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12733(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12734(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12735(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12736(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12737(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12738(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12739(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12740(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12741(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12742(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12743(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12744(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12745(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12746(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12747(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12748(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12749(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12750(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12751(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12752(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12753(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12754(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12755(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12756(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12757(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12758(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12759(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12760(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12761(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12762(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12763(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12764(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12765(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12766(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12767(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12768(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12769(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12770(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12771(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12772(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12773(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12774(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12775(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12776(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12777(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12778(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12779(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12780(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12781(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12782(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12783(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12784(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12785(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12786(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12787(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12788(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12789(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12790(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12791(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12792(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12793(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12794(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12795(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12796(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12797(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12798(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12799(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12800(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12801(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12802(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12803(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12804(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12805(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12806(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12807(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12808(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12809(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12810(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12811(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12812(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12813(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12814(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12815(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12816(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12817(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12818(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12819(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12820(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12821(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12822(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12823(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12824(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12825(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12826(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12827(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12828(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12829(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12830(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12831(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12832(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12833(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12834(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12835(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12836(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12837(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12838(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12839(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12840(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12841(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12842(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12843(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12844(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12845(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12846(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12847(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12848(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12849(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12850(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12851(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12852(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12853(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12854(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12855(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12856(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12857(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12858(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12859(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12860(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12861(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12862(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12863(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12864(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12865(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12866(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12867(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12868(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12869(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12870(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12871(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12872(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12873(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12874(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12875(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12876(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12877(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12878(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12879(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12880(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12881(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12882(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12883(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12884(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12885(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12886(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12887(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12888(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12889(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12890(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12891(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12892(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12893(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12894(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12895(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12896(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12897(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12898(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12899(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12900(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12901(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12902(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12903(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12904(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12905(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12906(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12907(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12908(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12909(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12910(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12911(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12912(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12913(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12914(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12915(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12916(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12917(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12918(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12919(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12920(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12921(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12922(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12923(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12924(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12925(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12926(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12927(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12928(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12929(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12930(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12931(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12932(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration12933(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration12934(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration12935(clk,q);
input clk;
output q;
    specparam [ "str" : 1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration12936(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration12937(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12938(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12939(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12940(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12941(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12942(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12943(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12944(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12945(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12946(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12947(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12948(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12949(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12950(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12951(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12952(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12953(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12954(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12955(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12956(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12957(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12958(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12959(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12960(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12961(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12962(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12963(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12964(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12965(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12966(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12967(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12968(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12969(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12970(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12971(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12972(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12973(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12974(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12975(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12976(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12977(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12978(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12979(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12980(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12981(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12982(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12983(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12984(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12985(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12986(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12987(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12988(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12989(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12990(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12991(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration12992(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration12993(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration12994(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration12995(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration12996(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration12997(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration12998(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration12999(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13000(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13001(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13002(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13003(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13004(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13005(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13006(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13007(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13008(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13009(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration13010(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13011(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13012(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13013(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13014(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13015(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13016(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13017(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13018(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13019(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13020(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13021(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13022(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13023(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13024(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13025(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13026(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13027(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13028(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13029(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13030(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13031(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13032(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13033(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13034(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13035(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13036(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13037(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13038(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13039(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13040(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13041(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13042(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13043(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13044(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13045(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13046(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13047(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13048(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13049(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13050(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13051(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13052(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13053(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13054(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13055(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13056(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13057(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13058(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13059(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13060(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13061(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13062(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13063(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13064(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13065(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13066(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13067(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13068(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13069(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13070(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13071(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13072(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13073(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13074(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13075(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13076(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13077(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13078(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13079(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13080(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13081(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13082(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration13083(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13084(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13085(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13086(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13087(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13088(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13089(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13090(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13091(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13092(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13093(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13094(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13095(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13096(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13097(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13098(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13099(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13100(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13101(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13102(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13103(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13104(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13105(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13106(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13107(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13108(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13109(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13110(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13111(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13112(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13113(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13114(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13115(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13116(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13117(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13118(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13119(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13120(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13121(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13122(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13123(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13124(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13125(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13126(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13127(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13128(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13129(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13130(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13131(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13132(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13133(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13134(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13135(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13136(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13137(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13138(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13139(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13140(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13141(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13142(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13143(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13144(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13145(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13146(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13147(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13148(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13149(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13150(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13151(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13152(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13153(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13154(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13155(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13156(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13157(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13158(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13159(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13160(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13161(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13162(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13163(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13164(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13165(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13166(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13167(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13168(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13169(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13170(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13171(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13172(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13173(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13174(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13175(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13176(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13177(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13178(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13179(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13180(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13181(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13182(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13183(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13184(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13185(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13186(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13187(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13188(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13189(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13190(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13191(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13192(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13193(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13194(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13195(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13196(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13197(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13198(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13199(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13200(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13201(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13202(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13203(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13204(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13205(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13206(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13207(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13208(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13209(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13210(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13211(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13212(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13213(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13214(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13215(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13216(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13217(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13218(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13219(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13220(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13221(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13222(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13223(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13224(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13225(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13226(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13227(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13228(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration13229(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13230(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13231(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13232(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13233(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13234(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13235(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13236(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13237(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13238(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13239(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13240(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13241(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13242(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13243(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13244(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13245(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13246(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13247(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13248(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13249(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13250(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13251(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13252(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13253(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13254(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13255(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13256(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13257(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13258(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13259(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13260(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13261(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13262(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13263(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13264(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13265(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13266(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13267(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13268(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13269(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13270(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13271(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13272(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13273(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13274(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13275(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13276(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13277(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13278(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13279(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13280(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13281(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13282(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13283(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13284(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13285(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13286(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13287(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13288(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13289(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13290(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13291(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13292(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13293(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13294(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13295(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13296(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13297(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13298(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13299(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13300(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13301(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13302(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13303(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13304(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13305(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13306(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13307(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13308(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13309(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13310(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13311(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13312(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13313(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13314(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13315(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13316(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13317(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13318(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13319(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13320(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13321(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13322(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13323(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13324(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13325(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13326(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13327(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13328(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13329(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13330(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13331(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13332(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13333(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13334(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13335(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13336(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13337(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13338(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13339(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13340(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13341(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13342(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13343(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13344(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13345(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13346(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13347(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13348(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13349(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13350(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13351(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13352(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13353(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13354(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13355(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13356(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13357(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13358(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13359(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13360(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13361(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13362(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13363(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13364(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13365(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13366(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13367(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13368(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13369(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13370(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13371(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13372(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13373(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13374(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13375(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13376(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13377(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13378(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13379(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13380(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13381(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13382(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13383(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13384(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13385(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13386(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13387(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13388(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13389(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13390(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13391(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13392(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13393(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13394(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13395(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13396(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13397(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13398(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13399(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13400(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13401(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13402(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13403(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13404(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13405(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13406(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13407(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13408(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13409(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13410(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13411(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13412(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13413(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13414(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13415(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13416(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13417(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13418(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13419(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13420(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13421(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13422(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13423(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13424(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13425(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13426(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13427(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13428(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13429(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13430(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13431(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13432(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13433(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13434(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13435(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13436(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13437(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13438(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13439(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13440(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13441(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13442(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13443(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13444(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13445(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13446(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13447(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13448(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13449(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13450(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13451(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13452(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13453(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13454(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13455(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13456(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13457(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13458(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13459(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13460(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13461(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13462(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13463(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13464(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13465(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13466(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13467(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13468(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13469(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13470(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13471(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13472(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13473(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13474(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13475(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13476(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13477(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13478(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13479(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13480(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13481(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13482(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13483(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13484(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13485(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13486(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13487(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13488(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13489(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13490(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13491(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13492(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13493(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13494(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13495(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13496(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13497(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13498(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13499(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13500(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13501(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13502(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13503(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13504(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13505(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13506(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13507(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13508(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13509(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13510(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13511(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13512(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13513(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13514(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13515(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13516(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13517(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13518(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13519(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13520(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration13521(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration13522(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration13523(clk,q);
input clk;
output q;
    specparam [ "str" : +1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration13524(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration13525(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13526(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13527(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13528(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13529(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13530(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13531(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13532(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13533(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13534(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13535(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13536(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13537(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13538(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13539(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13540(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13541(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13542(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13543(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13544(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13545(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13546(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13547(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13548(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13549(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13550(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13551(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13552(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13553(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13554(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13555(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13556(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13557(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13558(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13559(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13560(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13561(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13562(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13563(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13564(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13565(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13566(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13567(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13568(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13569(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13570(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13571(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13572(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13573(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13574(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13575(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13576(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13577(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13578(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13579(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13580(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13581(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13582(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13583(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13584(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13585(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13586(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13587(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13588(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13589(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13590(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13591(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13592(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13593(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13594(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13595(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13596(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13597(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration13598(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13599(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13600(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13601(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13602(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13603(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13604(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13605(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13606(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13607(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13608(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13609(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13610(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13611(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13612(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13613(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13614(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13615(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13616(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13617(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13618(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13619(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13620(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13621(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13622(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13623(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13624(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13625(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13626(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13627(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13628(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13629(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13630(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13631(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13632(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13633(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13634(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13635(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13636(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13637(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13638(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13639(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13640(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13641(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13642(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13643(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13644(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13645(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13646(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13647(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13648(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13649(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13650(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13651(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13652(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13653(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13654(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13655(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13656(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13657(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13658(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13659(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13660(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13661(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13662(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13663(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13664(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13665(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13666(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13667(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13668(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13669(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13670(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration13671(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13672(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13673(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13674(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13675(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13676(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13677(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13678(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13679(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13680(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13681(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13682(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13683(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13684(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13685(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13686(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13687(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13688(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13689(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13690(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13691(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13692(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13693(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13694(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13695(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13696(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13697(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13698(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13699(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13700(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13701(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13702(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13703(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13704(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13705(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13706(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13707(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13708(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13709(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13710(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13711(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13712(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13713(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13714(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13715(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13716(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13717(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13718(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13719(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13720(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13721(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13722(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13723(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13724(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13725(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13726(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13727(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13728(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13729(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13730(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13731(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13732(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13733(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13734(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13735(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13736(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13737(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13738(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13739(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13740(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13741(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13742(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13743(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13744(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13745(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13746(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13747(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13748(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13749(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13750(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13751(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13752(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13753(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13754(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13755(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13756(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13757(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13758(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13759(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13760(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13761(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13762(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13763(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13764(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13765(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13766(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13767(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13768(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13769(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13770(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13771(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13772(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13773(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13774(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13775(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13776(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13777(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13778(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13779(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13780(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13781(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13782(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13783(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13784(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13785(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13786(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13787(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13788(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13789(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13790(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13791(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13792(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13793(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13794(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13795(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13796(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13797(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13798(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13799(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13800(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13801(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13802(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13803(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13804(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13805(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13806(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13807(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13808(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13809(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13810(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13811(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13812(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13813(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13814(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13815(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13816(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration13817(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13818(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13819(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13820(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13821(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13822(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13823(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13824(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13825(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13826(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13827(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13828(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13829(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13830(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13831(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13832(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13833(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13834(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13835(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13836(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13837(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13838(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13839(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13840(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13841(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13842(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13843(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13844(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13845(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13846(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13847(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13848(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13849(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13850(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13851(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13852(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13853(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13854(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13855(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13856(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13857(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13858(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13859(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13860(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13861(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13862(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13863(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13864(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13865(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13866(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13867(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13868(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13869(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13870(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13871(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13872(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13873(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13874(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13875(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13876(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13877(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13878(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13879(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13880(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13881(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13882(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13883(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13884(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13885(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13886(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13887(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13888(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13889(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13890(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13891(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13892(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13893(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13894(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13895(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13896(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13897(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13898(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13899(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13900(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13901(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13902(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13903(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13904(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13905(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13906(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13907(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13908(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13909(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13910(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13911(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13912(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13913(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13914(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13915(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13916(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13917(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13918(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13919(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13920(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13921(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13922(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13923(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13924(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13925(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13926(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13927(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13928(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13929(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13930(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13931(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13932(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13933(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13934(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13935(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13936(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13937(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13938(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13939(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13940(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13941(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13942(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13943(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13944(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13945(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13946(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13947(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13948(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13949(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13950(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13951(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13952(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13953(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13954(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13955(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13956(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13957(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13958(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13959(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13960(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13961(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13962(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13963(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13964(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13965(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13966(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13967(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13968(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13969(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13970(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13971(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13972(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13973(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13974(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13975(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13976(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13977(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13978(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13979(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13980(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13981(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13982(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13983(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13984(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13985(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13986(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13987(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13988(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13989(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13990(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13991(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration13992(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration13993(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration13994(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration13995(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration13996(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration13997(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration13998(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration13999(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14000(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14001(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14002(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14003(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14004(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14005(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14006(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14007(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14008(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14009(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14010(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14011(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14012(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14013(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14014(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14015(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14016(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14017(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14018(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14019(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14020(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14021(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14022(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14023(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14024(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14025(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14026(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14027(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14028(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14029(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14030(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14031(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14032(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14033(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14034(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14035(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14036(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14037(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14038(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14039(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14040(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14041(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14042(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14043(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14044(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14045(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14046(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14047(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14048(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14049(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14050(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14051(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14052(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14053(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14054(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14055(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14056(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14057(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14058(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14059(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14060(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14061(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14062(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14063(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14064(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14065(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14066(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14067(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14068(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14069(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14070(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14071(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14072(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14073(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14074(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14075(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14076(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14077(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14078(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14079(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14080(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14081(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14082(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14083(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14084(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14085(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14086(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14087(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14088(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14089(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14090(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14091(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14092(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14093(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14094(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14095(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14096(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14097(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14098(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14099(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14100(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14101(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14102(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14103(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14104(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14105(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14106(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14107(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14108(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration14109(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration14110(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration14111(clk,q);
input clk;
output q;
    specparam [ "str" : 2-1 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration14112(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration14113(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14114(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14115(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14116(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14117(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14118(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14119(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14120(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14121(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14122(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14123(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14124(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14125(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14126(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14127(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14128(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14129(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14130(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14131(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14132(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14133(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14134(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14135(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14136(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14137(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14138(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14139(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14140(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14141(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14142(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14143(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14144(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14145(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14146(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14147(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14148(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14149(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14150(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14151(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14152(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14153(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14154(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14155(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14156(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14157(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14158(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14159(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14160(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14161(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14162(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14163(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14164(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14165(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14166(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14167(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14168(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14169(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14170(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14171(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14172(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14173(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14174(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14175(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14176(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14177(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14178(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14179(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14180(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14181(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14182(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14183(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14184(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14185(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration14186(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14187(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14188(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14189(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14190(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14191(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14192(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14193(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14194(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14195(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14196(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14197(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14198(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14199(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14200(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14201(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14202(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14203(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14204(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14205(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14206(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14207(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14208(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14209(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14210(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14211(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14212(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14213(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14214(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14215(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14216(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14217(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14218(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14219(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14220(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14221(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14222(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14223(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14224(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14225(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14226(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14227(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14228(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14229(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14230(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14231(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14232(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14233(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14234(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14235(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14236(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14237(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14238(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14239(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14240(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14241(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14242(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14243(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14244(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14245(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14246(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14247(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14248(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14249(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14250(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14251(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14252(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14253(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14254(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14255(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14256(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14257(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14258(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration14259(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14260(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14261(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14262(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14263(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14264(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14265(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14266(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14267(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14268(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14269(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14270(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14271(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14272(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14273(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14274(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14275(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14276(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14277(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14278(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14279(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14280(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14281(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14282(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14283(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14284(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14285(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14286(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14287(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14288(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14289(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14290(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14291(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14292(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14293(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14294(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14295(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14296(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14297(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14298(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14299(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14300(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14301(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14302(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14303(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14304(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14305(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14306(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14307(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14308(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14309(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14310(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14311(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14312(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14313(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14314(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14315(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14316(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14317(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14318(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14319(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14320(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14321(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14322(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14323(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14324(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14325(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14326(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14327(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14328(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14329(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14330(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14331(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14332(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14333(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14334(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14335(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14336(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14337(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14338(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14339(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14340(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14341(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14342(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14343(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14344(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14345(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14346(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14347(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14348(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14349(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14350(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14351(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14352(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14353(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14354(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14355(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14356(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14357(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14358(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14359(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14360(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14361(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14362(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14363(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14364(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14365(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14366(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14367(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14368(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14369(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14370(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14371(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14372(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14373(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14374(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14375(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14376(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14377(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14378(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14379(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14380(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14381(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14382(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14383(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14384(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14385(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14386(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14387(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14388(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14389(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14390(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14391(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14392(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14393(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14394(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14395(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14396(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14397(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14398(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14399(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14400(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14401(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14402(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14403(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14404(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration14405(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14406(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14407(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14408(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14409(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14410(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14411(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14412(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14413(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14414(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14415(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14416(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14417(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14418(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14419(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14420(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14421(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14422(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14423(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14424(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14425(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14426(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14427(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14428(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14429(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14430(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14431(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14432(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14433(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14434(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14435(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14436(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14437(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14438(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14439(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14440(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14441(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14442(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14443(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14444(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14445(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14446(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14447(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14448(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14449(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14450(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14451(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14452(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14453(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14454(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14455(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14456(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14457(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14458(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14459(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14460(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14461(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14462(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14463(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14464(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14465(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14466(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14467(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14468(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14469(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14470(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14471(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14472(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14473(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14474(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14475(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14476(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14477(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14478(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14479(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14480(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14481(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14482(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14483(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14484(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14485(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14486(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14487(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14488(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14489(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14490(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14491(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14492(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14493(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14494(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14495(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14496(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14497(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14498(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14499(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14500(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14501(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14502(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14503(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14504(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14505(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14506(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14507(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14508(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14509(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14510(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14511(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14512(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14513(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14514(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14515(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14516(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14517(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14518(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14519(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14520(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14521(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14522(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14523(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14524(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14525(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14526(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14527(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14528(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14529(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14530(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14531(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14532(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14533(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14534(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14535(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14536(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14537(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14538(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14539(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14540(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14541(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14542(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14543(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14544(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14545(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14546(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14547(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14548(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14549(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14550(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14551(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14552(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14553(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14554(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14555(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14556(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14557(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14558(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14559(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14560(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14561(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14562(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14563(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14564(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14565(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14566(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14567(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14568(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14569(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14570(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14571(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14572(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14573(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14574(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14575(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14576(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14577(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14578(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14579(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14580(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14581(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14582(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14583(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14584(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14585(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14586(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14587(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14588(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14589(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14590(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14591(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14592(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14593(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14594(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14595(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14596(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14597(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14598(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14599(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14600(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14601(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14602(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14603(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14604(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14605(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14606(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14607(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14608(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14609(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14610(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14611(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14612(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14613(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14614(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14615(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14616(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14617(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14618(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14619(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14620(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14621(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14622(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14623(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14624(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14625(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14626(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14627(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14628(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14629(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14630(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14631(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14632(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14633(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14634(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14635(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14636(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14637(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14638(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14639(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14640(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14641(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14642(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14643(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14644(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14645(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14646(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14647(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14648(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14649(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14650(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14651(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14652(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14653(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14654(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14655(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14656(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14657(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14658(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14659(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14660(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14661(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14662(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14663(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14664(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14665(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14666(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14667(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14668(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14669(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14670(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14671(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14672(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14673(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14674(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14675(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14676(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14677(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14678(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14679(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14680(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14681(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14682(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14683(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14684(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14685(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14686(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14687(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14688(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14689(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14690(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14691(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14692(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14693(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14694(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14695(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14696(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration14697(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration14698(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration14699(clk,q);
input clk;
output q;
    specparam [ "str" : 1?2:3 ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration14700(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2;
endmodule
//author : andreib
module specparam_declaration14701(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14702(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14703(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14704(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14705(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14706(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14707(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14708(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14709(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14710(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14711(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14712(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14713(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14714(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14715(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14716(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14717(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14718(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14719(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14720(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14721(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14722(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14723(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14724(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14725(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14726(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14727(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14728(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14729(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14730(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14731(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14732(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14733(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14734(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14735(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14736(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14737(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14738(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14739(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14740(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14741(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14742(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14743(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14744(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14745(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14746(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14747(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14748(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14749(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14750(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14751(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14752(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14753(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14754(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14755(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14756(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14757(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14758(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14759(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14760(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14761(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14762(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14763(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14764(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14765(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14766(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14767(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14768(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14769(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14770(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14771(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14772(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14773(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1;
endmodule
//author : andreib
module specparam_declaration14774(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14775(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14776(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14777(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14778(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14779(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14780(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14781(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14782(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14783(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14784(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14785(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14786(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14787(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14788(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14789(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14790(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14791(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14792(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14793(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14794(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14795(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14796(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14797(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14798(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14799(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14800(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14801(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14802(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14803(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14804(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14805(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14806(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14807(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14808(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14809(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14810(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14811(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14812(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14813(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14814(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14815(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14816(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14817(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14818(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14819(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14820(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14821(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14822(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14823(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14824(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14825(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14826(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14827(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14828(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14829(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14830(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14831(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14832(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14833(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14834(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14835(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14836(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14837(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14838(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14839(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14840(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14841(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14842(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14843(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14844(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14845(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14846(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1;
endmodule
//author : andreib
module specparam_declaration14847(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14848(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14849(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14850(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14851(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14852(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14853(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14854(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14855(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14856(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14857(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14858(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14859(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14860(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14861(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14862(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14863(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14864(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14865(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14866(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14867(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14868(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14869(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14870(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14871(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14872(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14873(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14874(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14875(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14876(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14877(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14878(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14879(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14880(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14881(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14882(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14883(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14884(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14885(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14886(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14887(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14888(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14889(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14890(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14891(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14892(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14893(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14894(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14895(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14896(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14897(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14898(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14899(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14900(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14901(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14902(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14903(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14904(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14905(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14906(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14907(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14908(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14909(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14910(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14911(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14912(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14913(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14914(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14915(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14916(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14917(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14918(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 2-1 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14919(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14920(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14921(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14922(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14923(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14924(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14925(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14926(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14927(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14928(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14929(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14930(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14931(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14932(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14933(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14934(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14935(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14936(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14937(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14938(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14939(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14940(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14941(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14942(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14943(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14944(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14945(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14946(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14947(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14948(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14949(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14950(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14951(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14952(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14953(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14954(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14955(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14956(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14957(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14958(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14959(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14960(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14961(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14962(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14963(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14964(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14965(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14966(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14967(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14968(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14969(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14970(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14971(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14972(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14973(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14974(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14975(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14976(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14977(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14978(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14979(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14980(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14981(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14982(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14983(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14984(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14985(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14986(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14987(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14988(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14989(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14990(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration14991(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration14992(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str";
endmodule
//author : andreib
module specparam_declaration14993(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration14994(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration14995(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration14996(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration14997(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration14998(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration14999(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15000(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15001(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15002(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15003(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15004(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15005(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15006(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15007(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15008(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15009(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15010(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15011(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15012(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15013(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15014(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15015(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15016(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15017(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15018(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15019(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15020(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15021(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15022(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15023(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15024(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15025(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15026(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15027(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15028(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15029(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15030(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15031(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15032(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15033(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15034(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15035(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15036(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15037(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15038(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15039(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15040(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15041(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15042(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15043(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15044(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15045(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15046(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15047(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15048(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15049(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15050(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15051(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15052(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15053(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15054(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15055(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15056(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15057(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15058(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15059(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15060(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15061(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15062(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15063(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15064(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = "str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15065(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15066(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15067(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15068(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15069(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15070(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15071(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15072(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15073(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15074(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15075(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15076(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15077(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15078(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15079(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15080(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15081(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15082(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15083(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15084(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15085(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15086(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15087(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15088(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15089(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15090(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15091(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15092(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15093(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15094(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15095(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15096(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15097(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15098(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15099(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15100(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15101(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15102(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15103(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15104(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15105(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15106(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15107(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15108(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15109(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15110(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15111(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15112(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15113(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15114(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15115(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15116(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15117(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15118(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15119(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15120(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15121(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15122(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15123(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15124(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15125(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15126(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15127(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15128(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15129(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15130(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15131(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15132(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15133(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15134(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15135(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15136(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15137(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1:2:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15138(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15139(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15140(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15141(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15142(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15143(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15144(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15145(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15146(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15147(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15148(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15149(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15150(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15151(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15152(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15153(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15154(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15155(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15156(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15157(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15158(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15159(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15160(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15161(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15162(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15163(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15164(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15165(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15166(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15167(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15168(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15169(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15170(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15171(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15172(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15173(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15174(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15175(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15176(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15177(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15178(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15179(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15180(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15181(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15182(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15183(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15184(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15185(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15186(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15187(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15188(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15189(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15190(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15191(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15192(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15193(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15194(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15195(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15196(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15197(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15198(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15199(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15200(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15201(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15202(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15203(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15204(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15205(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15206(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15207(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15208(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15209(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15210(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = +1:2-1:3 , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15211(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15212(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15213(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15214(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15215(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15216(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15217(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15218(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15219(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15220(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15221(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15222(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15223(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15224(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15225(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15226(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15227(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15228(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15229(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15230(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15231(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15232(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15233(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15234(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15235(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15236(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15237(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15238(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15239(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15240(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15241(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15242(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15243(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 2-1 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15244(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15245(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15246(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15247(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15248(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15249(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15250(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15251(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15252(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15253(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15254(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15255(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15256(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15257(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15258(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15259(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = "str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15260(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15261(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15262(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15263(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15264(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15265(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15266(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15267(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1:2:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15268(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15269(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15270(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15271(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15272(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15273(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15274(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15275(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = +1:2-1:3 , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15276(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2;
endmodule
//author : andreib
module specparam_declaration15277(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1;
endmodule
//author : andreib
module specparam_declaration15278(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 2-1;
endmodule
//author : andreib
module specparam_declaration15279(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3;
endmodule
//author : andreib
module specparam_declaration15280(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = "str";
endmodule
//author : andreib
module specparam_declaration15281(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1:2:3;
endmodule
//author : andreib
module specparam_declaration15282(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = +1:2-1:3;
endmodule
//author : andreib
module specparam_declaration15283(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] test_specparam_0 = 1?2:3:+2:"str" , test_specparam_1 = 1?2:3:+2:"str" , test_specparam_2 = 1?2:3:+2:"str";
endmodule
//author : andreib
module specparam_declaration15284(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] PATHPULSE$=( 2 );
endmodule
//author : andreib
module specparam_declaration15285(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] PATHPULSE$=( 2 , 8 );
endmodule
//author : andreib
module specparam_declaration15286(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] PATHPULSE$clk$q= ( 2 );
endmodule
//author : andreib
module specparam_declaration15287(clk,q);
input clk;
output q;
    specparam [ "str" : "str" ] PATHPULSE$clk$q= ( 2 , 8 );
endmodule
