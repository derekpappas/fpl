-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./utop_cslc_generated/code/vhdl/u21.vhd
-- FILE GENERATED ON : Sat Mar 14 19:03:19 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u21\ is
  port(\ifcrc2_reset\ : in csl_bit;
       \ifcrc2_clock\ : in csl_bit;
       \pin1\ : in csl_bit_vector(10#8# - 10#1# downto 10#0#);
       \pin2\ : in csl_bit_vector(10#8# - 10#1# downto 10#0#);
       \pout\ : out csl_bit_vector(10#36# - 10#1# downto 10#0#));
begin
end entity;

architecture \u21_logic\ of \u21\ is
begin
end architecture;

