-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./msi_rx_cslc_generated/code/vhdl/ddr_buf_ctrl.vhd
-- FILE GENERATED ON : Tue Jun 17 01:23:46 2008
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity \ddr_buf_ctrl\ is
  port(\lbdummy2\ : in std_logic;
       \dc_dbcdummy5\ : in std_logic);
begin
end entity;

architecture \ddr_buf_ctrl_logic\ of \ddr_buf_ctrl\ is
end architecture;

