// Test type: always statement - loop_statement - 1 attribute instance
// Vparser rule name:
// Author: andreib
module alwcon17;
reg [7:0]a,b;
always (*b*)forever a=2;
endmodule
