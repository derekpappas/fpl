// Test type: Octal Numbers - x digit in octal value
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a=9'o1xX;
endmodule
