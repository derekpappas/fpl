// Test type: conditional_statement - if(expr) null else null
// Vparser rule name:
// Author: andreib
module conditional_statement3;
reg a,b,c;
initial if(a==b) ;
else ;
endmodule
