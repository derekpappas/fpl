//st0.vh