// Test type: Real numbers - all numbers part6
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=1234567890e9;
endmodule
