// Test type: Strings - Void String
// Vparser rule name:
// Author: andreib
module stringtest;
reg [8*32:1] stringvar;
initial begin
stringvar = "";
end
endmodule
