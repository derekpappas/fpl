`include "defines.v"

module cap();
// Location of source csl unit: file name = IPX2400.csl line number = 113
  `include "cap.logic.v"
endmodule

