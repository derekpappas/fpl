// Test type: Octal Numbers - spaces between size, base and value
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a=24 'o 23454761;
endmodule
