--THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
--COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
--OUTPUT FILE NAME  : x.vh
--FILE GENERATED ON : Fri Jul 30 07:13:06 2010

y.vhd
x.vhd
stim_expect_mem_template.vhd
tb.vhd
