`include "defines.v"

module hash();
// Location of source csl unit: file name = IPX2400.csl line number = 101
  `include "hash.logic.v"
endmodule

