`include "defines.v"

module proc(in);
// Location of source csl unit: file name = connect_output_to_input_u_to_u.csl line number = 2
  input [32 - 1:0] in;
  `include "proc.logic.v"
endmodule

