// Test type: Decimal Numbers - z digit variation
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=5'd?;
endmodule
