module hello_pli ();
  	 
initial begin
   $hello_2;
  // #10 $finish;
end
  	  
endmodule 