//test type : module_or_generate_item ::= always_construct
//vparser rule name : 
//author : Codrin
module test_0360(x,y);
 input x;
 output y;
 wire x;
 reg y;
 (* debug = 0 *)
 always @(x)
  y = x;
endmodule
