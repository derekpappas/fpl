// Test type: Continuous assignment - pl1, st0 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous391;
wire a;
assign (pull1, strong0) a=1'b1;
endmodule
