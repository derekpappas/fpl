// Test type: case_statement - casez - expression,expression,expression:null
// Vparser rule name:
// Author: andreib
module case_statement45;
reg a,b;
initial casez(a)
	4'bzZ?0,4'b0001,4'b0010:;
	endcase
endmodule
