`include "defines.v"

module r1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 286
  output [1 - 1:0] ar_sa0_s10;
  q1 q10(.ar_sa0_s10(ar_sa0_s10));
  `include "r1.logic.vh"
endmodule

