//this is a celldefine legal test
`celldefine //mycell
module mymodule;
endmodule

