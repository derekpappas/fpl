  --THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
--COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
--OUTPUT FILE NAME  : a0.vhd
--FILE GENERATED ON : Fri Aug 27 02:46:55 2010


library ieee ; 
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all; 
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;
 
use work.csl_util_package.all;

entity a0 is 
-- Location of source csl unit: file name = temp.csl line number = 1
  
        sa0  : in csl_bit_vector (0 downto 0)
 );
end a0 ; 

 architecture  arch_a0 of a0 is 

 begin 

 end  arch_a0 ; 
