`resetall
`default_nettype tri
module x;
endmodule
`resetall
