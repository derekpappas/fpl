// Test type: Decimal Numbers - lower case z digit
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=5'dz;
endmodule
