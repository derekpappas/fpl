`default_nettype tri
module yyy;
`include "../legal/default_nettype06.v"
wire x;
`default_nettype none
endmodule
