// Test type: initial statement - task_enable - no attribute instance
// Vparser rule name:
// Author: andreib
module initcon37;
reg a;
task test_task;
;
endtask
initial test_task;
endmodule
