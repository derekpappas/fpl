`include "defines.v"

module usb_analog_phy();
// Location of source csl unit: file name = generated/vizzini_core.csl line number = 156
  `include "usb_analog_phy.logic.v"
endmodule

