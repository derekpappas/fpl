a.vhd
b.vhd
