`include "defines.v"

module d0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 19
  input [1 - 1:0] ar_sa0_s10;
  c0 c0(.ar_sa0_s10(ar_sa0_s10));
  `include "d0.logic.vh"
endmodule

