//this is a celldefine legal test
/**/`celldefine//
module mod;
/**//***//**/`celldefine/***///sa
module mymodule;
endmodule
/****/`endcelldefine//haha
wire x;
/*hihi*/endmodule
/**/`endcelldefine//
