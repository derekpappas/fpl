// Test type: procedural continuous assignment - force net assignment
// Vparser rule name:
// Author: andreib
module procedural_continuous_assignment4;
wire a;
initial force a=1;
endmodule
