`include "defines.v"

module u_control();
// Location of source csl unit: file name = mbist_datapath.csl line number = 193
  endmodule

