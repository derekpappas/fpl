r_pc.vhd
r_caddr.vhd
m_im.vhd
rf.vhd
m_rom.vhd
u_es.vhd
u_ir.vhd
u_alu.vhd
r_ha.vhd
r_status.vhd
u_control.vhd
u_mbist.vhd
