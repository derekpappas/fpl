`include "defines.v"

module k0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 71
  input [1 - 1:0] ar_sa0_s10;
  j0 j0(.ar_sa0_s10(ar_sa0_s10));
  `include "k0.logic.vh"
endmodule

