-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./top_cslc_generated/code/vhdl/u_a.vhd
-- FILE GENERATED ON : Wed Mar 11 20:22:38 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u_a\ is
  port(\ck\ : in csl_bit;
       \reset\ : in csl_bit;
       \p_a_in\ : in csl_bit_vector(10#8# - 10#1# downto 10#0#);
       \p_a_out\ : out csl_bit_vector(10#8# - 10#1# downto 10#0#));
begin
end entity;

architecture \u_a_logic\ of \u_a\ is
begin
end architecture;

