//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : data_tcm.v
//FILE GENERATED ON : Wed Jul  9 20:26:20 2008

`include "defines.v"

module data_tcm();
// Location of source csl unit: file name = generated/mitch.csl line number = 33
  `include "data_tcm.logic.v"
endmodule

