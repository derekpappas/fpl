//this is a celldefine legal test
`resetall
module mod;
`celldefine
module mymodule;
endmodule
endmodule
`timescale 1ms/1fs

`endcelldefine
