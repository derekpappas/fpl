--THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
--COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
--OUTPUT FILE NAME  : a1.vhd
--FILE GENERATED ON : Fri Aug 27 02:46:56 2010


library ieee ; 
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all; 
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;
 
use work.csl_util_package.all;

entity a1 is 

 port ( -- Location of source csl unit: file name = temp.csl line number = 182

s10: out csl_bit_vector (0 downto 0)
 );
end a1 ; 

 architecture  arch_a1 of a1 is 

ar_sa0_s10 : in   csl_bit_vector(0 downto 0) 
 begin 

 end  arch_a1 ; 
