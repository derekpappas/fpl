-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./v_top_cslc_generated/code/vhdl/io_cell.vhd
-- FILE GENERATED ON : Tue Sep 30 16:36:13 2008
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \io_cell\ is
  port(\pad_in\ : out csl_bit;
       \pad_out\ : in csl_bit;
       \pad_en\ : in csl_bit;
       \pad_pin\ : inout csl_bit);
begin
end entity;

architecture \io_cell_logic\ of \io_cell\ is
begin
end architecture;

