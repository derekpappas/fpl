//test type : block_item_declaration ::= time list_of_block_variable_identifiers;
//vparser rule name : 
//author : Codrin
module test_0510;
  (* timeset, timer = "start" *)
  time start, tend, tpause;
endmodule
