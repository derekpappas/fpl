a.vhd
b.vhd
stim_expect_mem_template.vhd
tb.vhd
