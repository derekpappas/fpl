// Test type: Continuous assignment - list_of_net_assignments - 3 elements
// Vparser rule name:
// Author: andreib
module continuous3;
wire a,b,c;
assign a=1'b1, b=1'b0, c=1'd2;
endmodule
