a1.vhd
b1.vhd
