// Test type: conditional_statement - if(expr) null
// Vparser rule name:
// Author: andreib
module conditional_statement1;
reg a,b,c;
initial if(a==b) ;
endmodule
