// Test type: conditional_statement - if(expr) statement else null
// Vparser rule name:
// Author: andreib
module conditional_statement5;
reg a,b,c;
initial if(a==b) c=1;
else ;
endmodule
