//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : eth_io.v
//FILE GENERATED ON : Thu Jun 19 15:32:42 2008

`include "defines.v"

module eth_io();
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 25
  `include "eth_io.logic.v"
endmodule

