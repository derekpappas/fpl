//test type : module_or_generate_item ::= initial_construct
//vparser rule name : 
//author : Codrin
module test_0350;
 reg x;
 (* debug = 1, errors = 0 *)
 initial
  x = 1'b0;
endmodule
