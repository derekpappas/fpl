//test type : port_declaration
//vparser rule name : 
//author : Codrin
module declaration_0110(x);
 (* a , b = 1 *) output x;
endmodule
