// Test type: Octal Numbers - underscore within size and value
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a=1_2'o12__34;
endmodule
