// Test type: Continuous assignment - st1, sup0 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous316;
wire a;
assign (strong1, supply0) a=1'b1;
endmodule
