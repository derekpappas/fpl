-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./u_mbist_cslc_generated/code/vhdl/u_arith.vhd
-- FILE GENERATED ON : Wed Nov 18 19:49:32 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u_arith\ is
  port(\ifc_op0_op1\ : in csl_bit_vector(10#15# downto 10#0#);
       \ifc_op0_op2\ : in csl_bit_vector(10#15# downto 10#0#);
       \ifc_sel0_sel\ : in csl_bit_vector(10#3# downto 10#0#);
       \ifc_out0_o\ : out csl_bit_vector(10#15# downto 10#0#);
       \cin\ : in csl_bit;
       \cout\ : out csl_bit);
begin
end entity;

architecture \u_arith_logic\ of \u_arith\ is
begin
end architecture;

