// Test type: Binary Numbers - Size with underscores
// Vparser rule name: Numbers
// Author: andreib
module binary_num;
wire a;
assign a=1_5'b1011011011;
endmodule
