// Test type: Hex Numbers - spaces between size, base and value
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=8 'h 2A;
endmodule
