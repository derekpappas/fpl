`include "defines.v"

module c0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 13
  input [1 - 1:0] ar_sa0_s10;
  b0 b0(.ar_sa0_s10(ar_sa0_s10));
  `include "c0.logic.vh"
endmodule

