//test type : {constant_expression concatenation}
//vparser rule name : 
//author : Bogdan Mereghea
module multiple_concatenation1;
    wire a;
    assign a = {0{1'b1}};
endmodule
