u_a.vhd
u_b.vhd
u_c.vhd
u_d.vhd
u_top.vhd
