`include "defines.v"

module p0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 107
  input [1 - 1:0] ar_sa0_s10;
  o0 o0(.ar_sa0_s10(ar_sa0_s10));
  `include "p0.logic.vh"
endmodule

