// Test type: Decimal Numbers - upper case decimal base
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=5'D16;
endmodule
