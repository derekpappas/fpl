// Test type: Octal Numbers - variation of sign/base letter case
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a=9'sO123;
endmodule
