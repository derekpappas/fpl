//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : fabric_add.v
//FILE GENERATED ON : Wed Jul  9 20:26:20 2008

`include "defines.v"

module fabric_add();
// Location of source csl unit: file name = generated/mitch.csl line number = 19
  `include "fabric_add.logic.v"
endmodule

