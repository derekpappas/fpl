//test type : port_declaration
//vparser rule name : 
//author : Codrin
module declaration_0120(x);
 (* a = 2 , b, c = 0 *) output x;
endmodule
