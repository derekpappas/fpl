// Test type: Continuous assignment - h1, sup0 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous676;
wire a;
assign (highz1, supply0) a=1'b1;
endmodule
