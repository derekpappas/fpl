// Test type: Continuous assignment - wk0, h1 - list_of_net_assignments - 2 elements
// Vparser rule name:
// Author: andreib
module continuous542;
wire a,b;
assign (weak0, highz1) a=1'b1, b=1'b0;
endmodule
