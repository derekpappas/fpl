//test type : module_declaration
//vparser rule name : 
//author : Codrin
(* a *)
(* a = 1 *)
(* a, b *)
(* a = 1, b *)
module declaration_030;
endmodule
