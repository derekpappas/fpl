
module new_sigs;

parameter signed p1 = 0;
parameter [31:0] p2 = 0;
parameter signed [31:0] p3 = 0;
parameter integer p4 = 0;
parameter real p5 = 0;
parameter realtime p6 = 0;
parameter time p7 = 0;


realtime rt;
trior t_or;

endmodule
