// Test type: Continuous assignment - wk1, st0 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous451;
wire a;
assign (weak1, strong0) a=1'b1;
endmodule
