module hwb30(x,z);
    input [30:1] x;
    output z;

    wire [4:0] sum;

    assign sum =
	{4'b0,x[30]} +
	{4'b0,x[29]} +
	{4'b0,x[28]} +
	{4'b0,x[27]} +
	{4'b0,x[26]} +
	{4'b0,x[25]} +
	{4'b0,x[24]} +
	{4'b0,x[23]} +
	{4'b0,x[22]} +
	{4'b0,x[21]} +
	{4'b0,x[20]} +
	{4'b0,x[19]} +
	{4'b0,x[18]} +
	{4'b0,x[17]} +
	{4'b0,x[16]} +
	{4'b0,x[15]} +
	{4'b0,x[14]} +
	{4'b0,x[13]} +
	{4'b0,x[12]} +
	{4'b0,x[11]} +
	{4'b0,x[10]} +
	{4'b0,x[9]} +
	{4'b0,x[8]} +
	{4'b0,x[7]} +
	{4'b0,x[6]} +
	{4'b0,x[5]} +
	{4'b0,x[4]} +
	{4'b0,x[3]} +
	{4'b0,x[2]} +
	{4'b0,x[1]};

    assign z = 
	x[30] & (sum == 30) |
	x[29] & (sum == 29) |
	x[28] & (sum == 28) |
	x[27] & (sum == 27) |
	x[26] & (sum == 26) |
	x[25] & (sum == 25) |
	x[24] & (sum == 24) |
	x[23] & (sum == 23) |
	x[22] & (sum == 22) |
	x[21] & (sum == 21) |
	x[20] & (sum == 20) |
	x[19] & (sum == 19) |
	x[18] & (sum == 18) |
	x[17] & (sum == 17) |
	x[16] & (sum == 16) |
	x[15] & (sum == 15) |
	x[14] & (sum == 14) |
	x[13] & (sum == 13) |
	x[12] & (sum == 12) |
	x[11] & (sum == 11) |
	x[10] & (sum == 10) |
	x[9] & (sum == 9) |
	x[8] & (sum == 8) |
	x[7] & (sum == 7) |
	x[6] & (sum == 6) |
	x[5] & (sum == 5) |
	x[4] & (sum == 4) |
	x[3] & (sum == 3) |
	x[2] & (sum == 2) |
	x[1] & (sum == 1);

endmodule // hwb
