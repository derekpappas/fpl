//test type : task_item_declaration ::= inout_declaration
//vparser rule name : 
//author : Codrin
//fixed by: Gabrield
module test_0440;
 (* carry, text = "error" *)
 task string;
  inout a;
  ;
 endtask
endmodule
