// Test type: delay_control - delay_value - real number
// Vparser rule name:
// Author: andreib
module delay_control2;
reg a;
initial #1e1 a=1'b1;
endmodule
