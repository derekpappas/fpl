// Test type: Real numbers - real number with underscore
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=27___4.32;
endmodule
