//test type : number binary_operator_** hierarchical_identifier
//vparser rule name : 
//author : Bogdan Mereghea
module binary_operator187;
    reg a, b;
    initial begin
        a = 1'b1 ** b;
    end
endmodule
