// Test type: delay_or_event_control - delay_control - mintypmax
// Vparser rule name:
// Author: andreib
module delay_or_event_control2;
reg a;
initial #(4:5:6) a=1'b1;
endmodule
