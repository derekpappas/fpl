// Test type: procedural continuous assignment - release net assignment
// Vparser rule name:
// Author: andreib
module procedural_continuous_assignment6;
wire a;
initial release a;
endmodule
