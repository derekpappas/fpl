// Test type: Continuous assignment - pl0, wk1 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous181;
wire a;
assign (pull0, weak1) a=1'b1;
endmodule
