`include "defines.v"

module j1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 238
  output [1 - 1:0] ar_sa0_s10;
  i1 i10(.ar_sa0_s10(ar_sa0_s10));
  `include "j1.logic.vh"
endmodule

