`include "defines.v"

module sramctrl();
// Location of source csl unit: file name = IPX2400.csl line number = 89
  `include "sramctrl.logic.v"
endmodule

