// Test type: procedural continuous assignment - release variable assignment
// Vparser rule name:
// Author: andreib
module procedural_continuous_assignment5;
reg a;
initial release a;
endmodule
