u_mem.vhd
u_top.vhd
