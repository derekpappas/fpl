//Primitive Instantiation and Instances: gate_instantiation = enable_gatetype ... ;
//tests by GabrielD
module gate_instantiation_enable_gatetype0;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype1;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype2;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype3;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype4;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype6;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype7;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype8;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype9;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype10;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype12;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype13;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype14;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype15;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype16;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype18;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype19;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype20;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype21;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype22;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype24;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype25;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype26;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype27;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype28;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype30;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype31;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype32;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype33;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype34;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype36;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype37;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype38;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype39;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype40;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype42;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype43;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype44;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype45;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype46;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype48;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype49;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype50;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype51;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype52;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype54;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype55;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype56;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype57;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype58;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype60;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype61;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype62;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype63;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype64;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype66;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype67;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype68;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype69;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype70;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype72;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype73;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype74;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype75;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype76;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype78;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype79;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype80;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype81;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype82;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( strong1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype84;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype85;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype86;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype87;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype88;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype90;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype91;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype92;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype93;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype94;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype96;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype97;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype98;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype99;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype100;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype102;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype103;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype104;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype105;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype106;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( weak1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype108;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype109;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype110;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype111;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype112;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype114;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype115;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype116;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype117;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype118;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype120;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype121;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype122;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype123;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype124;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype126;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype127;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype128;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype129;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype130;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype132;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype133;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype134;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype135;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype136;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype138;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype139;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype140;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype141;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype142;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype144;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype145;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype146;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype147;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype148;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype150;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype151;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype152;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype153;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype154;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype156;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, strong1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype157;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype158;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype159;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype160;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype162;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype163;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype164;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype165;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype166;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype168;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, weak1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype169;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype170;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype171;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype172;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype174;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype175;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype176;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype177;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype178;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz0, weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype180;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, supply0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype181;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype182;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype183;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype184;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype186;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype187;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype188;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype189;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype190;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype192;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, pull0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype193;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype194;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype195;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype196;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype198;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype199;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype200;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype201;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype202;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif0 (highz1, pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype204;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype205;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype206;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype207;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype208;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype210;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype211;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype212;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype213;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype214;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype216;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype217;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype218;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype219;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype220;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype222;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype223;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype224;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype225;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype226;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype228;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype229;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype230;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype231;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype232;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype234;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype235;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype236;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype237;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype238;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype240;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype241;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype242;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype243;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype244;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype246;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype247;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype248;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype249;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype250;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype252;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype253;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype254;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype255;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype256;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype258;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype259;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype260;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype261;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype262;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype264;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype265;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype266;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype267;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype268;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype270;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype271;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype272;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype273;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype274;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype276;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype277;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype278;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype279;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype280;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype282;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype283;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype284;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype285;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype286;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( strong1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype288;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype289;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype290;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype291;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype292;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype294;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype295;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype296;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype297;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype298;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype300;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype301;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype302;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype303;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype304;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype306;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype307;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype308;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype309;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype310;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( weak1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype312;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype313;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype314;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype315;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype316;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype318;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype319;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype320;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype321;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype322;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype324;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype325;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype326;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype327;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype328;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype330;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype331;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype332;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype333;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype334;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype336;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype337;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype338;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype339;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype340;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype342;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype343;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype344;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype345;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype346;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype348;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype349;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype350;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype351;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype352;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype354;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype355;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype356;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype357;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype358;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype360;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, strong1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype361;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype362;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype363;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype364;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype366;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype367;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype368;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype369;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype370;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype372;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, weak1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype373;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype374;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype375;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype376;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype378;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype379;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype380;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype381;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype382;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz0, weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype384;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, supply0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype385;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype386;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype387;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype388;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype390;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype391;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype392;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype393;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype394;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype396;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, pull0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype397;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype398;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype399;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype400;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype402;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype403;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype404;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype405;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype406;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  bufif1 (highz1, pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype408;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype409;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype410;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype411;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype412;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype414;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype415;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype416;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype417;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype418;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype420;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype421;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype422;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype423;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype424;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype426;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype427;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype428;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype429;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype430;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype432;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype433;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype434;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype435;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype436;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype438;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype439;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype440;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype441;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype442;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype444;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype445;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype446;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype447;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype448;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype450;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype451;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype452;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype453;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype454;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype456;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype457;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype458;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype459;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype460;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype462;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype463;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype464;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype465;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype466;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype468;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype469;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype470;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype471;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype472;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype474;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype475;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype476;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype477;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype478;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype480;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype481;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype482;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype483;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype484;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype486;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype487;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype488;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype489;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype490;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( strong1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype492;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype493;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype494;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype495;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype496;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype498;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype499;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype500;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype501;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype502;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype504;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype505;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype506;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype507;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype508;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype510;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype511;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype512;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype513;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype514;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( weak1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype516;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype517;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype518;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype519;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype520;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype522;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype523;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype524;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype525;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype526;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype528;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype529;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype530;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype531;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype532;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype534;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype535;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype536;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype537;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype538;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype540;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype541;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype542;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype543;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype544;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype546;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype547;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype548;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype549;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype550;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype552;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype553;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype554;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype555;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype556;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype558;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype559;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype560;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype561;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype562;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype564;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, strong1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype565;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype566;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype567;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype568;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype570;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype571;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype572;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype573;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype574;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype576;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, weak1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype577;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype578;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype579;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype580;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype582;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype583;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype584;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype585;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype586;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz0, weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype588;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, supply0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype589;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype590;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype591;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype592;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype594;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype595;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype596;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype597;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype598;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype600;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, pull0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype601;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype602;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype603;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype604;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype606;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype607;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype608;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype609;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype610;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif0 (highz1, pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype612;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype613;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype614;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype615;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype616;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype618;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype619;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype620;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype621;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype622;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype624;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype625;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype626;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype627;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype628;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype630;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype631;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype632;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype633;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype634;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype636;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype637;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype638;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype639;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype640;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype642;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype643;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype644;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype645;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype646;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype648;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype649;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype650;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype651;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype652;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype654;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype655;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype656;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype657;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype658;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype660;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype661;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype662;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype663;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype664;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype666;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype667;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype668;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype669;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype670;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 , weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype672;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype673;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype674;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype675;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype676;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype678;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype679;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype680;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype681;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype682;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype684;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype685;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype686;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype687;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype688;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype690;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype691;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype692;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype693;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype694;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( strong1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype696;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype697;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype698;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype699;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype700;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype702;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype703;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype704;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype705;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype706;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype708;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype709;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype710;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype711;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype712;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype714;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype715;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype716;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype717;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype718;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( weak1 , pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype720;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype721;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype722;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype723;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype724;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype726;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype727;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype728;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype729;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype730;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype732;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype733;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype734;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype735;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype736;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype738;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype739;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype740;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype741;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype742;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype744;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype745;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype746;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype747;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype748;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype750;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype751;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype752;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype753;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype754;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( supply0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype756;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype757;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype758;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype759;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype760;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype762;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype763;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype764;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype765;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype766;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 ( pull0 ,highz1) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype768;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, strong1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype769;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype770;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, strong1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype771;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype772;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, strong1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype774;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype775;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype776;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, strong1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype777;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype778;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, strong1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype780;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, weak1 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype781;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype782;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, weak1 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype783;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype784;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, weak1 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype786;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype787;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype788;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, weak1 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype789;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype790;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz0, weak1 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype791;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, supply0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype793;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype794;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, supply0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype795;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype796;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, supply0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype799;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype800;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, supply0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype801;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype802;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, supply0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype804;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, pull0 ) (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype805;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype806;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, pull0 ) (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype807;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype808;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, pull0 ) name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype810;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype811;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype812;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, pull0 ) #3 (output_terminal,input_terminal,ncontrol_terminal) , name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype813;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
module gate_instantiation_enable_gatetype814;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  notif1 (highz1, pull0 ) #3 name_of_gate_instance (output_terminal,input_terminal,ncontrol_terminal) , (output_terminal,input_terminal,ncontrol_terminal) ;
endmodule
