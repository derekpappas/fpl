module mygrandparents;
`define x
`ifdef x
  `define x \
\
\
reg x3;
reg x33;
  `define y endmodule
`endif

`x
`y
