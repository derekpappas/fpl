-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./c_cslc_generated/code/vhdl/a.vhd
-- FILE GENERATED ON : Fri Nov 27 06:35:43 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \a\ is
  port(\ifc00_p_m\ : in csl_bit_vector(10#78# - 10#1# downto 10#0#);
       \ifc00_p_n\ : out csl_bit_vector(10#64# - 10#1# downto 10#0#);
       \ifc00_p_o\ : in csl_bit_vector(10#78# - 10#1# downto 10#0#);
       \p_n\ : inout csl_bit_vector(10#64# - 10#1# downto 10#0#));
begin
end entity;

architecture \a_logic\ of \a\ is
begin
end architecture;

