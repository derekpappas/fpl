// Test type: Octal Numbers - all numbers
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a=24'o01234567;
endmodule
