// Test type: Hex Numbers - ? (z) digit
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=12'h7??;
endmodule
