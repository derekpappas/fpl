`include "defines.v"

module xpi();
// Location of source csl unit: file name = IPX2400.csl line number = 232
  `include "xpi.logic.v"
endmodule

