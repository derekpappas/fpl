// Test type: Real numbers - all numbers part4
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=1234567890e67;
endmodule
