`include "defines.v"

module ctrlstore();
// Location of source csl unit: file name = IPX2400.csl line number = 28
  `include "ctrlstore.logic.v"
endmodule

