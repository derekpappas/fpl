// Test type: Continuous assignment - wk0, h1 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous541;
wire a;
assign (weak0, highz1) a=1'b1;
endmodule
