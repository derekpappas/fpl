`ifndef CTU_SYNC
`define CTU_SYNC

module ctu_synchronizer;
endmodule

module ctu_synch_ref_jl;
endmodule

module ctu_or2;
endmodule

module ctu_inv;
endmodule

module ctu_nor2;
endmodule

module ctu_and2;
endmodule

module ctu_dft_jtag_tap;
endmodule

module ctu_mux21;
endmodule

module ctu_jtag_clk_sel_0_0_ff;
endmodule

module ctu_jtag_clk_sel_1_0_ff;
endmodule

module ctu_jtag_clk_sel_0_1_ff;
endmodule

`endif
