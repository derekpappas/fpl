// Test type: Binary Numbers - with ? digits
// Vparser rule name: Numbers
// Author: andreib
module binary_num;
wire a;
assign a=5'b011??;
endmodule
