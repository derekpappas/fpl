//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : i2c_lba.v
//FILE GENERATED ON : Tue Jun 17 01:23:46 2008

`include "defines.v"

module i2c_lba(lbadummy3,
               lbdummy2);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 29
  input lbdummy2;
  output lbadummy3;
  `include "i2c_lba.logic.v"
endmodule

