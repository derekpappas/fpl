-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./u_mbist_cslc_generated/code/vhdl/u_mux41.vhd
-- FILE GENERATED ON : Wed Nov 18 19:49:32 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u_mux41\ is
  port(\in0\ : in csl_bit_vector(10#15# downto 10#0#);
       \in1\ : in csl_bit_vector(10#15# downto 10#0#);
       \in2\ : in csl_bit_vector(10#15# downto 10#0#);
       \in3\ : in csl_bit_vector(10#15# downto 10#0#);
       \sel\ : in csl_bit_vector(10#4# - 10#1# downto 10#0#);
       \ifc_out0_o\ : out csl_bit_vector(10#15# downto 10#0#));
begin
end entity;

architecture \u_mux41_logic\ of \u_mux41\ is
begin
end architecture;

