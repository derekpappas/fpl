// Test type: Hex Numbers - underscore within size and value
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=1_6'hC2_d3_;
endmodule
