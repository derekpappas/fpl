//test type : module_or_generate_item ::= module_or_generate_item_declaration (task_declaration)
//vparser rule name : 
//author : Codrin
//fixed by: Gabrield
module test_0240;
 (* tasklist *)
 task foo;
  ;
 endtask
endmodule
