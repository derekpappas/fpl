//cd.vh