// Test type: Continuous assignment - h0, sup1 - list_of_net_assignments - 2 elements
// Vparser rule name:
// Author: andreib
module continuous617;
wire a,b;
assign (highz0, supply1) a=1'b1, b=1'b0;
endmodule
