//test type : block_item_declaration ::= reg[signed][range] list_of_block_variable_identifiers;
//vparser rule name : 
//author : Codrin
module test_0490;
  (* debug, size *)
  reg [7:0] bus, data, address;
endmodule
