// Test type: Decimal Numbers - upper case signed and lower case decimal base
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=5'Sd2___9;
endmodule
