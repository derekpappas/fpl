// Test type: Strings - 1 char tring
// Vparser rule name:
// Author: andreib
module stringtest;
reg [8*32:1] stringvar;
initial begin
stringvar = "a";
end
endmodule
