`include "defines.v"

module m_rom();
// Location of source csl unit: file name = mbist_datapath.csl line number = 110
// The depth of memory module m_rom is of illegal type. Depth set to 1.
// The width of memory module m_rom is of illegal type. Width set to 1.
  endmodule

