`include "defines.v"

module c1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 195
  output [1 - 1:0] ar_sa0_s10;
  b1 b10(.ar_sa0_s10(ar_sa0_s10));
  `include "c1.logic.vh"
endmodule

