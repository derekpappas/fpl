// Test type: Continuous assignment - sup1, pl0 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous286;
wire a;
assign (supply1, pull0) a=1'b1;
endmodule
