-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./proc_ring_cslc_generated/code/vhdl/fabric_dma.vhd
-- FILE GENERATED ON : Wed Jul  9 20:26:20 2008
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \fabric_dma\ is
  port(\sbfdstart\ : in csl_bit;
       \sbfdbusy\ : out csl_bit);
begin
end entity;

architecture \fabric_dma_logic\ of \fabric_dma\ is
begin
end architecture;

