`include "defines.v"

module opmux();
// Location of source csl unit: file name = IPX2400.csl line number = 61
  `include "opmux.logic.v"
endmodule

