module testbench_inout_declaration;
    inout_declaration0 inout_declaration_instance0();
    inout_declaration1 inout_declaration_instance1();
    inout_declaration2 inout_declaration_instance2();
    inout_declaration3 inout_declaration_instance3();
    inout_declaration4 inout_declaration_instance4();
    inout_declaration5 inout_declaration_instance5();
    inout_declaration6 inout_declaration_instance6();
    inout_declaration7 inout_declaration_instance7();
    inout_declaration8 inout_declaration_instance8();
    inout_declaration9 inout_declaration_instance9();
    inout_declaration10 inout_declaration_instance10();
    inout_declaration11 inout_declaration_instance11();
    inout_declaration12 inout_declaration_instance12();
    inout_declaration13 inout_declaration_instance13();
    inout_declaration14 inout_declaration_instance14();
    inout_declaration15 inout_declaration_instance15();
    inout_declaration16 inout_declaration_instance16();
    inout_declaration17 inout_declaration_instance17();
    inout_declaration18 inout_declaration_instance18();
    inout_declaration19 inout_declaration_instance19();
    inout_declaration20 inout_declaration_instance20();
    inout_declaration21 inout_declaration_instance21();
    inout_declaration22 inout_declaration_instance22();
    inout_declaration23 inout_declaration_instance23();
    inout_declaration24 inout_declaration_instance24();
    inout_declaration25 inout_declaration_instance25();
    inout_declaration26 inout_declaration_instance26();
    inout_declaration27 inout_declaration_instance27();
    inout_declaration28 inout_declaration_instance28();
    inout_declaration29 inout_declaration_instance29();
    inout_declaration30 inout_declaration_instance30();
    inout_declaration31 inout_declaration_instance31();
    inout_declaration32 inout_declaration_instance32();
    inout_declaration33 inout_declaration_instance33();
    inout_declaration34 inout_declaration_instance34();
    inout_declaration35 inout_declaration_instance35();
    inout_declaration36 inout_declaration_instance36();
    inout_declaration37 inout_declaration_instance37();
    inout_declaration38 inout_declaration_instance38();
    inout_declaration39 inout_declaration_instance39();
    inout_declaration40 inout_declaration_instance40();
    inout_declaration41 inout_declaration_instance41();
    inout_declaration42 inout_declaration_instance42();
    inout_declaration43 inout_declaration_instance43();
    inout_declaration44 inout_declaration_instance44();
    inout_declaration45 inout_declaration_instance45();
    inout_declaration46 inout_declaration_instance46();
    inout_declaration47 inout_declaration_instance47();
    inout_declaration48 inout_declaration_instance48();
    inout_declaration49 inout_declaration_instance49();
    inout_declaration50 inout_declaration_instance50();
    inout_declaration51 inout_declaration_instance51();
    inout_declaration52 inout_declaration_instance52();
    inout_declaration53 inout_declaration_instance53();
    inout_declaration54 inout_declaration_instance54();
    inout_declaration55 inout_declaration_instance55();
    inout_declaration56 inout_declaration_instance56();
    inout_declaration57 inout_declaration_instance57();
    inout_declaration58 inout_declaration_instance58();
    inout_declaration59 inout_declaration_instance59();
    inout_declaration60 inout_declaration_instance60();
    inout_declaration61 inout_declaration_instance61();
    inout_declaration62 inout_declaration_instance62();
    inout_declaration63 inout_declaration_instance63();
    inout_declaration64 inout_declaration_instance64();
    inout_declaration65 inout_declaration_instance65();
    inout_declaration66 inout_declaration_instance66();
    inout_declaration67 inout_declaration_instance67();
    inout_declaration68 inout_declaration_instance68();
    inout_declaration69 inout_declaration_instance69();
    inout_declaration70 inout_declaration_instance70();
    inout_declaration71 inout_declaration_instance71();
    inout_declaration72 inout_declaration_instance72();
    inout_declaration73 inout_declaration_instance73();
    inout_declaration74 inout_declaration_instance74();
    inout_declaration75 inout_declaration_instance75();
    inout_declaration76 inout_declaration_instance76();
    inout_declaration77 inout_declaration_instance77();
    inout_declaration78 inout_declaration_instance78();
    inout_declaration79 inout_declaration_instance79();
    inout_declaration80 inout_declaration_instance80();
    inout_declaration81 inout_declaration_instance81();
    inout_declaration82 inout_declaration_instance82();
    inout_declaration83 inout_declaration_instance83();
    inout_declaration84 inout_declaration_instance84();
    inout_declaration85 inout_declaration_instance85();
    inout_declaration86 inout_declaration_instance86();
    inout_declaration87 inout_declaration_instance87();
    inout_declaration88 inout_declaration_instance88();
    inout_declaration89 inout_declaration_instance89();
    inout_declaration90 inout_declaration_instance90();
    inout_declaration91 inout_declaration_instance91();
    inout_declaration92 inout_declaration_instance92();
    inout_declaration93 inout_declaration_instance93();
    inout_declaration94 inout_declaration_instance94();
    inout_declaration95 inout_declaration_instance95();
    inout_declaration96 inout_declaration_instance96();
    inout_declaration97 inout_declaration_instance97();
    inout_declaration98 inout_declaration_instance98();
    inout_declaration99 inout_declaration_instance99();
    inout_declaration100 inout_declaration_instance100();
    inout_declaration101 inout_declaration_instance101();
    inout_declaration102 inout_declaration_instance102();
    inout_declaration103 inout_declaration_instance103();
    inout_declaration104 inout_declaration_instance104();
    inout_declaration105 inout_declaration_instance105();
    inout_declaration106 inout_declaration_instance106();
    inout_declaration107 inout_declaration_instance107();
    inout_declaration108 inout_declaration_instance108();
    inout_declaration109 inout_declaration_instance109();
    inout_declaration110 inout_declaration_instance110();
    inout_declaration111 inout_declaration_instance111();
    inout_declaration112 inout_declaration_instance112();
    inout_declaration113 inout_declaration_instance113();
    inout_declaration114 inout_declaration_instance114();
    inout_declaration115 inout_declaration_instance115();
    inout_declaration116 inout_declaration_instance116();
    inout_declaration117 inout_declaration_instance117();
    inout_declaration118 inout_declaration_instance118();
    inout_declaration119 inout_declaration_instance119();
    inout_declaration120 inout_declaration_instance120();
    inout_declaration121 inout_declaration_instance121();
    inout_declaration122 inout_declaration_instance122();
    inout_declaration123 inout_declaration_instance123();
    inout_declaration124 inout_declaration_instance124();
    inout_declaration125 inout_declaration_instance125();
    inout_declaration126 inout_declaration_instance126();
    inout_declaration127 inout_declaration_instance127();
    inout_declaration128 inout_declaration_instance128();
    inout_declaration129 inout_declaration_instance129();
    inout_declaration130 inout_declaration_instance130();
    inout_declaration131 inout_declaration_instance131();
    inout_declaration132 inout_declaration_instance132();
    inout_declaration133 inout_declaration_instance133();
    inout_declaration134 inout_declaration_instance134();
    inout_declaration135 inout_declaration_instance135();
    inout_declaration136 inout_declaration_instance136();
    inout_declaration137 inout_declaration_instance137();
    inout_declaration138 inout_declaration_instance138();
    inout_declaration139 inout_declaration_instance139();
    inout_declaration140 inout_declaration_instance140();
    inout_declaration141 inout_declaration_instance141();
    inout_declaration142 inout_declaration_instance142();
    inout_declaration143 inout_declaration_instance143();
    inout_declaration144 inout_declaration_instance144();
    inout_declaration145 inout_declaration_instance145();
    inout_declaration146 inout_declaration_instance146();
    inout_declaration147 inout_declaration_instance147();
    inout_declaration148 inout_declaration_instance148();
    inout_declaration149 inout_declaration_instance149();
    inout_declaration150 inout_declaration_instance150();
    inout_declaration151 inout_declaration_instance151();
    inout_declaration152 inout_declaration_instance152();
    inout_declaration153 inout_declaration_instance153();
    inout_declaration154 inout_declaration_instance154();
    inout_declaration155 inout_declaration_instance155();
    inout_declaration156 inout_declaration_instance156();
    inout_declaration157 inout_declaration_instance157();
    inout_declaration158 inout_declaration_instance158();
    inout_declaration159 inout_declaration_instance159();
    inout_declaration160 inout_declaration_instance160();
    inout_declaration161 inout_declaration_instance161();
    inout_declaration162 inout_declaration_instance162();
    inout_declaration163 inout_declaration_instance163();
    inout_declaration164 inout_declaration_instance164();
    inout_declaration165 inout_declaration_instance165();
    inout_declaration166 inout_declaration_instance166();
    inout_declaration167 inout_declaration_instance167();
    inout_declaration168 inout_declaration_instance168();
    inout_declaration169 inout_declaration_instance169();
    inout_declaration170 inout_declaration_instance170();
    inout_declaration171 inout_declaration_instance171();
    inout_declaration172 inout_declaration_instance172();
    inout_declaration173 inout_declaration_instance173();
    inout_declaration174 inout_declaration_instance174();
    inout_declaration175 inout_declaration_instance175();
    inout_declaration176 inout_declaration_instance176();
    inout_declaration177 inout_declaration_instance177();
    inout_declaration178 inout_declaration_instance178();
    inout_declaration179 inout_declaration_instance179();
    inout_declaration180 inout_declaration_instance180();
    inout_declaration181 inout_declaration_instance181();
    inout_declaration182 inout_declaration_instance182();
    inout_declaration183 inout_declaration_instance183();
    inout_declaration184 inout_declaration_instance184();
    inout_declaration185 inout_declaration_instance185();
    inout_declaration186 inout_declaration_instance186();
    inout_declaration187 inout_declaration_instance187();
    inout_declaration188 inout_declaration_instance188();
    inout_declaration189 inout_declaration_instance189();
    inout_declaration190 inout_declaration_instance190();
    inout_declaration191 inout_declaration_instance191();
    inout_declaration192 inout_declaration_instance192();
    inout_declaration193 inout_declaration_instance193();
    inout_declaration194 inout_declaration_instance194();
    inout_declaration195 inout_declaration_instance195();
    inout_declaration196 inout_declaration_instance196();
    inout_declaration197 inout_declaration_instance197();
    inout_declaration198 inout_declaration_instance198();
    inout_declaration199 inout_declaration_instance199();
    inout_declaration200 inout_declaration_instance200();
    inout_declaration201 inout_declaration_instance201();
    inout_declaration202 inout_declaration_instance202();
    inout_declaration203 inout_declaration_instance203();
    inout_declaration204 inout_declaration_instance204();
    inout_declaration205 inout_declaration_instance205();
    inout_declaration206 inout_declaration_instance206();
    inout_declaration207 inout_declaration_instance207();
    inout_declaration208 inout_declaration_instance208();
    inout_declaration209 inout_declaration_instance209();
    inout_declaration210 inout_declaration_instance210();
    inout_declaration211 inout_declaration_instance211();
    inout_declaration212 inout_declaration_instance212();
    inout_declaration213 inout_declaration_instance213();
    inout_declaration214 inout_declaration_instance214();
    inout_declaration215 inout_declaration_instance215();
    inout_declaration216 inout_declaration_instance216();
    inout_declaration217 inout_declaration_instance217();
    inout_declaration218 inout_declaration_instance218();
    inout_declaration219 inout_declaration_instance219();
    inout_declaration220 inout_declaration_instance220();
    inout_declaration221 inout_declaration_instance221();
    inout_declaration222 inout_declaration_instance222();
    inout_declaration223 inout_declaration_instance223();
    inout_declaration224 inout_declaration_instance224();
    inout_declaration225 inout_declaration_instance225();
    inout_declaration226 inout_declaration_instance226();
    inout_declaration227 inout_declaration_instance227();
    inout_declaration228 inout_declaration_instance228();
    inout_declaration229 inout_declaration_instance229();
    inout_declaration230 inout_declaration_instance230();
    inout_declaration231 inout_declaration_instance231();
    inout_declaration232 inout_declaration_instance232();
    inout_declaration233 inout_declaration_instance233();
    inout_declaration234 inout_declaration_instance234();
    inout_declaration235 inout_declaration_instance235();
    inout_declaration236 inout_declaration_instance236();
    inout_declaration237 inout_declaration_instance237();
    inout_declaration238 inout_declaration_instance238();
    inout_declaration239 inout_declaration_instance239();
    inout_declaration240 inout_declaration_instance240();
    inout_declaration241 inout_declaration_instance241();
    inout_declaration242 inout_declaration_instance242();
    inout_declaration243 inout_declaration_instance243();
    inout_declaration244 inout_declaration_instance244();
    inout_declaration245 inout_declaration_instance245();
    inout_declaration246 inout_declaration_instance246();
    inout_declaration247 inout_declaration_instance247();
    inout_declaration248 inout_declaration_instance248();
    inout_declaration249 inout_declaration_instance249();
    inout_declaration250 inout_declaration_instance250();
    inout_declaration251 inout_declaration_instance251();
    inout_declaration252 inout_declaration_instance252();
    inout_declaration253 inout_declaration_instance253();
    inout_declaration254 inout_declaration_instance254();
    inout_declaration255 inout_declaration_instance255();
    inout_declaration256 inout_declaration_instance256();
    inout_declaration257 inout_declaration_instance257();
    inout_declaration258 inout_declaration_instance258();
    inout_declaration259 inout_declaration_instance259();
    inout_declaration260 inout_declaration_instance260();
    inout_declaration261 inout_declaration_instance261();
    inout_declaration262 inout_declaration_instance262();
    inout_declaration263 inout_declaration_instance263();
    inout_declaration264 inout_declaration_instance264();
    inout_declaration265 inout_declaration_instance265();
    inout_declaration266 inout_declaration_instance266();
    inout_declaration267 inout_declaration_instance267();
    inout_declaration268 inout_declaration_instance268();
    inout_declaration269 inout_declaration_instance269();
    inout_declaration270 inout_declaration_instance270();
    inout_declaration271 inout_declaration_instance271();
    inout_declaration272 inout_declaration_instance272();
    inout_declaration273 inout_declaration_instance273();
    inout_declaration274 inout_declaration_instance274();
    inout_declaration275 inout_declaration_instance275();
    inout_declaration276 inout_declaration_instance276();
    inout_declaration277 inout_declaration_instance277();
    inout_declaration278 inout_declaration_instance278();
    inout_declaration279 inout_declaration_instance279();
    inout_declaration280 inout_declaration_instance280();
    inout_declaration281 inout_declaration_instance281();
    inout_declaration282 inout_declaration_instance282();
    inout_declaration283 inout_declaration_instance283();
    inout_declaration284 inout_declaration_instance284();
    inout_declaration285 inout_declaration_instance285();
    inout_declaration286 inout_declaration_instance286();
    inout_declaration287 inout_declaration_instance287();
    inout_declaration288 inout_declaration_instance288();
    inout_declaration289 inout_declaration_instance289();
    inout_declaration290 inout_declaration_instance290();
    inout_declaration291 inout_declaration_instance291();
    inout_declaration292 inout_declaration_instance292();
    inout_declaration293 inout_declaration_instance293();
    inout_declaration294 inout_declaration_instance294();
    inout_declaration295 inout_declaration_instance295();
    inout_declaration296 inout_declaration_instance296();
    inout_declaration297 inout_declaration_instance297();
    inout_declaration298 inout_declaration_instance298();
    inout_declaration299 inout_declaration_instance299();
    inout_declaration300 inout_declaration_instance300();
    inout_declaration301 inout_declaration_instance301();
    inout_declaration302 inout_declaration_instance302();
    inout_declaration303 inout_declaration_instance303();
    inout_declaration304 inout_declaration_instance304();
    inout_declaration305 inout_declaration_instance305();
    inout_declaration306 inout_declaration_instance306();
    inout_declaration307 inout_declaration_instance307();
    inout_declaration308 inout_declaration_instance308();
    inout_declaration309 inout_declaration_instance309();
    inout_declaration310 inout_declaration_instance310();
    inout_declaration311 inout_declaration_instance311();
    inout_declaration312 inout_declaration_instance312();
    inout_declaration313 inout_declaration_instance313();
    inout_declaration314 inout_declaration_instance314();
    inout_declaration315 inout_declaration_instance315();
    inout_declaration316 inout_declaration_instance316();
    inout_declaration317 inout_declaration_instance317();
    inout_declaration318 inout_declaration_instance318();
    inout_declaration319 inout_declaration_instance319();
    inout_declaration320 inout_declaration_instance320();
    inout_declaration321 inout_declaration_instance321();
    inout_declaration322 inout_declaration_instance322();
    inout_declaration323 inout_declaration_instance323();
    inout_declaration324 inout_declaration_instance324();
    inout_declaration325 inout_declaration_instance325();
    inout_declaration326 inout_declaration_instance326();
    inout_declaration327 inout_declaration_instance327();
    inout_declaration328 inout_declaration_instance328();
    inout_declaration329 inout_declaration_instance329();
    inout_declaration330 inout_declaration_instance330();
    inout_declaration331 inout_declaration_instance331();
    inout_declaration332 inout_declaration_instance332();
    inout_declaration333 inout_declaration_instance333();
    inout_declaration334 inout_declaration_instance334();
    inout_declaration335 inout_declaration_instance335();
    inout_declaration336 inout_declaration_instance336();
    inout_declaration337 inout_declaration_instance337();
    inout_declaration338 inout_declaration_instance338();
    inout_declaration339 inout_declaration_instance339();
    inout_declaration340 inout_declaration_instance340();
    inout_declaration341 inout_declaration_instance341();
    inout_declaration342 inout_declaration_instance342();
    inout_declaration343 inout_declaration_instance343();
    inout_declaration344 inout_declaration_instance344();
    inout_declaration345 inout_declaration_instance345();
    inout_declaration346 inout_declaration_instance346();
    inout_declaration347 inout_declaration_instance347();
    inout_declaration348 inout_declaration_instance348();
    inout_declaration349 inout_declaration_instance349();
    inout_declaration350 inout_declaration_instance350();
    inout_declaration351 inout_declaration_instance351();
    inout_declaration352 inout_declaration_instance352();
    inout_declaration353 inout_declaration_instance353();
    inout_declaration354 inout_declaration_instance354();
    inout_declaration355 inout_declaration_instance355();
    inout_declaration356 inout_declaration_instance356();
    inout_declaration357 inout_declaration_instance357();
    inout_declaration358 inout_declaration_instance358();
    inout_declaration359 inout_declaration_instance359();
    inout_declaration360 inout_declaration_instance360();
    inout_declaration361 inout_declaration_instance361();
    inout_declaration362 inout_declaration_instance362();
    inout_declaration363 inout_declaration_instance363();
    inout_declaration364 inout_declaration_instance364();
    inout_declaration365 inout_declaration_instance365();
    inout_declaration366 inout_declaration_instance366();
    inout_declaration367 inout_declaration_instance367();
    inout_declaration368 inout_declaration_instance368();
    inout_declaration369 inout_declaration_instance369();
    inout_declaration370 inout_declaration_instance370();
    inout_declaration371 inout_declaration_instance371();
    inout_declaration372 inout_declaration_instance372();
    inout_declaration373 inout_declaration_instance373();
    inout_declaration374 inout_declaration_instance374();
    inout_declaration375 inout_declaration_instance375();
    inout_declaration376 inout_declaration_instance376();
    inout_declaration377 inout_declaration_instance377();
    inout_declaration378 inout_declaration_instance378();
    inout_declaration379 inout_declaration_instance379();
    inout_declaration380 inout_declaration_instance380();
    inout_declaration381 inout_declaration_instance381();
    inout_declaration382 inout_declaration_instance382();
    inout_declaration383 inout_declaration_instance383();
    inout_declaration384 inout_declaration_instance384();
    inout_declaration385 inout_declaration_instance385();
    inout_declaration386 inout_declaration_instance386();
    inout_declaration387 inout_declaration_instance387();
    inout_declaration388 inout_declaration_instance388();
    inout_declaration389 inout_declaration_instance389();
    inout_declaration390 inout_declaration_instance390();
    inout_declaration391 inout_declaration_instance391();
    inout_declaration392 inout_declaration_instance392();
    inout_declaration393 inout_declaration_instance393();
    inout_declaration394 inout_declaration_instance394();
    inout_declaration395 inout_declaration_instance395();
    inout_declaration396 inout_declaration_instance396();
    inout_declaration397 inout_declaration_instance397();
    inout_declaration398 inout_declaration_instance398();
    inout_declaration399 inout_declaration_instance399();
    inout_declaration400 inout_declaration_instance400();
    inout_declaration401 inout_declaration_instance401();
    inout_declaration402 inout_declaration_instance402();
    inout_declaration403 inout_declaration_instance403();
    inout_declaration404 inout_declaration_instance404();
    inout_declaration405 inout_declaration_instance405();
    inout_declaration406 inout_declaration_instance406();
    inout_declaration407 inout_declaration_instance407();
    inout_declaration408 inout_declaration_instance408();
    inout_declaration409 inout_declaration_instance409();
    inout_declaration410 inout_declaration_instance410();
    inout_declaration411 inout_declaration_instance411();
    inout_declaration412 inout_declaration_instance412();
    inout_declaration413 inout_declaration_instance413();
    inout_declaration414 inout_declaration_instance414();
    inout_declaration415 inout_declaration_instance415();
    inout_declaration416 inout_declaration_instance416();
    inout_declaration417 inout_declaration_instance417();
    inout_declaration418 inout_declaration_instance418();
    inout_declaration419 inout_declaration_instance419();
    inout_declaration420 inout_declaration_instance420();
    inout_declaration421 inout_declaration_instance421();
    inout_declaration422 inout_declaration_instance422();
    inout_declaration423 inout_declaration_instance423();
    inout_declaration424 inout_declaration_instance424();
    inout_declaration425 inout_declaration_instance425();
    inout_declaration426 inout_declaration_instance426();
    inout_declaration427 inout_declaration_instance427();
    inout_declaration428 inout_declaration_instance428();
    inout_declaration429 inout_declaration_instance429();
    inout_declaration430 inout_declaration_instance430();
    inout_declaration431 inout_declaration_instance431();
    inout_declaration432 inout_declaration_instance432();
    inout_declaration433 inout_declaration_instance433();
    inout_declaration434 inout_declaration_instance434();
    inout_declaration435 inout_declaration_instance435();
    inout_declaration436 inout_declaration_instance436();
    inout_declaration437 inout_declaration_instance437();
    inout_declaration438 inout_declaration_instance438();
    inout_declaration439 inout_declaration_instance439();
    inout_declaration440 inout_declaration_instance440();
    inout_declaration441 inout_declaration_instance441();
    inout_declaration442 inout_declaration_instance442();
    inout_declaration443 inout_declaration_instance443();
    inout_declaration444 inout_declaration_instance444();
    inout_declaration445 inout_declaration_instance445();
    inout_declaration446 inout_declaration_instance446();
    inout_declaration447 inout_declaration_instance447();
    inout_declaration448 inout_declaration_instance448();
    inout_declaration449 inout_declaration_instance449();
    inout_declaration450 inout_declaration_instance450();
    inout_declaration451 inout_declaration_instance451();
    inout_declaration452 inout_declaration_instance452();
    inout_declaration453 inout_declaration_instance453();
    inout_declaration454 inout_declaration_instance454();
    inout_declaration455 inout_declaration_instance455();
    inout_declaration456 inout_declaration_instance456();
    inout_declaration457 inout_declaration_instance457();
    inout_declaration458 inout_declaration_instance458();
    inout_declaration459 inout_declaration_instance459();
    inout_declaration460 inout_declaration_instance460();
    inout_declaration461 inout_declaration_instance461();
    inout_declaration462 inout_declaration_instance462();
    inout_declaration463 inout_declaration_instance463();
    inout_declaration464 inout_declaration_instance464();
    inout_declaration465 inout_declaration_instance465();
    inout_declaration466 inout_declaration_instance466();
    inout_declaration467 inout_declaration_instance467();
    inout_declaration468 inout_declaration_instance468();
    inout_declaration469 inout_declaration_instance469();
    inout_declaration470 inout_declaration_instance470();
    inout_declaration471 inout_declaration_instance471();
    inout_declaration472 inout_declaration_instance472();
    inout_declaration473 inout_declaration_instance473();
    inout_declaration474 inout_declaration_instance474();
    inout_declaration475 inout_declaration_instance475();
    inout_declaration476 inout_declaration_instance476();
    inout_declaration477 inout_declaration_instance477();
    inout_declaration478 inout_declaration_instance478();
    inout_declaration479 inout_declaration_instance479();
    inout_declaration480 inout_declaration_instance480();
    inout_declaration481 inout_declaration_instance481();
    inout_declaration482 inout_declaration_instance482();
    inout_declaration483 inout_declaration_instance483();
    inout_declaration484 inout_declaration_instance484();
    inout_declaration485 inout_declaration_instance485();
    inout_declaration486 inout_declaration_instance486();
    inout_declaration487 inout_declaration_instance487();
    inout_declaration488 inout_declaration_instance488();
    inout_declaration489 inout_declaration_instance489();
    inout_declaration490 inout_declaration_instance490();
    inout_declaration491 inout_declaration_instance491();
    inout_declaration492 inout_declaration_instance492();
    inout_declaration493 inout_declaration_instance493();
    inout_declaration494 inout_declaration_instance494();
    inout_declaration495 inout_declaration_instance495();
    inout_declaration496 inout_declaration_instance496();
    inout_declaration497 inout_declaration_instance497();
    inout_declaration498 inout_declaration_instance498();
    inout_declaration499 inout_declaration_instance499();
    inout_declaration500 inout_declaration_instance500();
    inout_declaration501 inout_declaration_instance501();
    inout_declaration502 inout_declaration_instance502();
    inout_declaration503 inout_declaration_instance503();
    inout_declaration504 inout_declaration_instance504();
    inout_declaration505 inout_declaration_instance505();
    inout_declaration506 inout_declaration_instance506();
    inout_declaration507 inout_declaration_instance507();
    inout_declaration508 inout_declaration_instance508();
    inout_declaration509 inout_declaration_instance509();
    inout_declaration510 inout_declaration_instance510();
    inout_declaration511 inout_declaration_instance511();
    inout_declaration512 inout_declaration_instance512();
    inout_declaration513 inout_declaration_instance513();
    inout_declaration514 inout_declaration_instance514();
    inout_declaration515 inout_declaration_instance515();
    inout_declaration516 inout_declaration_instance516();
    inout_declaration517 inout_declaration_instance517();
    inout_declaration518 inout_declaration_instance518();
    inout_declaration519 inout_declaration_instance519();
    inout_declaration520 inout_declaration_instance520();
    inout_declaration521 inout_declaration_instance521();
    inout_declaration522 inout_declaration_instance522();
    inout_declaration523 inout_declaration_instance523();
    inout_declaration524 inout_declaration_instance524();
    inout_declaration525 inout_declaration_instance525();
    inout_declaration526 inout_declaration_instance526();
    inout_declaration527 inout_declaration_instance527();
    inout_declaration528 inout_declaration_instance528();
    inout_declaration529 inout_declaration_instance529();
    inout_declaration530 inout_declaration_instance530();
    inout_declaration531 inout_declaration_instance531();
    inout_declaration532 inout_declaration_instance532();
    inout_declaration533 inout_declaration_instance533();
    inout_declaration534 inout_declaration_instance534();
    inout_declaration535 inout_declaration_instance535();
    inout_declaration536 inout_declaration_instance536();
    inout_declaration537 inout_declaration_instance537();
    inout_declaration538 inout_declaration_instance538();
    inout_declaration539 inout_declaration_instance539();
    inout_declaration540 inout_declaration_instance540();
    inout_declaration541 inout_declaration_instance541();
    inout_declaration542 inout_declaration_instance542();
    inout_declaration543 inout_declaration_instance543();
    inout_declaration544 inout_declaration_instance544();
    inout_declaration545 inout_declaration_instance545();
    inout_declaration546 inout_declaration_instance546();
    inout_declaration547 inout_declaration_instance547();
    inout_declaration548 inout_declaration_instance548();
    inout_declaration549 inout_declaration_instance549();
    inout_declaration550 inout_declaration_instance550();
    inout_declaration551 inout_declaration_instance551();
    inout_declaration552 inout_declaration_instance552();
    inout_declaration553 inout_declaration_instance553();
    inout_declaration554 inout_declaration_instance554();
    inout_declaration555 inout_declaration_instance555();
    inout_declaration556 inout_declaration_instance556();
    inout_declaration557 inout_declaration_instance557();
    inout_declaration558 inout_declaration_instance558();
    inout_declaration559 inout_declaration_instance559();
    inout_declaration560 inout_declaration_instance560();
    inout_declaration561 inout_declaration_instance561();
    inout_declaration562 inout_declaration_instance562();
    inout_declaration563 inout_declaration_instance563();
    inout_declaration564 inout_declaration_instance564();
    inout_declaration565 inout_declaration_instance565();
    inout_declaration566 inout_declaration_instance566();
    inout_declaration567 inout_declaration_instance567();
    inout_declaration568 inout_declaration_instance568();
    inout_declaration569 inout_declaration_instance569();
    inout_declaration570 inout_declaration_instance570();
    inout_declaration571 inout_declaration_instance571();
endmodule
//@
//author : andreib
module inout_declaration0( abc,ABC ); inout abc,ABC;
endmodule
//author : andreib
module inout_declaration1( abc,ABC ); inout [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration2( abc,ABC ); inout [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration3( abc,ABC ); inout [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration4( abc,ABC ); inout [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration5( abc,ABC ); inout [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration6( abc,ABC ); inout [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration7( abc,ABC ); inout [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration8( abc,ABC ); inout [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration9( abc,ABC ); inout [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration10( abc,ABC ); inout [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration11( abc,ABC ); inout [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration12( abc,ABC ); inout [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration13( abc,ABC ); inout [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration14( abc,ABC ); inout [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration15( abc,ABC ); inout [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration16( abc,ABC ); inout [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration17( abc,ABC ); inout [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration18( abc,ABC ); inout [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration19( abc,ABC ); inout [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration20( abc,ABC ); inout [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration21( abc,ABC ); inout [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration22( abc,ABC ); inout [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration23( abc,ABC ); inout [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration24( abc,ABC ); inout [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration25( abc,ABC ); inout [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration26( abc,ABC ); inout signed abc,ABC;
endmodule
//author : andreib
module inout_declaration27( abc,ABC ); inout signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration28( abc,ABC ); inout signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration29( abc,ABC ); inout signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration30( abc,ABC ); inout signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration31( abc,ABC ); inout signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration32( abc,ABC ); inout signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration33( abc,ABC ); inout signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration34( abc,ABC ); inout signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration35( abc,ABC ); inout signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration36( abc,ABC ); inout signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration37( abc,ABC ); inout signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration38( abc,ABC ); inout signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration39( abc,ABC ); inout signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration40( abc,ABC ); inout signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration41( abc,ABC ); inout signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration42( abc,ABC ); inout signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration43( abc,ABC ); inout signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration44( abc,ABC ); inout signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration45( abc,ABC ); inout signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration46( abc,ABC ); inout signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration47( abc,ABC ); inout signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration48( abc,ABC ); inout signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration49( abc,ABC ); inout signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration50( abc,ABC ); inout signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration51( abc,ABC ); inout signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration52( abc,ABC ); inout supply0 abc,ABC;
endmodule
//author : andreib
module inout_declaration53( abc,ABC ); inout supply0 [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration54( abc,ABC ); inout supply0 [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration55( abc,ABC ); inout supply0 [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration56( abc,ABC ); inout supply0 [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration57( abc,ABC ); inout supply0 [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration58( abc,ABC ); inout supply0 [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration59( abc,ABC ); inout supply0 [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration60( abc,ABC ); inout supply0 [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration61( abc,ABC ); inout supply0 [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration62( abc,ABC ); inout supply0 [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration63( abc,ABC ); inout supply0 [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration64( abc,ABC ); inout supply0 [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration65( abc,ABC ); inout supply0 [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration66( abc,ABC ); inout supply0 [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration67( abc,ABC ); inout supply0 [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration68( abc,ABC ); inout supply0 [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration69( abc,ABC ); inout supply0 [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration70( abc,ABC ); inout supply0 [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration71( abc,ABC ); inout supply0 [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration72( abc,ABC ); inout supply0 [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration73( abc,ABC ); inout supply0 [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration74( abc,ABC ); inout supply0 [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration75( abc,ABC ); inout supply0 [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration76( abc,ABC ); inout supply0 [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration77( abc,ABC ); inout supply0 [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration78( abc,ABC ); inout supply0 signed abc,ABC;
endmodule
//author : andreib
module inout_declaration79( abc,ABC ); inout supply0 signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration80( abc,ABC ); inout supply0 signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration81( abc,ABC ); inout supply0 signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration82( abc,ABC ); inout supply0 signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration83( abc,ABC ); inout supply0 signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration84( abc,ABC ); inout supply0 signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration85( abc,ABC ); inout supply0 signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration86( abc,ABC ); inout supply0 signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration87( abc,ABC ); inout supply0 signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration88( abc,ABC ); inout supply0 signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration89( abc,ABC ); inout supply0 signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration90( abc,ABC ); inout supply0 signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration91( abc,ABC ); inout supply0 signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration92( abc,ABC ); inout supply0 signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration93( abc,ABC ); inout supply0 signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration94( abc,ABC ); inout supply0 signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration95( abc,ABC ); inout supply0 signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration96( abc,ABC ); inout supply0 signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration97( abc,ABC ); inout supply0 signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration98( abc,ABC ); inout supply0 signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration99( abc,ABC ); inout supply0 signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration100( abc,ABC ); inout supply0 signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration101( abc,ABC ); inout supply0 signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration102( abc,ABC ); inout supply0 signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration103( abc,ABC ); inout supply0 signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration104( abc,ABC ); inout supply1 abc,ABC;
endmodule
//author : andreib
module inout_declaration105( abc,ABC ); inout supply1 [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration106( abc,ABC ); inout supply1 [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration107( abc,ABC ); inout supply1 [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration108( abc,ABC ); inout supply1 [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration109( abc,ABC ); inout supply1 [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration110( abc,ABC ); inout supply1 [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration111( abc,ABC ); inout supply1 [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration112( abc,ABC ); inout supply1 [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration113( abc,ABC ); inout supply1 [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration114( abc,ABC ); inout supply1 [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration115( abc,ABC ); inout supply1 [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration116( abc,ABC ); inout supply1 [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration117( abc,ABC ); inout supply1 [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration118( abc,ABC ); inout supply1 [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration119( abc,ABC ); inout supply1 [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration120( abc,ABC ); inout supply1 [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration121( abc,ABC ); inout supply1 [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration122( abc,ABC ); inout supply1 [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration123( abc,ABC ); inout supply1 [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration124( abc,ABC ); inout supply1 [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration125( abc,ABC ); inout supply1 [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration126( abc,ABC ); inout supply1 [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration127( abc,ABC ); inout supply1 [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration128( abc,ABC ); inout supply1 [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration129( abc,ABC ); inout supply1 [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration130( abc,ABC ); inout supply1 signed abc,ABC;
endmodule
//author : andreib
module inout_declaration131( abc,ABC ); inout supply1 signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration132( abc,ABC ); inout supply1 signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration133( abc,ABC ); inout supply1 signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration134( abc,ABC ); inout supply1 signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration135( abc,ABC ); inout supply1 signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration136( abc,ABC ); inout supply1 signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration137( abc,ABC ); inout supply1 signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration138( abc,ABC ); inout supply1 signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration139( abc,ABC ); inout supply1 signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration140( abc,ABC ); inout supply1 signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration141( abc,ABC ); inout supply1 signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration142( abc,ABC ); inout supply1 signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration143( abc,ABC ); inout supply1 signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration144( abc,ABC ); inout supply1 signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration145( abc,ABC ); inout supply1 signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration146( abc,ABC ); inout supply1 signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration147( abc,ABC ); inout supply1 signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration148( abc,ABC ); inout supply1 signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration149( abc,ABC ); inout supply1 signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration150( abc,ABC ); inout supply1 signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration151( abc,ABC ); inout supply1 signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration152( abc,ABC ); inout supply1 signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration153( abc,ABC ); inout supply1 signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration154( abc,ABC ); inout supply1 signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration155( abc,ABC ); inout supply1 signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration156( abc,ABC ); inout tri abc,ABC;
endmodule
//author : andreib
module inout_declaration157( abc,ABC ); inout tri [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration158( abc,ABC ); inout tri [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration159( abc,ABC ); inout tri [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration160( abc,ABC ); inout tri [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration161( abc,ABC ); inout tri [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration162( abc,ABC ); inout tri [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration163( abc,ABC ); inout tri [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration164( abc,ABC ); inout tri [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration165( abc,ABC ); inout tri [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration166( abc,ABC ); inout tri [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration167( abc,ABC ); inout tri [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration168( abc,ABC ); inout tri [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration169( abc,ABC ); inout tri [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration170( abc,ABC ); inout tri [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration171( abc,ABC ); inout tri [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration172( abc,ABC ); inout tri [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration173( abc,ABC ); inout tri [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration174( abc,ABC ); inout tri [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration175( abc,ABC ); inout tri [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration176( abc,ABC ); inout tri [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration177( abc,ABC ); inout tri [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration178( abc,ABC ); inout tri [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration179( abc,ABC ); inout tri [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration180( abc,ABC ); inout tri [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration181( abc,ABC ); inout tri [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration182( abc,ABC ); inout tri signed abc,ABC;
endmodule
//author : andreib
module inout_declaration183( abc,ABC ); inout tri signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration184( abc,ABC ); inout tri signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration185( abc,ABC ); inout tri signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration186( abc,ABC ); inout tri signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration187( abc,ABC ); inout tri signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration188( abc,ABC ); inout tri signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration189( abc,ABC ); inout tri signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration190( abc,ABC ); inout tri signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration191( abc,ABC ); inout tri signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration192( abc,ABC ); inout tri signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration193( abc,ABC ); inout tri signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration194( abc,ABC ); inout tri signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration195( abc,ABC ); inout tri signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration196( abc,ABC ); inout tri signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration197( abc,ABC ); inout tri signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration198( abc,ABC ); inout tri signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration199( abc,ABC ); inout tri signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration200( abc,ABC ); inout tri signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration201( abc,ABC ); inout tri signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration202( abc,ABC ); inout tri signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration203( abc,ABC ); inout tri signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration204( abc,ABC ); inout tri signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration205( abc,ABC ); inout tri signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration206( abc,ABC ); inout tri signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration207( abc,ABC ); inout tri signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration208( abc,ABC ); inout triand abc,ABC;
endmodule
//author : andreib
module inout_declaration209( abc,ABC ); inout triand [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration210( abc,ABC ); inout triand [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration211( abc,ABC ); inout triand [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration212( abc,ABC ); inout triand [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration213( abc,ABC ); inout triand [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration214( abc,ABC ); inout triand [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration215( abc,ABC ); inout triand [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration216( abc,ABC ); inout triand [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration217( abc,ABC ); inout triand [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration218( abc,ABC ); inout triand [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration219( abc,ABC ); inout triand [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration220( abc,ABC ); inout triand [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration221( abc,ABC ); inout triand [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration222( abc,ABC ); inout triand [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration223( abc,ABC ); inout triand [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration224( abc,ABC ); inout triand [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration225( abc,ABC ); inout triand [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration226( abc,ABC ); inout triand [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration227( abc,ABC ); inout triand [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration228( abc,ABC ); inout triand [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration229( abc,ABC ); inout triand [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration230( abc,ABC ); inout triand [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration231( abc,ABC ); inout triand [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration232( abc,ABC ); inout triand [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration233( abc,ABC ); inout triand [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration234( abc,ABC ); inout triand signed abc,ABC;
endmodule
//author : andreib
module inout_declaration235( abc,ABC ); inout triand signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration236( abc,ABC ); inout triand signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration237( abc,ABC ); inout triand signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration238( abc,ABC ); inout triand signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration239( abc,ABC ); inout triand signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration240( abc,ABC ); inout triand signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration241( abc,ABC ); inout triand signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration242( abc,ABC ); inout triand signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration243( abc,ABC ); inout triand signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration244( abc,ABC ); inout triand signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration245( abc,ABC ); inout triand signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration246( abc,ABC ); inout triand signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration247( abc,ABC ); inout triand signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration248( abc,ABC ); inout triand signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration249( abc,ABC ); inout triand signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration250( abc,ABC ); inout triand signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration251( abc,ABC ); inout triand signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration252( abc,ABC ); inout triand signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration253( abc,ABC ); inout triand signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration254( abc,ABC ); inout triand signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration255( abc,ABC ); inout triand signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration256( abc,ABC ); inout triand signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration257( abc,ABC ); inout triand signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration258( abc,ABC ); inout triand signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration259( abc,ABC ); inout triand signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration260( abc,ABC ); inout trior abc,ABC;
endmodule
//author : andreib
module inout_declaration261( abc,ABC ); inout trior [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration262( abc,ABC ); inout trior [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration263( abc,ABC ); inout trior [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration264( abc,ABC ); inout trior [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration265( abc,ABC ); inout trior [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration266( abc,ABC ); inout trior [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration267( abc,ABC ); inout trior [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration268( abc,ABC ); inout trior [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration269( abc,ABC ); inout trior [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration270( abc,ABC ); inout trior [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration271( abc,ABC ); inout trior [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration272( abc,ABC ); inout trior [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration273( abc,ABC ); inout trior [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration274( abc,ABC ); inout trior [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration275( abc,ABC ); inout trior [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration276( abc,ABC ); inout trior [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration277( abc,ABC ); inout trior [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration278( abc,ABC ); inout trior [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration279( abc,ABC ); inout trior [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration280( abc,ABC ); inout trior [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration281( abc,ABC ); inout trior [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration282( abc,ABC ); inout trior [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration283( abc,ABC ); inout trior [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration284( abc,ABC ); inout trior [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration285( abc,ABC ); inout trior [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration286( abc,ABC ); inout trior signed abc,ABC;
endmodule
//author : andreib
module inout_declaration287( abc,ABC ); inout trior signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration288( abc,ABC ); inout trior signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration289( abc,ABC ); inout trior signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration290( abc,ABC ); inout trior signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration291( abc,ABC ); inout trior signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration292( abc,ABC ); inout trior signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration293( abc,ABC ); inout trior signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration294( abc,ABC ); inout trior signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration295( abc,ABC ); inout trior signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration296( abc,ABC ); inout trior signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration297( abc,ABC ); inout trior signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration298( abc,ABC ); inout trior signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration299( abc,ABC ); inout trior signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration300( abc,ABC ); inout trior signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration301( abc,ABC ); inout trior signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration302( abc,ABC ); inout trior signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration303( abc,ABC ); inout trior signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration304( abc,ABC ); inout trior signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration305( abc,ABC ); inout trior signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration306( abc,ABC ); inout trior signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration307( abc,ABC ); inout trior signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration308( abc,ABC ); inout trior signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration309( abc,ABC ); inout trior signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration310( abc,ABC ); inout trior signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration311( abc,ABC ); inout trior signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration312( abc,ABC ); inout tri0 abc,ABC;
endmodule
//author : andreib
module inout_declaration313( abc,ABC ); inout tri0 [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration314( abc,ABC ); inout tri0 [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration315( abc,ABC ); inout tri0 [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration316( abc,ABC ); inout tri0 [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration317( abc,ABC ); inout tri0 [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration318( abc,ABC ); inout tri0 [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration319( abc,ABC ); inout tri0 [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration320( abc,ABC ); inout tri0 [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration321( abc,ABC ); inout tri0 [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration322( abc,ABC ); inout tri0 [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration323( abc,ABC ); inout tri0 [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration324( abc,ABC ); inout tri0 [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration325( abc,ABC ); inout tri0 [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration326( abc,ABC ); inout tri0 [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration327( abc,ABC ); inout tri0 [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration328( abc,ABC ); inout tri0 [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration329( abc,ABC ); inout tri0 [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration330( abc,ABC ); inout tri0 [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration331( abc,ABC ); inout tri0 [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration332( abc,ABC ); inout tri0 [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration333( abc,ABC ); inout tri0 [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration334( abc,ABC ); inout tri0 [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration335( abc,ABC ); inout tri0 [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration336( abc,ABC ); inout tri0 [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration337( abc,ABC ); inout tri0 [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration338( abc,ABC ); inout tri0 signed abc,ABC;
endmodule
//author : andreib
module inout_declaration339( abc,ABC ); inout tri0 signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration340( abc,ABC ); inout tri0 signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration341( abc,ABC ); inout tri0 signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration342( abc,ABC ); inout tri0 signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration343( abc,ABC ); inout tri0 signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration344( abc,ABC ); inout tri0 signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration345( abc,ABC ); inout tri0 signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration346( abc,ABC ); inout tri0 signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration347( abc,ABC ); inout tri0 signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration348( abc,ABC ); inout tri0 signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration349( abc,ABC ); inout tri0 signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration350( abc,ABC ); inout tri0 signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration351( abc,ABC ); inout tri0 signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration352( abc,ABC ); inout tri0 signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration353( abc,ABC ); inout tri0 signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration354( abc,ABC ); inout tri0 signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration355( abc,ABC ); inout tri0 signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration356( abc,ABC ); inout tri0 signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration357( abc,ABC ); inout tri0 signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration358( abc,ABC ); inout tri0 signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration359( abc,ABC ); inout tri0 signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration360( abc,ABC ); inout tri0 signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration361( abc,ABC ); inout tri0 signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration362( abc,ABC ); inout tri0 signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration363( abc,ABC ); inout tri0 signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration364( abc,ABC ); inout tri1 abc,ABC;
endmodule
//author : andreib
module inout_declaration365( abc,ABC ); inout tri1 [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration366( abc,ABC ); inout tri1 [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration367( abc,ABC ); inout tri1 [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration368( abc,ABC ); inout tri1 [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration369( abc,ABC ); inout tri1 [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration370( abc,ABC ); inout tri1 [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration371( abc,ABC ); inout tri1 [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration372( abc,ABC ); inout tri1 [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration373( abc,ABC ); inout tri1 [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration374( abc,ABC ); inout tri1 [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration375( abc,ABC ); inout tri1 [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration376( abc,ABC ); inout tri1 [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration377( abc,ABC ); inout tri1 [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration378( abc,ABC ); inout tri1 [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration379( abc,ABC ); inout tri1 [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration380( abc,ABC ); inout tri1 [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration381( abc,ABC ); inout tri1 [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration382( abc,ABC ); inout tri1 [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration383( abc,ABC ); inout tri1 [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration384( abc,ABC ); inout tri1 [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration385( abc,ABC ); inout tri1 [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration386( abc,ABC ); inout tri1 [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration387( abc,ABC ); inout tri1 [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration388( abc,ABC ); inout tri1 [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration389( abc,ABC ); inout tri1 [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration390( abc,ABC ); inout tri1 signed abc,ABC;
endmodule
//author : andreib
module inout_declaration391( abc,ABC ); inout tri1 signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration392( abc,ABC ); inout tri1 signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration393( abc,ABC ); inout tri1 signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration394( abc,ABC ); inout tri1 signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration395( abc,ABC ); inout tri1 signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration396( abc,ABC ); inout tri1 signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration397( abc,ABC ); inout tri1 signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration398( abc,ABC ); inout tri1 signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration399( abc,ABC ); inout tri1 signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration400( abc,ABC ); inout tri1 signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration401( abc,ABC ); inout tri1 signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration402( abc,ABC ); inout tri1 signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration403( abc,ABC ); inout tri1 signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration404( abc,ABC ); inout tri1 signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration405( abc,ABC ); inout tri1 signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration406( abc,ABC ); inout tri1 signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration407( abc,ABC ); inout tri1 signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration408( abc,ABC ); inout tri1 signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration409( abc,ABC ); inout tri1 signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration410( abc,ABC ); inout tri1 signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration411( abc,ABC ); inout tri1 signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration412( abc,ABC ); inout tri1 signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration413( abc,ABC ); inout tri1 signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration414( abc,ABC ); inout tri1 signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration415( abc,ABC ); inout tri1 signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration416( abc,ABC ); inout wire abc,ABC;
endmodule
//author : andreib
module inout_declaration417( abc,ABC ); inout wire [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration418( abc,ABC ); inout wire [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration419( abc,ABC ); inout wire [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration420( abc,ABC ); inout wire [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration421( abc,ABC ); inout wire [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration422( abc,ABC ); inout wire [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration423( abc,ABC ); inout wire [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration424( abc,ABC ); inout wire [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration425( abc,ABC ); inout wire [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration426( abc,ABC ); inout wire [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration427( abc,ABC ); inout wire [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration428( abc,ABC ); inout wire [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration429( abc,ABC ); inout wire [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration430( abc,ABC ); inout wire [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration431( abc,ABC ); inout wire [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration432( abc,ABC ); inout wire [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration433( abc,ABC ); inout wire [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration434( abc,ABC ); inout wire [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration435( abc,ABC ); inout wire [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration436( abc,ABC ); inout wire [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration437( abc,ABC ); inout wire [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration438( abc,ABC ); inout wire [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration439( abc,ABC ); inout wire [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration440( abc,ABC ); inout wire [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration441( abc,ABC ); inout wire [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration442( abc,ABC ); inout wire signed abc,ABC;
endmodule
//author : andreib
module inout_declaration443( abc,ABC ); inout wire signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration444( abc,ABC ); inout wire signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration445( abc,ABC ); inout wire signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration446( abc,ABC ); inout wire signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration447( abc,ABC ); inout wire signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration448( abc,ABC ); inout wire signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration449( abc,ABC ); inout wire signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration450( abc,ABC ); inout wire signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration451( abc,ABC ); inout wire signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration452( abc,ABC ); inout wire signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration453( abc,ABC ); inout wire signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration454( abc,ABC ); inout wire signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration455( abc,ABC ); inout wire signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration456( abc,ABC ); inout wire signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration457( abc,ABC ); inout wire signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration458( abc,ABC ); inout wire signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration459( abc,ABC ); inout wire signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration460( abc,ABC ); inout wire signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration461( abc,ABC ); inout wire signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration462( abc,ABC ); inout wire signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration463( abc,ABC ); inout wire signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration464( abc,ABC ); inout wire signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration465( abc,ABC ); inout wire signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration466( abc,ABC ); inout wire signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration467( abc,ABC ); inout wire signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration468( abc,ABC ); inout wand abc,ABC;
endmodule
//author : andreib
module inout_declaration469( abc,ABC ); inout wand [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration470( abc,ABC ); inout wand [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration471( abc,ABC ); inout wand [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration472( abc,ABC ); inout wand [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration473( abc,ABC ); inout wand [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration474( abc,ABC ); inout wand [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration475( abc,ABC ); inout wand [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration476( abc,ABC ); inout wand [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration477( abc,ABC ); inout wand [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration478( abc,ABC ); inout wand [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration479( abc,ABC ); inout wand [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration480( abc,ABC ); inout wand [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration481( abc,ABC ); inout wand [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration482( abc,ABC ); inout wand [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration483( abc,ABC ); inout wand [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration484( abc,ABC ); inout wand [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration485( abc,ABC ); inout wand [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration486( abc,ABC ); inout wand [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration487( abc,ABC ); inout wand [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration488( abc,ABC ); inout wand [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration489( abc,ABC ); inout wand [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration490( abc,ABC ); inout wand [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration491( abc,ABC ); inout wand [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration492( abc,ABC ); inout wand [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration493( abc,ABC ); inout wand [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration494( abc,ABC ); inout wand signed abc,ABC;
endmodule
//author : andreib
module inout_declaration495( abc,ABC ); inout wand signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration496( abc,ABC ); inout wand signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration497( abc,ABC ); inout wand signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration498( abc,ABC ); inout wand signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration499( abc,ABC ); inout wand signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration500( abc,ABC ); inout wand signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration501( abc,ABC ); inout wand signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration502( abc,ABC ); inout wand signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration503( abc,ABC ); inout wand signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration504( abc,ABC ); inout wand signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration505( abc,ABC ); inout wand signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration506( abc,ABC ); inout wand signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration507( abc,ABC ); inout wand signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration508( abc,ABC ); inout wand signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration509( abc,ABC ); inout wand signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration510( abc,ABC ); inout wand signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration511( abc,ABC ); inout wand signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration512( abc,ABC ); inout wand signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration513( abc,ABC ); inout wand signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration514( abc,ABC ); inout wand signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration515( abc,ABC ); inout wand signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration516( abc,ABC ); inout wand signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration517( abc,ABC ); inout wand signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration518( abc,ABC ); inout wand signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration519( abc,ABC ); inout wand signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration520( abc,ABC ); inout wor abc,ABC;
endmodule
//author : andreib
module inout_declaration521( abc,ABC ); inout wor [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration522( abc,ABC ); inout wor [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration523( abc,ABC ); inout wor [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration524( abc,ABC ); inout wor [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration525( abc,ABC ); inout wor [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration526( abc,ABC ); inout wor [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration527( abc,ABC ); inout wor [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration528( abc,ABC ); inout wor [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration529( abc,ABC ); inout wor [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration530( abc,ABC ); inout wor [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration531( abc,ABC ); inout wor [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration532( abc,ABC ); inout wor [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration533( abc,ABC ); inout wor [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration534( abc,ABC ); inout wor [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration535( abc,ABC ); inout wor [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration536( abc,ABC ); inout wor [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration537( abc,ABC ); inout wor [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration538( abc,ABC ); inout wor [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration539( abc,ABC ); inout wor [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration540( abc,ABC ); inout wor [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration541( abc,ABC ); inout wor [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration542( abc,ABC ); inout wor [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration543( abc,ABC ); inout wor [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration544( abc,ABC ); inout wor [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration545( abc,ABC ); inout wor [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration546( abc,ABC ); inout wor signed abc,ABC;
endmodule
//author : andreib
module inout_declaration547( abc,ABC ); inout wor signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration548( abc,ABC ); inout wor signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration549( abc,ABC ); inout wor signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration550( abc,ABC ); inout wor signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration551( abc,ABC ); inout wor signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration552( abc,ABC ); inout wor signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration553( abc,ABC ); inout wor signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration554( abc,ABC ); inout wor signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration555( abc,ABC ); inout wor signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration556( abc,ABC ); inout wor signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration557( abc,ABC ); inout wor signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration558( abc,ABC ); inout wor signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration559( abc,ABC ); inout wor signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration560( abc,ABC ); inout wor signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration561( abc,ABC ); inout wor signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration562( abc,ABC ); inout wor signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration563( abc,ABC ); inout wor signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration564( abc,ABC ); inout wor signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration565( abc,ABC ); inout wor signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration566( abc,ABC ); inout wor signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module inout_declaration567( abc,ABC ); inout wor signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration568( abc,ABC ); inout wor signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration569( abc,ABC ); inout wor signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration570( abc,ABC ); inout wor signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module inout_declaration571( abc,ABC ); inout wor signed [ "str" : "str" ] abc,ABC;
endmodule
