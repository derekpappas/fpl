// Test type: Hex Numbers - x digit
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=12'h2xX;
endmodule
