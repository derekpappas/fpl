-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./msi_rx_cslc_generated/code/vhdl/mfd_sec.vhd
-- FILE GENERATED ON : Tue Jun 17 01:23:46 2008
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity \mfd_sec\ is
  port(\lbadummy3\ : in std_logic);
begin
end entity;

architecture \mfd_sec_logic\ of \mfd_sec\ is
end architecture;

