`include "defines.v"

module m1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 256
  output [1 - 1:0] ar_sa0_s10;
  l1 l10(.ar_sa0_s10(ar_sa0_s10));
  `include "m1.logic.vh"
endmodule

