//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : sd_flash.v
//FILE GENERATED ON : Tue Jun 17 01:23:46 2008

`include "defines.v"

module sd_flash(lbadummy3);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 20
  input lbadummy3;
  `include "sd_flash.logic.v"
endmodule

