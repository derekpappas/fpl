//test type : module_or_generate_item ::= module_or_generate_item_declaration (reg_declaration)
//vparser rule name : 
//author : Codrin
module test_0150;
 (* fsm_state *) reg [7:0] state1;
endmodule
