-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./u_mbist_cslc_generated/code/vhdl/u_cmp.vhd
-- FILE GENERATED ON : Wed Nov 18 19:49:32 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u_cmp\ is
  port(\ifc_op_cmp_op1\ : in csl_bit_vector(10#15# downto 10#0#);
       \ifc_op_cmp_op2\ : in csl_bit_vector(10#15# downto 10#0#);
       \res\ : out csl_bit);
begin
end entity;

architecture \u_cmp_logic\ of \u_cmp\ is
begin
end architecture;

