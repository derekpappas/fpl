//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC CSL COMPILER
//COPYRIGHT (c) 2005, 2006 FastpathLogic Inc

`define br 0
`define alu 1
`define mem 2
module enum_test();
endmodule

