// Dummy by Claudiu

module MUX4_32;
endmodule

module TRIBUF_32;
endmodule

module PHI1_LATCH_EN_32;
endmodule

module MUX2_32;
endmodule

module PHI1_LATCH_EN_30;
endmodule

module PHI2_LATCH_EN_30;
endmodule

module MUX3_30;
endmodule

module PHI2_LATCH_EN_32;
endmodule

module MUX3_32;
endmodule

module COMP_6;
endmodule

module ADD_6;
endmodule

module MUX2_6;
endmodule

module PHI1_LATCH_6;
endmodule

module PHI2_LATCH_6;
endmodule

module PHI2_LATCH_7;
endmodule

module MUX2_7;
endmodule

module PHI1_LATCH_EN_7;
endmodule

module PHI2_LATCH_EN_7;
endmodule


module PHI2_LATCH_26;
endmodule

module MUX2_26;
endmodule

module PHI1_LATCH_EN_26;
endmodule

module PHI2_LATCH_EN_26;
endmodule

module PHI2_LATCH_24;
endmodule

module MUX2_24;
endmodule

module PHI1_LATCH_EN_24;
endmodule

module PHI2_LATCH_EN_24;
endmodule

module ADD_30;
endmodule

module MUX2_30;
endmodule

module PHI1_LATCH_30;
endmodule

module MUX2_10;
endmodule

module MUX2_20;
endmodule

module PHI1_LATCH_20;
endmodule

module PHI2_LATCH_20;
endmodule

module PHI2_LATCH_EN_10;
endmodule

module PHI1_LATCH_10;
endmodule

module MUX5_30;
endmodule

module PHI2_LATCH_30;
endmodule
