-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./top_cslc_generated/code/vhdl/u21.vhd
-- FILE GENERATED ON : Tue Mar 10 20:48:07 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u21\ is
  port(\ifc_in1_pi1\ : in csl_bit_vector(10#2# - 10#1# downto 10#0#);
       \ifc_in1_pi2\ : in csl_bit_vector(10#4# - 10#1# downto 10#0#);
       \ifc_in1_pi3\ : in csl_bit);
begin
end entity;

architecture \u21_logic\ of \u21\ is
begin
end architecture;

