// Test type: net_assignment - string
// Vparser rule name:
// Author: andreib
module netasign9;
wire a;
assign a="test_string";
endmodule
