// Test type: seq_block - begin - end
// Vparser rule name:
// Author: andreib
module seq_block1;
initial begin end
endmodule
