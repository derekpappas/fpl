u.vhd
