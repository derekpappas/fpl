u12.vhd
u11.vhd
u21.vhd
ubc.vhd
uabc.vhd
utop.vhd
