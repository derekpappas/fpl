`include "defines.v"

module u();
// Location of source csl unit: file name = RISC_ISA.csl line number = 8
  `include "u.logic.v"
endmodule

