// Test type: always statement - system_task_enable - no attribute instance
// Vparser rule name:
// Author: andreib
module alwcon34;
reg a;
always a=$random;
endmodule
