// Test type: delay_or_event_control - delay_control - delay_value
// Vparser rule name:
// Author: andreib
module delay_or_event_control1;
reg a;
initial #10 a=1'b1;
endmodule
