`include "defines.v"

module n0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 95
  input [1 - 1:0] ar_sa0_s10;
  m0 m0(.ar_sa0_s10(ar_sa0_s10));
  `include "n0.logic.vh"
endmodule

