`include "defines.v"

module pcictrl();
// Location of source csl unit: file name = IPX2400.csl line number = 107
  `include "pcictrl.logic.v"
endmodule

