// Test type: Binary Numbers - signed base letter case variation
// Vparser rule name: Numbers
// Author: andreib
module binary_num;
wire a;
assign a=3'sB101;
endmodule
