//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : eth_tx.v
//FILE GENERATED ON : Tue Jun 17 01:23:46 2008

`include "defines.v"

module eth_tx();
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 46
  `include "eth_tx.logic.v"
endmodule

