  --THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
--COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
--OUTPUT FILE NAME  : a.vhd
--FILE GENERATED ON : Wed Jan 20 06:20:06 2010


library ieee ; 
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all; 
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;
 
use work.csl_util_package.all;

entity a is 

-- Location of source csl unit: file name = assign10.csl line number = 11
           <= (:);
     <= ;
end a ; 

 architecture  arch_a of a is 
 begin 

 end  arch_a ; 
