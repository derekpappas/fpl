//st2.vh