//test type : block_item_declaration ::= realtime list_of_block_variable_identifiers;
//vparser rule name : 
//author : Codrin
module test_0530;
  (* reset, start_timers, ends = 1 *)
  realtime regfile[1:64], rtime;
endmodule
