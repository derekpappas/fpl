// Test type: initial statement - nonblocking_assignment - no attribute instance
// Vparser rule name:
// Author: andreib
module initcon19;
reg [7:0]a;
initial a<=2;
endmodule
