`include "defines.v"

module h1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 226
  output [1 - 1:0] ar_sa0_s10;
  g1 g10(.ar_sa0_s10(ar_sa0_s10));
  `include "h1.logic.vh"
endmodule

