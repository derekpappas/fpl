// Test type: Constant Expression - primary - param
// Vparser rule name:
// Author: andreib
module constantexpression;
parameter test=1;
reg[test:0] a;
endmodule
