//rn_logic.vh
