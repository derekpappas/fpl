-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./utop_cslc_generated/code/vhdl/usu.vhd
-- FILE GENERATED ON : Sat Mar 14 18:38:34 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \usu\ is
  port(\ifcsu0_iin\ : in csl_bit_vector(10#16# - 10#1# downto 10#0#);
       \ifcsu0_iout\ : out csl_bit_vector(10#16# - 10#1# downto 10#0#));
begin
end entity;

architecture \usu_logic\ of \usu\ is
begin
end architecture;

