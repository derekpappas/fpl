// Test type: net_assignment - unary operator, no attribute instance
// Vparser rule name:
// Author: andreib
module netasign2;
wire a;
assign a=^2;
endmodule
