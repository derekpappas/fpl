//test type : hierarchical_identifier binary_operator_&& hierarchical_identifier
//vparser rule name : 
//author : Bogdan Mereghea
module binary_operator10;
    wire a, b, c;
    assign a = b && c;
endmodule
