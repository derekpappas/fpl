`include "defines.v"

module u2();
// Location of source csl unit: file name = ar16.csl line number = 39
  `include "u2.logic.v"
endmodule

