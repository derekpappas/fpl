`define MAX 200
//parameter r = 20;
module tets;
    `define MIN 100
    parameter p = 10;
endmodule