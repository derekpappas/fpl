// Test type: always statement - procedural_continuous_assign - no attribute instance
// Vparser rule name:
// Author: andreib
module alwcon25;
reg [7:0]a;
always 
assign a=2;
endmodule
