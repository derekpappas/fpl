-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./msi_rx_cslc_generated/code/vhdl/mfd_sec.vhd
-- FILE GENERATED ON : Thu Jun 19 15:32:42 2008
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \mfd_sec\ is
  port(\lbdummy3\ : in csl_bit);
begin
end entity;

architecture \mfd_sec_logic\ of \mfd_sec\ is
begin
end architecture;

