u.vhd
top1.vhd
