// Test type: Continuous assignment - sup1, h0 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous556;
wire a;
assign (supply1, highz0) a=1'b1;
endmodule
