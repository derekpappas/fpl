

module top();

a a();
b b();

endmodule