`include "defines.v"

module x0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 165
  input [1 - 1:0] ar_sa0_s10;
  w0 w0(.ar_sa0_s10(ar_sa0_s10));
  `include "x0.logic.vh"
endmodule

