u1.vhd
u2.vhd
top.vhd
top1.vhd
