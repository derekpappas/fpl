usb_tm_packetizer.vhd
usb_tm_dispatcher.vhd
fab.vhd
usb_transaction_mgr.vhd
usb_protocol_mgr.vhd
uart.vhd
uart_mgr.vhd
usb_phy.vhd
fifo_regs.vhd
fab_filter.vhd
RAM.vhd
i2c.vhd
avalon_bridge.vhd
f_core.vhd
