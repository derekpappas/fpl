module x;
   reg _389000_389000 ; 
   reg __389000_389000;
   reg _389001_389001 ; 
   reg __389001_389001;
   reg _389002_389002 ; 
   reg __389002_389002;
   reg _389003_389003 ; 
   reg __389003_389003;
   reg _389004_389004 ; 
   reg __389004_389004;
   reg _389005_389005 ; 
   reg __389005_389005;
   reg _389006_389006 ; 
   reg __389006_389006;
   reg _389007_389007 ; 
   reg __389007_389007;
   reg _389008_389008 ; 
   reg __389008_389008;
   reg _389009_389009 ; 
   reg __389009_389009;
   reg _389010_389010 ; 
   reg __389010_389010;
   reg _389011_389011 ; 
   reg __389011_389011;
   reg _389012_389012 ; 
   reg __389012_389012;
   reg _389013_389013 ; 
   reg __389013_389013;
   reg _389014_389014 ; 
   reg __389014_389014;
   reg _389015_389015 ; 
   reg __389015_389015;
   reg _389016_389016 ; 
   reg __389016_389016;
   reg _389017_389017 ; 
   reg __389017_389017;
   reg _389018_389018 ; 
   reg __389018_389018;
   reg _389019_389019 ; 
   reg __389019_389019;
   reg _389020_389020 ; 
   reg __389020_389020;
   reg _389021_389021 ; 
   reg __389021_389021;
   reg _389022_389022 ; 
   reg __389022_389022;
   reg _389023_389023 ; 
   reg __389023_389023;
   reg _389024_389024 ; 
   reg __389024_389024;
   reg _389025_389025 ; 
   reg __389025_389025;
   reg _389026_389026 ; 
   reg __389026_389026;
   reg _389027_389027 ; 
   reg __389027_389027;
   reg _389028_389028 ; 
   reg __389028_389028;
   reg _389029_389029 ; 
   reg __389029_389029;
   reg _389030_389030 ; 
   reg __389030_389030;
   reg _389031_389031 ; 
   reg __389031_389031;
   reg _389032_389032 ; 
   reg __389032_389032;
   reg _389033_389033 ; 
   reg __389033_389033;
   reg _389034_389034 ; 
   reg __389034_389034;
   reg _389035_389035 ; 
   reg __389035_389035;
   reg _389036_389036 ; 
   reg __389036_389036;
   reg _389037_389037 ; 
   reg __389037_389037;
   reg _389038_389038 ; 
   reg __389038_389038;
   reg _389039_389039 ; 
   reg __389039_389039;
   reg _389040_389040 ; 
   reg __389040_389040;
   reg _389041_389041 ; 
   reg __389041_389041;
   reg _389042_389042 ; 
   reg __389042_389042;
   reg _389043_389043 ; 
   reg __389043_389043;
   reg _389044_389044 ; 
   reg __389044_389044;
   reg _389045_389045 ; 
   reg __389045_389045;
   reg _389046_389046 ; 
   reg __389046_389046;
   reg _389047_389047 ; 
   reg __389047_389047;
   reg _389048_389048 ; 
   reg __389048_389048;
   reg _389049_389049 ; 
   reg __389049_389049;
   reg _389050_389050 ; 
   reg __389050_389050;
   reg _389051_389051 ; 
   reg __389051_389051;
   reg _389052_389052 ; 
   reg __389052_389052;
   reg _389053_389053 ; 
   reg __389053_389053;
   reg _389054_389054 ; 
   reg __389054_389054;
   reg _389055_389055 ; 
   reg __389055_389055;
   reg _389056_389056 ; 
   reg __389056_389056;
   reg _389057_389057 ; 
   reg __389057_389057;
   reg _389058_389058 ; 
   reg __389058_389058;
   reg _389059_389059 ; 
   reg __389059_389059;
   reg _389060_389060 ; 
   reg __389060_389060;
   reg _389061_389061 ; 
   reg __389061_389061;
   reg _389062_389062 ; 
   reg __389062_389062;
   reg _389063_389063 ; 
   reg __389063_389063;
   reg _389064_389064 ; 
   reg __389064_389064;
   reg _389065_389065 ; 
   reg __389065_389065;
   reg _389066_389066 ; 
   reg __389066_389066;
   reg _389067_389067 ; 
   reg __389067_389067;
   reg _389068_389068 ; 
   reg __389068_389068;
   reg _389069_389069 ; 
   reg __389069_389069;
   reg _389070_389070 ; 
   reg __389070_389070;
   reg _389071_389071 ; 
   reg __389071_389071;
   reg _389072_389072 ; 
   reg __389072_389072;
   reg _389073_389073 ; 
   reg __389073_389073;
   reg _389074_389074 ; 
   reg __389074_389074;
   reg _389075_389075 ; 
   reg __389075_389075;
   reg _389076_389076 ; 
   reg __389076_389076;
   reg _389077_389077 ; 
   reg __389077_389077;
   reg _389078_389078 ; 
   reg __389078_389078;
   reg _389079_389079 ; 
   reg __389079_389079;
   reg _389080_389080 ; 
   reg __389080_389080;
   reg _389081_389081 ; 
   reg __389081_389081;
   reg _389082_389082 ; 
   reg __389082_389082;
   reg _389083_389083 ; 
   reg __389083_389083;
   reg _389084_389084 ; 
   reg __389084_389084;
   reg _389085_389085 ; 
   reg __389085_389085;
   reg _389086_389086 ; 
   reg __389086_389086;
   reg _389087_389087 ; 
   reg __389087_389087;
   reg _389088_389088 ; 
   reg __389088_389088;
   reg _389089_389089 ; 
   reg __389089_389089;
   reg _389090_389090 ; 
   reg __389090_389090;
   reg _389091_389091 ; 
   reg __389091_389091;
   reg _389092_389092 ; 
   reg __389092_389092;
   reg _389093_389093 ; 
   reg __389093_389093;
   reg _389094_389094 ; 
   reg __389094_389094;
   reg _389095_389095 ; 
   reg __389095_389095;
   reg _389096_389096 ; 
   reg __389096_389096;
   reg _389097_389097 ; 
   reg __389097_389097;
   reg _389098_389098 ; 
   reg __389098_389098;
   reg _389099_389099 ; 
   reg __389099_389099;
   reg _389100_389100 ; 
   reg __389100_389100;
   reg _389101_389101 ; 
   reg __389101_389101;
   reg _389102_389102 ; 
   reg __389102_389102;
   reg _389103_389103 ; 
   reg __389103_389103;
   reg _389104_389104 ; 
   reg __389104_389104;
   reg _389105_389105 ; 
   reg __389105_389105;
   reg _389106_389106 ; 
   reg __389106_389106;
   reg _389107_389107 ; 
   reg __389107_389107;
   reg _389108_389108 ; 
   reg __389108_389108;
   reg _389109_389109 ; 
   reg __389109_389109;
   reg _389110_389110 ; 
   reg __389110_389110;
   reg _389111_389111 ; 
   reg __389111_389111;
   reg _389112_389112 ; 
   reg __389112_389112;
   reg _389113_389113 ; 
   reg __389113_389113;
   reg _389114_389114 ; 
   reg __389114_389114;
   reg _389115_389115 ; 
   reg __389115_389115;
   reg _389116_389116 ; 
   reg __389116_389116;
   reg _389117_389117 ; 
   reg __389117_389117;
   reg _389118_389118 ; 
   reg __389118_389118;
   reg _389119_389119 ; 
   reg __389119_389119;
   reg _389120_389120 ; 
   reg __389120_389120;
   reg _389121_389121 ; 
   reg __389121_389121;
   reg _389122_389122 ; 
   reg __389122_389122;
   reg _389123_389123 ; 
   reg __389123_389123;
   reg _389124_389124 ; 
   reg __389124_389124;
   reg _389125_389125 ; 
   reg __389125_389125;
   reg _389126_389126 ; 
   reg __389126_389126;
   reg _389127_389127 ; 
   reg __389127_389127;
   reg _389128_389128 ; 
   reg __389128_389128;
   reg _389129_389129 ; 
   reg __389129_389129;
   reg _389130_389130 ; 
   reg __389130_389130;
   reg _389131_389131 ; 
   reg __389131_389131;
   reg _389132_389132 ; 
   reg __389132_389132;
   reg _389133_389133 ; 
   reg __389133_389133;
   reg _389134_389134 ; 
   reg __389134_389134;
   reg _389135_389135 ; 
   reg __389135_389135;
   reg _389136_389136 ; 
   reg __389136_389136;
   reg _389137_389137 ; 
   reg __389137_389137;
   reg _389138_389138 ; 
   reg __389138_389138;
   reg _389139_389139 ; 
   reg __389139_389139;
   reg _389140_389140 ; 
   reg __389140_389140;
   reg _389141_389141 ; 
   reg __389141_389141;
   reg _389142_389142 ; 
   reg __389142_389142;
   reg _389143_389143 ; 
   reg __389143_389143;
   reg _389144_389144 ; 
   reg __389144_389144;
   reg _389145_389145 ; 
   reg __389145_389145;
   reg _389146_389146 ; 
   reg __389146_389146;
   reg _389147_389147 ; 
   reg __389147_389147;
   reg _389148_389148 ; 
   reg __389148_389148;
   reg _389149_389149 ; 
   reg __389149_389149;
   reg _389150_389150 ; 
   reg __389150_389150;
   reg _389151_389151 ; 
   reg __389151_389151;
   reg _389152_389152 ; 
   reg __389152_389152;
   reg _389153_389153 ; 
   reg __389153_389153;
   reg _389154_389154 ; 
   reg __389154_389154;
   reg _389155_389155 ; 
   reg __389155_389155;
   reg _389156_389156 ; 
   reg __389156_389156;
   reg _389157_389157 ; 
   reg __389157_389157;
   reg _389158_389158 ; 
   reg __389158_389158;
   reg _389159_389159 ; 
   reg __389159_389159;
   reg _389160_389160 ; 
   reg __389160_389160;
   reg _389161_389161 ; 
   reg __389161_389161;
   reg _389162_389162 ; 
   reg __389162_389162;
   reg _389163_389163 ; 
   reg __389163_389163;
   reg _389164_389164 ; 
   reg __389164_389164;
   reg _389165_389165 ; 
   reg __389165_389165;
   reg _389166_389166 ; 
   reg __389166_389166;
   reg _389167_389167 ; 
   reg __389167_389167;
   reg _389168_389168 ; 
   reg __389168_389168;
   reg _389169_389169 ; 
   reg __389169_389169;
   reg _389170_389170 ; 
   reg __389170_389170;
   reg _389171_389171 ; 
   reg __389171_389171;
   reg _389172_389172 ; 
   reg __389172_389172;
   reg _389173_389173 ; 
   reg __389173_389173;
   reg _389174_389174 ; 
   reg __389174_389174;
   reg _389175_389175 ; 
   reg __389175_389175;
   reg _389176_389176 ; 
   reg __389176_389176;
   reg _389177_389177 ; 
   reg __389177_389177;
   reg _389178_389178 ; 
   reg __389178_389178;
   reg _389179_389179 ; 
   reg __389179_389179;
   reg _389180_389180 ; 
   reg __389180_389180;
   reg _389181_389181 ; 
   reg __389181_389181;
   reg _389182_389182 ; 
   reg __389182_389182;
   reg _389183_389183 ; 
   reg __389183_389183;
   reg _389184_389184 ; 
   reg __389184_389184;
   reg _389185_389185 ; 
   reg __389185_389185;
   reg _389186_389186 ; 
   reg __389186_389186;
   reg _389187_389187 ; 
   reg __389187_389187;
   reg _389188_389188 ; 
   reg __389188_389188;
   reg _389189_389189 ; 
   reg __389189_389189;
   reg _389190_389190 ; 
   reg __389190_389190;
   reg _389191_389191 ; 
   reg __389191_389191;
   reg _389192_389192 ; 
   reg __389192_389192;
   reg _389193_389193 ; 
   reg __389193_389193;
   reg _389194_389194 ; 
   reg __389194_389194;
   reg _389195_389195 ; 
   reg __389195_389195;
   reg _389196_389196 ; 
   reg __389196_389196;
   reg _389197_389197 ; 
   reg __389197_389197;
   reg _389198_389198 ; 
   reg __389198_389198;
   reg _389199_389199 ; 
   reg __389199_389199;
   reg _389200_389200 ; 
   reg __389200_389200;
   reg _389201_389201 ; 
   reg __389201_389201;
   reg _389202_389202 ; 
   reg __389202_389202;
   reg _389203_389203 ; 
   reg __389203_389203;
   reg _389204_389204 ; 
   reg __389204_389204;
   reg _389205_389205 ; 
   reg __389205_389205;
   reg _389206_389206 ; 
   reg __389206_389206;
   reg _389207_389207 ; 
   reg __389207_389207;
   reg _389208_389208 ; 
   reg __389208_389208;
   reg _389209_389209 ; 
   reg __389209_389209;
   reg _389210_389210 ; 
   reg __389210_389210;
   reg _389211_389211 ; 
   reg __389211_389211;
   reg _389212_389212 ; 
   reg __389212_389212;
   reg _389213_389213 ; 
   reg __389213_389213;
   reg _389214_389214 ; 
   reg __389214_389214;
   reg _389215_389215 ; 
   reg __389215_389215;
   reg _389216_389216 ; 
   reg __389216_389216;
   reg _389217_389217 ; 
   reg __389217_389217;
   reg _389218_389218 ; 
   reg __389218_389218;
   reg _389219_389219 ; 
   reg __389219_389219;
   reg _389220_389220 ; 
   reg __389220_389220;
   reg _389221_389221 ; 
   reg __389221_389221;
   reg _389222_389222 ; 
   reg __389222_389222;
   reg _389223_389223 ; 
   reg __389223_389223;
   reg _389224_389224 ; 
   reg __389224_389224;
   reg _389225_389225 ; 
   reg __389225_389225;
   reg _389226_389226 ; 
   reg __389226_389226;
   reg _389227_389227 ; 
   reg __389227_389227;
   reg _389228_389228 ; 
   reg __389228_389228;
   reg _389229_389229 ; 
   reg __389229_389229;
   reg _389230_389230 ; 
   reg __389230_389230;
   reg _389231_389231 ; 
   reg __389231_389231;
   reg _389232_389232 ; 
   reg __389232_389232;
   reg _389233_389233 ; 
   reg __389233_389233;
   reg _389234_389234 ; 
   reg __389234_389234;
   reg _389235_389235 ; 
   reg __389235_389235;
   reg _389236_389236 ; 
   reg __389236_389236;
   reg _389237_389237 ; 
   reg __389237_389237;
   reg _389238_389238 ; 
   reg __389238_389238;
   reg _389239_389239 ; 
   reg __389239_389239;
   reg _389240_389240 ; 
   reg __389240_389240;
   reg _389241_389241 ; 
   reg __389241_389241;
   reg _389242_389242 ; 
   reg __389242_389242;
   reg _389243_389243 ; 
   reg __389243_389243;
   reg _389244_389244 ; 
   reg __389244_389244;
   reg _389245_389245 ; 
   reg __389245_389245;
   reg _389246_389246 ; 
   reg __389246_389246;
   reg _389247_389247 ; 
   reg __389247_389247;
   reg _389248_389248 ; 
   reg __389248_389248;
   reg _389249_389249 ; 
   reg __389249_389249;
   reg _389250_389250 ; 
   reg __389250_389250;
   reg _389251_389251 ; 
   reg __389251_389251;
   reg _389252_389252 ; 
   reg __389252_389252;
   reg _389253_389253 ; 
   reg __389253_389253;
   reg _389254_389254 ; 
   reg __389254_389254;
   reg _389255_389255 ; 
   reg __389255_389255;
   reg _389256_389256 ; 
   reg __389256_389256;
   reg _389257_389257 ; 
   reg __389257_389257;
   reg _389258_389258 ; 
   reg __389258_389258;
   reg _389259_389259 ; 
   reg __389259_389259;
   reg _389260_389260 ; 
   reg __389260_389260;
   reg _389261_389261 ; 
   reg __389261_389261;
   reg _389262_389262 ; 
   reg __389262_389262;
   reg _389263_389263 ; 
   reg __389263_389263;
   reg _389264_389264 ; 
   reg __389264_389264;
   reg _389265_389265 ; 
   reg __389265_389265;
   reg _389266_389266 ; 
   reg __389266_389266;
   reg _389267_389267 ; 
   reg __389267_389267;
   reg _389268_389268 ; 
   reg __389268_389268;
   reg _389269_389269 ; 
   reg __389269_389269;
   reg _389270_389270 ; 
   reg __389270_389270;
   reg _389271_389271 ; 
   reg __389271_389271;
   reg _389272_389272 ; 
   reg __389272_389272;
   reg _389273_389273 ; 
   reg __389273_389273;
   reg _389274_389274 ; 
   reg __389274_389274;
   reg _389275_389275 ; 
   reg __389275_389275;
   reg _389276_389276 ; 
   reg __389276_389276;
   reg _389277_389277 ; 
   reg __389277_389277;
   reg _389278_389278 ; 
   reg __389278_389278;
   reg _389279_389279 ; 
   reg __389279_389279;
   reg _389280_389280 ; 
   reg __389280_389280;
   reg _389281_389281 ; 
   reg __389281_389281;
   reg _389282_389282 ; 
   reg __389282_389282;
   reg _389283_389283 ; 
   reg __389283_389283;
   reg _389284_389284 ; 
   reg __389284_389284;
   reg _389285_389285 ; 
   reg __389285_389285;
   reg _389286_389286 ; 
   reg __389286_389286;
   reg _389287_389287 ; 
   reg __389287_389287;
   reg _389288_389288 ; 
   reg __389288_389288;
   reg _389289_389289 ; 
   reg __389289_389289;
   reg _389290_389290 ; 
   reg __389290_389290;
   reg _389291_389291 ; 
   reg __389291_389291;
   reg _389292_389292 ; 
   reg __389292_389292;
   reg _389293_389293 ; 
   reg __389293_389293;
   reg _389294_389294 ; 
   reg __389294_389294;
   reg _389295_389295 ; 
   reg __389295_389295;
   reg _389296_389296 ; 
   reg __389296_389296;
   reg _389297_389297 ; 
   reg __389297_389297;
   reg _389298_389298 ; 
   reg __389298_389298;
   reg _389299_389299 ; 
   reg __389299_389299;
   reg _389300_389300 ; 
   reg __389300_389300;
   reg _389301_389301 ; 
   reg __389301_389301;
   reg _389302_389302 ; 
   reg __389302_389302;
   reg _389303_389303 ; 
   reg __389303_389303;
   reg _389304_389304 ; 
   reg __389304_389304;
   reg _389305_389305 ; 
   reg __389305_389305;
   reg _389306_389306 ; 
   reg __389306_389306;
   reg _389307_389307 ; 
   reg __389307_389307;
   reg _389308_389308 ; 
   reg __389308_389308;
   reg _389309_389309 ; 
   reg __389309_389309;
   reg _389310_389310 ; 
   reg __389310_389310;
   reg _389311_389311 ; 
   reg __389311_389311;
   reg _389312_389312 ; 
   reg __389312_389312;
   reg _389313_389313 ; 
   reg __389313_389313;
   reg _389314_389314 ; 
   reg __389314_389314;
   reg _389315_389315 ; 
   reg __389315_389315;
   reg _389316_389316 ; 
   reg __389316_389316;
   reg _389317_389317 ; 
   reg __389317_389317;
   reg _389318_389318 ; 
   reg __389318_389318;
   reg _389319_389319 ; 
   reg __389319_389319;
   reg _389320_389320 ; 
   reg __389320_389320;
   reg _389321_389321 ; 
   reg __389321_389321;
   reg _389322_389322 ; 
   reg __389322_389322;
   reg _389323_389323 ; 
   reg __389323_389323;
   reg _389324_389324 ; 
   reg __389324_389324;
   reg _389325_389325 ; 
   reg __389325_389325;
   reg _389326_389326 ; 
   reg __389326_389326;
   reg _389327_389327 ; 
   reg __389327_389327;
   reg _389328_389328 ; 
   reg __389328_389328;
   reg _389329_389329 ; 
   reg __389329_389329;
   reg _389330_389330 ; 
   reg __389330_389330;
   reg _389331_389331 ; 
   reg __389331_389331;
   reg _389332_389332 ; 
   reg __389332_389332;
   reg _389333_389333 ; 
   reg __389333_389333;
   reg _389334_389334 ; 
   reg __389334_389334;
   reg _389335_389335 ; 
   reg __389335_389335;
   reg _389336_389336 ; 
   reg __389336_389336;
   reg _389337_389337 ; 
   reg __389337_389337;
   reg _389338_389338 ; 
   reg __389338_389338;
   reg _389339_389339 ; 
   reg __389339_389339;
   reg _389340_389340 ; 
   reg __389340_389340;
   reg _389341_389341 ; 
   reg __389341_389341;
   reg _389342_389342 ; 
   reg __389342_389342;
   reg _389343_389343 ; 
   reg __389343_389343;
   reg _389344_389344 ; 
   reg __389344_389344;
   reg _389345_389345 ; 
   reg __389345_389345;
   reg _389346_389346 ; 
   reg __389346_389346;
   reg _389347_389347 ; 
   reg __389347_389347;
   reg _389348_389348 ; 
   reg __389348_389348;
   reg _389349_389349 ; 
   reg __389349_389349;
   reg _389350_389350 ; 
   reg __389350_389350;
   reg _389351_389351 ; 
   reg __389351_389351;
   reg _389352_389352 ; 
   reg __389352_389352;
   reg _389353_389353 ; 
   reg __389353_389353;
   reg _389354_389354 ; 
   reg __389354_389354;
   reg _389355_389355 ; 
   reg __389355_389355;
   reg _389356_389356 ; 
   reg __389356_389356;
   reg _389357_389357 ; 
   reg __389357_389357;
   reg _389358_389358 ; 
   reg __389358_389358;
   reg _389359_389359 ; 
   reg __389359_389359;
   reg _389360_389360 ; 
   reg __389360_389360;
   reg _389361_389361 ; 
   reg __389361_389361;
   reg _389362_389362 ; 
   reg __389362_389362;
   reg _389363_389363 ; 
   reg __389363_389363;
   reg _389364_389364 ; 
   reg __389364_389364;
   reg _389365_389365 ; 
   reg __389365_389365;
   reg _389366_389366 ; 
   reg __389366_389366;
   reg _389367_389367 ; 
   reg __389367_389367;
   reg _389368_389368 ; 
   reg __389368_389368;
   reg _389369_389369 ; 
   reg __389369_389369;
   reg _389370_389370 ; 
   reg __389370_389370;
   reg _389371_389371 ; 
   reg __389371_389371;
   reg _389372_389372 ; 
   reg __389372_389372;
   reg _389373_389373 ; 
   reg __389373_389373;
   reg _389374_389374 ; 
   reg __389374_389374;
   reg _389375_389375 ; 
   reg __389375_389375;
   reg _389376_389376 ; 
   reg __389376_389376;
   reg _389377_389377 ; 
   reg __389377_389377;
   reg _389378_389378 ; 
   reg __389378_389378;
   reg _389379_389379 ; 
   reg __389379_389379;
   reg _389380_389380 ; 
   reg __389380_389380;
   reg _389381_389381 ; 
   reg __389381_389381;
   reg _389382_389382 ; 
   reg __389382_389382;
   reg _389383_389383 ; 
   reg __389383_389383;
   reg _389384_389384 ; 
   reg __389384_389384;
   reg _389385_389385 ; 
   reg __389385_389385;
   reg _389386_389386 ; 
   reg __389386_389386;
   reg _389387_389387 ; 
   reg __389387_389387;
   reg _389388_389388 ; 
   reg __389388_389388;
   reg _389389_389389 ; 
   reg __389389_389389;
   reg _389390_389390 ; 
   reg __389390_389390;
   reg _389391_389391 ; 
   reg __389391_389391;
   reg _389392_389392 ; 
   reg __389392_389392;
   reg _389393_389393 ; 
   reg __389393_389393;
   reg _389394_389394 ; 
   reg __389394_389394;
   reg _389395_389395 ; 
   reg __389395_389395;
   reg _389396_389396 ; 
   reg __389396_389396;
   reg _389397_389397 ; 
   reg __389397_389397;
   reg _389398_389398 ; 
   reg __389398_389398;
   reg _389399_389399 ; 
   reg __389399_389399;
   reg _389400_389400 ; 
   reg __389400_389400;
   reg _389401_389401 ; 
   reg __389401_389401;
   reg _389402_389402 ; 
   reg __389402_389402;
   reg _389403_389403 ; 
   reg __389403_389403;
   reg _389404_389404 ; 
   reg __389404_389404;
   reg _389405_389405 ; 
   reg __389405_389405;
   reg _389406_389406 ; 
   reg __389406_389406;
   reg _389407_389407 ; 
   reg __389407_389407;
   reg _389408_389408 ; 
   reg __389408_389408;
   reg _389409_389409 ; 
   reg __389409_389409;
   reg _389410_389410 ; 
   reg __389410_389410;
   reg _389411_389411 ; 
   reg __389411_389411;
   reg _389412_389412 ; 
   reg __389412_389412;
   reg _389413_389413 ; 
   reg __389413_389413;
   reg _389414_389414 ; 
   reg __389414_389414;
   reg _389415_389415 ; 
   reg __389415_389415;
   reg _389416_389416 ; 
   reg __389416_389416;
   reg _389417_389417 ; 
   reg __389417_389417;
   reg _389418_389418 ; 
   reg __389418_389418;
   reg _389419_389419 ; 
   reg __389419_389419;
   reg _389420_389420 ; 
   reg __389420_389420;
   reg _389421_389421 ; 
   reg __389421_389421;
   reg _389422_389422 ; 
   reg __389422_389422;
   reg _389423_389423 ; 
   reg __389423_389423;
   reg _389424_389424 ; 
   reg __389424_389424;
   reg _389425_389425 ; 
   reg __389425_389425;
   reg _389426_389426 ; 
   reg __389426_389426;
   reg _389427_389427 ; 
   reg __389427_389427;
   reg _389428_389428 ; 
   reg __389428_389428;
   reg _389429_389429 ; 
   reg __389429_389429;
   reg _389430_389430 ; 
   reg __389430_389430;
   reg _389431_389431 ; 
   reg __389431_389431;
   reg _389432_389432 ; 
   reg __389432_389432;
   reg _389433_389433 ; 
   reg __389433_389433;
   reg _389434_389434 ; 
   reg __389434_389434;
   reg _389435_389435 ; 
   reg __389435_389435;
   reg _389436_389436 ; 
   reg __389436_389436;
   reg _389437_389437 ; 
   reg __389437_389437;
   reg _389438_389438 ; 
   reg __389438_389438;
   reg _389439_389439 ; 
   reg __389439_389439;
   reg _389440_389440 ; 
   reg __389440_389440;
   reg _389441_389441 ; 
   reg __389441_389441;
   reg _389442_389442 ; 
   reg __389442_389442;
   reg _389443_389443 ; 
   reg __389443_389443;
   reg _389444_389444 ; 
   reg __389444_389444;
   reg _389445_389445 ; 
   reg __389445_389445;
   reg _389446_389446 ; 
   reg __389446_389446;
   reg _389447_389447 ; 
   reg __389447_389447;
   reg _389448_389448 ; 
   reg __389448_389448;
   reg _389449_389449 ; 
   reg __389449_389449;
   reg _389450_389450 ; 
   reg __389450_389450;
   reg _389451_389451 ; 
   reg __389451_389451;
   reg _389452_389452 ; 
   reg __389452_389452;
   reg _389453_389453 ; 
   reg __389453_389453;
   reg _389454_389454 ; 
   reg __389454_389454;
   reg _389455_389455 ; 
   reg __389455_389455;
   reg _389456_389456 ; 
   reg __389456_389456;
   reg _389457_389457 ; 
   reg __389457_389457;
   reg _389458_389458 ; 
   reg __389458_389458;
   reg _389459_389459 ; 
   reg __389459_389459;
   reg _389460_389460 ; 
   reg __389460_389460;
   reg _389461_389461 ; 
   reg __389461_389461;
   reg _389462_389462 ; 
   reg __389462_389462;
   reg _389463_389463 ; 
   reg __389463_389463;
   reg _389464_389464 ; 
   reg __389464_389464;
   reg _389465_389465 ; 
   reg __389465_389465;
   reg _389466_389466 ; 
   reg __389466_389466;
   reg _389467_389467 ; 
   reg __389467_389467;
   reg _389468_389468 ; 
   reg __389468_389468;
   reg _389469_389469 ; 
   reg __389469_389469;
   reg _389470_389470 ; 
   reg __389470_389470;
   reg _389471_389471 ; 
   reg __389471_389471;
   reg _389472_389472 ; 
   reg __389472_389472;
   reg _389473_389473 ; 
   reg __389473_389473;
   reg _389474_389474 ; 
   reg __389474_389474;
   reg _389475_389475 ; 
   reg __389475_389475;
   reg _389476_389476 ; 
   reg __389476_389476;
   reg _389477_389477 ; 
   reg __389477_389477;
   reg _389478_389478 ; 
   reg __389478_389478;
   reg _389479_389479 ; 
   reg __389479_389479;
   reg _389480_389480 ; 
   reg __389480_389480;
   reg _389481_389481 ; 
   reg __389481_389481;
   reg _389482_389482 ; 
   reg __389482_389482;
   reg _389483_389483 ; 
   reg __389483_389483;
   reg _389484_389484 ; 
   reg __389484_389484;
   reg _389485_389485 ; 
   reg __389485_389485;
   reg _389486_389486 ; 
   reg __389486_389486;
   reg _389487_389487 ; 
   reg __389487_389487;
   reg _389488_389488 ; 
   reg __389488_389488;
   reg _389489_389489 ; 
   reg __389489_389489;
   reg _389490_389490 ; 
   reg __389490_389490;
   reg _389491_389491 ; 
   reg __389491_389491;
   reg _389492_389492 ; 
   reg __389492_389492;
   reg _389493_389493 ; 
   reg __389493_389493;
   reg _389494_389494 ; 
   reg __389494_389494;
   reg _389495_389495 ; 
   reg __389495_389495;
   reg _389496_389496 ; 
   reg __389496_389496;
   reg _389497_389497 ; 
   reg __389497_389497;
   reg _389498_389498 ; 
   reg __389498_389498;
   reg _389499_389499 ; 
   reg __389499_389499;
   reg _389500_389500 ; 
   reg __389500_389500;
   reg _389501_389501 ; 
   reg __389501_389501;
   reg _389502_389502 ; 
   reg __389502_389502;
   reg _389503_389503 ; 
   reg __389503_389503;
   reg _389504_389504 ; 
   reg __389504_389504;
   reg _389505_389505 ; 
   reg __389505_389505;
   reg _389506_389506 ; 
   reg __389506_389506;
   reg _389507_389507 ; 
   reg __389507_389507;
   reg _389508_389508 ; 
   reg __389508_389508;
   reg _389509_389509 ; 
   reg __389509_389509;
   reg _389510_389510 ; 
   reg __389510_389510;
   reg _389511_389511 ; 
   reg __389511_389511;
   reg _389512_389512 ; 
   reg __389512_389512;
   reg _389513_389513 ; 
   reg __389513_389513;
   reg _389514_389514 ; 
   reg __389514_389514;
   reg _389515_389515 ; 
   reg __389515_389515;
   reg _389516_389516 ; 
   reg __389516_389516;
   reg _389517_389517 ; 
   reg __389517_389517;
   reg _389518_389518 ; 
   reg __389518_389518;
   reg _389519_389519 ; 
   reg __389519_389519;
   reg _389520_389520 ; 
   reg __389520_389520;
   reg _389521_389521 ; 
   reg __389521_389521;
   reg _389522_389522 ; 
   reg __389522_389522;
   reg _389523_389523 ; 
   reg __389523_389523;
   reg _389524_389524 ; 
   reg __389524_389524;
   reg _389525_389525 ; 
   reg __389525_389525;
   reg _389526_389526 ; 
   reg __389526_389526;
   reg _389527_389527 ; 
   reg __389527_389527;
   reg _389528_389528 ; 
   reg __389528_389528;
   reg _389529_389529 ; 
   reg __389529_389529;
   reg _389530_389530 ; 
   reg __389530_389530;
   reg _389531_389531 ; 
   reg __389531_389531;
   reg _389532_389532 ; 
   reg __389532_389532;
   reg _389533_389533 ; 
   reg __389533_389533;
   reg _389534_389534 ; 
   reg __389534_389534;
   reg _389535_389535 ; 
   reg __389535_389535;
   reg _389536_389536 ; 
   reg __389536_389536;
   reg _389537_389537 ; 
   reg __389537_389537;
   reg _389538_389538 ; 
   reg __389538_389538;
   reg _389539_389539 ; 
   reg __389539_389539;
   reg _389540_389540 ; 
   reg __389540_389540;
   reg _389541_389541 ; 
   reg __389541_389541;
   reg _389542_389542 ; 
   reg __389542_389542;
   reg _389543_389543 ; 
   reg __389543_389543;
   reg _389544_389544 ; 
   reg __389544_389544;
   reg _389545_389545 ; 
   reg __389545_389545;
   reg _389546_389546 ; 
   reg __389546_389546;
   reg _389547_389547 ; 
   reg __389547_389547;
   reg _389548_389548 ; 
   reg __389548_389548;
   reg _389549_389549 ; 
   reg __389549_389549;
   reg _389550_389550 ; 
   reg __389550_389550;
   reg _389551_389551 ; 
   reg __389551_389551;
   reg _389552_389552 ; 
   reg __389552_389552;
   reg _389553_389553 ; 
   reg __389553_389553;
   reg _389554_389554 ; 
   reg __389554_389554;
   reg _389555_389555 ; 
   reg __389555_389555;
   reg _389556_389556 ; 
   reg __389556_389556;
   reg _389557_389557 ; 
   reg __389557_389557;
   reg _389558_389558 ; 
   reg __389558_389558;
   reg _389559_389559 ; 
   reg __389559_389559;
   reg _389560_389560 ; 
   reg __389560_389560;
   reg _389561_389561 ; 
   reg __389561_389561;
   reg _389562_389562 ; 
   reg __389562_389562;
   reg _389563_389563 ; 
   reg __389563_389563;
   reg _389564_389564 ; 
   reg __389564_389564;
   reg _389565_389565 ; 
   reg __389565_389565;
   reg _389566_389566 ; 
   reg __389566_389566;
   reg _389567_389567 ; 
   reg __389567_389567;
   reg _389568_389568 ; 
   reg __389568_389568;
   reg _389569_389569 ; 
   reg __389569_389569;
   reg _389570_389570 ; 
   reg __389570_389570;
   reg _389571_389571 ; 
   reg __389571_389571;
   reg _389572_389572 ; 
   reg __389572_389572;
   reg _389573_389573 ; 
   reg __389573_389573;
   reg _389574_389574 ; 
   reg __389574_389574;
   reg _389575_389575 ; 
   reg __389575_389575;
   reg _389576_389576 ; 
   reg __389576_389576;
   reg _389577_389577 ; 
   reg __389577_389577;
   reg _389578_389578 ; 
   reg __389578_389578;
   reg _389579_389579 ; 
   reg __389579_389579;
   reg _389580_389580 ; 
   reg __389580_389580;
   reg _389581_389581 ; 
   reg __389581_389581;
   reg _389582_389582 ; 
   reg __389582_389582;
   reg _389583_389583 ; 
   reg __389583_389583;
   reg _389584_389584 ; 
   reg __389584_389584;
   reg _389585_389585 ; 
   reg __389585_389585;
   reg _389586_389586 ; 
   reg __389586_389586;
   reg _389587_389587 ; 
   reg __389587_389587;
   reg _389588_389588 ; 
   reg __389588_389588;
   reg _389589_389589 ; 
   reg __389589_389589;
   reg _389590_389590 ; 
   reg __389590_389590;
   reg _389591_389591 ; 
   reg __389591_389591;
   reg _389592_389592 ; 
   reg __389592_389592;
   reg _389593_389593 ; 
   reg __389593_389593;
   reg _389594_389594 ; 
   reg __389594_389594;
   reg _389595_389595 ; 
   reg __389595_389595;
   reg _389596_389596 ; 
   reg __389596_389596;
   reg _389597_389597 ; 
   reg __389597_389597;
   reg _389598_389598 ; 
   reg __389598_389598;
   reg _389599_389599 ; 
   reg __389599_389599;
   reg _389600_389600 ; 
   reg __389600_389600;
   reg _389601_389601 ; 
   reg __389601_389601;
   reg _389602_389602 ; 
   reg __389602_389602;
   reg _389603_389603 ; 
   reg __389603_389603;
   reg _389604_389604 ; 
   reg __389604_389604;
   reg _389605_389605 ; 
   reg __389605_389605;
   reg _389606_389606 ; 
   reg __389606_389606;
   reg _389607_389607 ; 
   reg __389607_389607;
   reg _389608_389608 ; 
   reg __389608_389608;
   reg _389609_389609 ; 
   reg __389609_389609;
   reg _389610_389610 ; 
   reg __389610_389610;
   reg _389611_389611 ; 
   reg __389611_389611;
   reg _389612_389612 ; 
   reg __389612_389612;
   reg _389613_389613 ; 
   reg __389613_389613;
   reg _389614_389614 ; 
   reg __389614_389614;
   reg _389615_389615 ; 
   reg __389615_389615;
   reg _389616_389616 ; 
   reg __389616_389616;
   reg _389617_389617 ; 
   reg __389617_389617;
   reg _389618_389618 ; 
   reg __389618_389618;
   reg _389619_389619 ; 
   reg __389619_389619;
   reg _389620_389620 ; 
   reg __389620_389620;
   reg _389621_389621 ; 
   reg __389621_389621;
   reg _389622_389622 ; 
   reg __389622_389622;
   reg _389623_389623 ; 
   reg __389623_389623;
   reg _389624_389624 ; 
   reg __389624_389624;
   reg _389625_389625 ; 
   reg __389625_389625;
   reg _389626_389626 ; 
   reg __389626_389626;
   reg _389627_389627 ; 
   reg __389627_389627;
   reg _389628_389628 ; 
   reg __389628_389628;
   reg _389629_389629 ; 
   reg __389629_389629;
   reg _389630_389630 ; 
   reg __389630_389630;
   reg _389631_389631 ; 
   reg __389631_389631;
   reg _389632_389632 ; 
   reg __389632_389632;
   reg _389633_389633 ; 
   reg __389633_389633;
   reg _389634_389634 ; 
   reg __389634_389634;
   reg _389635_389635 ; 
   reg __389635_389635;
   reg _389636_389636 ; 
   reg __389636_389636;
   reg _389637_389637 ; 
   reg __389637_389637;
   reg _389638_389638 ; 
   reg __389638_389638;
   reg _389639_389639 ; 
   reg __389639_389639;
   reg _389640_389640 ; 
   reg __389640_389640;
   reg _389641_389641 ; 
   reg __389641_389641;
   reg _389642_389642 ; 
   reg __389642_389642;
   reg _389643_389643 ; 
   reg __389643_389643;
   reg _389644_389644 ; 
   reg __389644_389644;
   reg _389645_389645 ; 
   reg __389645_389645;
   reg _389646_389646 ; 
   reg __389646_389646;
   reg _389647_389647 ; 
   reg __389647_389647;
   reg _389648_389648 ; 
   reg __389648_389648;
   reg _389649_389649 ; 
   reg __389649_389649;
   reg _389650_389650 ; 
   reg __389650_389650;
   reg _389651_389651 ; 
   reg __389651_389651;
   reg _389652_389652 ; 
   reg __389652_389652;
   reg _389653_389653 ; 
   reg __389653_389653;
   reg _389654_389654 ; 
   reg __389654_389654;
   reg _389655_389655 ; 
   reg __389655_389655;
   reg _389656_389656 ; 
   reg __389656_389656;
   reg _389657_389657 ; 
   reg __389657_389657;
   reg _389658_389658 ; 
   reg __389658_389658;
   reg _389659_389659 ; 
   reg __389659_389659;
   reg _389660_389660 ; 
   reg __389660_389660;
   reg _389661_389661 ; 
   reg __389661_389661;
   reg _389662_389662 ; 
   reg __389662_389662;
   reg _389663_389663 ; 
   reg __389663_389663;
   reg _389664_389664 ; 
   reg __389664_389664;
   reg _389665_389665 ; 
   reg __389665_389665;
   reg _389666_389666 ; 
   reg __389666_389666;
   reg _389667_389667 ; 
   reg __389667_389667;
   reg _389668_389668 ; 
   reg __389668_389668;
   reg _389669_389669 ; 
   reg __389669_389669;
   reg _389670_389670 ; 
   reg __389670_389670;
   reg _389671_389671 ; 
   reg __389671_389671;
   reg _389672_389672 ; 
   reg __389672_389672;
   reg _389673_389673 ; 
   reg __389673_389673;
   reg _389674_389674 ; 
   reg __389674_389674;
   reg _389675_389675 ; 
   reg __389675_389675;
   reg _389676_389676 ; 
   reg __389676_389676;
   reg _389677_389677 ; 
   reg __389677_389677;
   reg _389678_389678 ; 
   reg __389678_389678;
   reg _389679_389679 ; 
   reg __389679_389679;
   reg _389680_389680 ; 
   reg __389680_389680;
   reg _389681_389681 ; 
   reg __389681_389681;
   reg _389682_389682 ; 
   reg __389682_389682;
   reg _389683_389683 ; 
   reg __389683_389683;
   reg _389684_389684 ; 
   reg __389684_389684;
   reg _389685_389685 ; 
   reg __389685_389685;
   reg _389686_389686 ; 
   reg __389686_389686;
   reg _389687_389687 ; 
   reg __389687_389687;
   reg _389688_389688 ; 
   reg __389688_389688;
   reg _389689_389689 ; 
   reg __389689_389689;
   reg _389690_389690 ; 
   reg __389690_389690;
   reg _389691_389691 ; 
   reg __389691_389691;
   reg _389692_389692 ; 
   reg __389692_389692;
   reg _389693_389693 ; 
   reg __389693_389693;
   reg _389694_389694 ; 
   reg __389694_389694;
   reg _389695_389695 ; 
   reg __389695_389695;
   reg _389696_389696 ; 
   reg __389696_389696;
   reg _389697_389697 ; 
   reg __389697_389697;
   reg _389698_389698 ; 
   reg __389698_389698;
   reg _389699_389699 ; 
   reg __389699_389699;
   reg _389700_389700 ; 
   reg __389700_389700;
   reg _389701_389701 ; 
   reg __389701_389701;
   reg _389702_389702 ; 
   reg __389702_389702;
   reg _389703_389703 ; 
   reg __389703_389703;
   reg _389704_389704 ; 
   reg __389704_389704;
   reg _389705_389705 ; 
   reg __389705_389705;
   reg _389706_389706 ; 
   reg __389706_389706;
   reg _389707_389707 ; 
   reg __389707_389707;
   reg _389708_389708 ; 
   reg __389708_389708;
   reg _389709_389709 ; 
   reg __389709_389709;
   reg _389710_389710 ; 
   reg __389710_389710;
   reg _389711_389711 ; 
   reg __389711_389711;
   reg _389712_389712 ; 
   reg __389712_389712;
   reg _389713_389713 ; 
   reg __389713_389713;
   reg _389714_389714 ; 
   reg __389714_389714;
   reg _389715_389715 ; 
   reg __389715_389715;
   reg _389716_389716 ; 
   reg __389716_389716;
   reg _389717_389717 ; 
   reg __389717_389717;
   reg _389718_389718 ; 
   reg __389718_389718;
   reg _389719_389719 ; 
   reg __389719_389719;
   reg _389720_389720 ; 
   reg __389720_389720;
   reg _389721_389721 ; 
   reg __389721_389721;
   reg _389722_389722 ; 
   reg __389722_389722;
   reg _389723_389723 ; 
   reg __389723_389723;
   reg _389724_389724 ; 
   reg __389724_389724;
   reg _389725_389725 ; 
   reg __389725_389725;
   reg _389726_389726 ; 
   reg __389726_389726;
   reg _389727_389727 ; 
   reg __389727_389727;
   reg _389728_389728 ; 
   reg __389728_389728;
   reg _389729_389729 ; 
   reg __389729_389729;
   reg _389730_389730 ; 
   reg __389730_389730;
   reg _389731_389731 ; 
   reg __389731_389731;
   reg _389732_389732 ; 
   reg __389732_389732;
   reg _389733_389733 ; 
   reg __389733_389733;
   reg _389734_389734 ; 
   reg __389734_389734;
   reg _389735_389735 ; 
   reg __389735_389735;
   reg _389736_389736 ; 
   reg __389736_389736;
   reg _389737_389737 ; 
   reg __389737_389737;
   reg _389738_389738 ; 
   reg __389738_389738;
   reg _389739_389739 ; 
   reg __389739_389739;
   reg _389740_389740 ; 
   reg __389740_389740;
   reg _389741_389741 ; 
   reg __389741_389741;
   reg _389742_389742 ; 
   reg __389742_389742;
   reg _389743_389743 ; 
   reg __389743_389743;
   reg _389744_389744 ; 
   reg __389744_389744;
   reg _389745_389745 ; 
   reg __389745_389745;
   reg _389746_389746 ; 
   reg __389746_389746;
   reg _389747_389747 ; 
   reg __389747_389747;
   reg _389748_389748 ; 
   reg __389748_389748;
   reg _389749_389749 ; 
   reg __389749_389749;
   reg _389750_389750 ; 
   reg __389750_389750;
   reg _389751_389751 ; 
   reg __389751_389751;
   reg _389752_389752 ; 
   reg __389752_389752;
   reg _389753_389753 ; 
   reg __389753_389753;
   reg _389754_389754 ; 
   reg __389754_389754;
   reg _389755_389755 ; 
   reg __389755_389755;
   reg _389756_389756 ; 
   reg __389756_389756;
   reg _389757_389757 ; 
   reg __389757_389757;
   reg _389758_389758 ; 
   reg __389758_389758;
   reg _389759_389759 ; 
   reg __389759_389759;
   reg _389760_389760 ; 
   reg __389760_389760;
   reg _389761_389761 ; 
   reg __389761_389761;
   reg _389762_389762 ; 
   reg __389762_389762;
   reg _389763_389763 ; 
   reg __389763_389763;
   reg _389764_389764 ; 
   reg __389764_389764;
   reg _389765_389765 ; 
   reg __389765_389765;
   reg _389766_389766 ; 
   reg __389766_389766;
   reg _389767_389767 ; 
   reg __389767_389767;
   reg _389768_389768 ; 
   reg __389768_389768;
   reg _389769_389769 ; 
   reg __389769_389769;
   reg _389770_389770 ; 
   reg __389770_389770;
   reg _389771_389771 ; 
   reg __389771_389771;
   reg _389772_389772 ; 
   reg __389772_389772;
   reg _389773_389773 ; 
   reg __389773_389773;
   reg _389774_389774 ; 
   reg __389774_389774;
   reg _389775_389775 ; 
   reg __389775_389775;
   reg _389776_389776 ; 
   reg __389776_389776;
   reg _389777_389777 ; 
   reg __389777_389777;
   reg _389778_389778 ; 
   reg __389778_389778;
   reg _389779_389779 ; 
   reg __389779_389779;
   reg _389780_389780 ; 
   reg __389780_389780;
   reg _389781_389781 ; 
   reg __389781_389781;
   reg _389782_389782 ; 
   reg __389782_389782;
   reg _389783_389783 ; 
   reg __389783_389783;
   reg _389784_389784 ; 
   reg __389784_389784;
   reg _389785_389785 ; 
   reg __389785_389785;
   reg _389786_389786 ; 
   reg __389786_389786;
   reg _389787_389787 ; 
   reg __389787_389787;
   reg _389788_389788 ; 
   reg __389788_389788;
   reg _389789_389789 ; 
   reg __389789_389789;
   reg _389790_389790 ; 
   reg __389790_389790;
   reg _389791_389791 ; 
   reg __389791_389791;
   reg _389792_389792 ; 
   reg __389792_389792;
   reg _389793_389793 ; 
   reg __389793_389793;
   reg _389794_389794 ; 
   reg __389794_389794;
   reg _389795_389795 ; 
   reg __389795_389795;
   reg _389796_389796 ; 
   reg __389796_389796;
   reg _389797_389797 ; 
   reg __389797_389797;
   reg _389798_389798 ; 
   reg __389798_389798;
   reg _389799_389799 ; 
   reg __389799_389799;
   reg _389800_389800 ; 
   reg __389800_389800;
   reg _389801_389801 ; 
   reg __389801_389801;
   reg _389802_389802 ; 
   reg __389802_389802;
   reg _389803_389803 ; 
   reg __389803_389803;
   reg _389804_389804 ; 
   reg __389804_389804;
   reg _389805_389805 ; 
   reg __389805_389805;
   reg _389806_389806 ; 
   reg __389806_389806;
   reg _389807_389807 ; 
   reg __389807_389807;
   reg _389808_389808 ; 
   reg __389808_389808;
   reg _389809_389809 ; 
   reg __389809_389809;
   reg _389810_389810 ; 
   reg __389810_389810;
   reg _389811_389811 ; 
   reg __389811_389811;
   reg _389812_389812 ; 
   reg __389812_389812;
   reg _389813_389813 ; 
   reg __389813_389813;
   reg _389814_389814 ; 
   reg __389814_389814;
   reg _389815_389815 ; 
   reg __389815_389815;
   reg _389816_389816 ; 
   reg __389816_389816;
   reg _389817_389817 ; 
   reg __389817_389817;
   reg _389818_389818 ; 
   reg __389818_389818;
   reg _389819_389819 ; 
   reg __389819_389819;
   reg _389820_389820 ; 
   reg __389820_389820;
   reg _389821_389821 ; 
   reg __389821_389821;
   reg _389822_389822 ; 
   reg __389822_389822;
   reg _389823_389823 ; 
   reg __389823_389823;
   reg _389824_389824 ; 
   reg __389824_389824;
   reg _389825_389825 ; 
   reg __389825_389825;
   reg _389826_389826 ; 
   reg __389826_389826;
   reg _389827_389827 ; 
   reg __389827_389827;
   reg _389828_389828 ; 
   reg __389828_389828;
   reg _389829_389829 ; 
   reg __389829_389829;
   reg _389830_389830 ; 
   reg __389830_389830;
   reg _389831_389831 ; 
   reg __389831_389831;
   reg _389832_389832 ; 
   reg __389832_389832;
   reg _389833_389833 ; 
   reg __389833_389833;
   reg _389834_389834 ; 
   reg __389834_389834;
   reg _389835_389835 ; 
   reg __389835_389835;
   reg _389836_389836 ; 
   reg __389836_389836;
   reg _389837_389837 ; 
   reg __389837_389837;
   reg _389838_389838 ; 
   reg __389838_389838;
   reg _389839_389839 ; 
   reg __389839_389839;
   reg _389840_389840 ; 
   reg __389840_389840;
   reg _389841_389841 ; 
   reg __389841_389841;
   reg _389842_389842 ; 
   reg __389842_389842;
   reg _389843_389843 ; 
   reg __389843_389843;
   reg _389844_389844 ; 
   reg __389844_389844;
   reg _389845_389845 ; 
   reg __389845_389845;
   reg _389846_389846 ; 
   reg __389846_389846;
   reg _389847_389847 ; 
   reg __389847_389847;
   reg _389848_389848 ; 
   reg __389848_389848;
   reg _389849_389849 ; 
   reg __389849_389849;
   reg _389850_389850 ; 
   reg __389850_389850;
   reg _389851_389851 ; 
   reg __389851_389851;
   reg _389852_389852 ; 
   reg __389852_389852;
   reg _389853_389853 ; 
   reg __389853_389853;
   reg _389854_389854 ; 
   reg __389854_389854;
   reg _389855_389855 ; 
   reg __389855_389855;
   reg _389856_389856 ; 
   reg __389856_389856;
   reg _389857_389857 ; 
   reg __389857_389857;
   reg _389858_389858 ; 
   reg __389858_389858;
   reg _389859_389859 ; 
   reg __389859_389859;
   reg _389860_389860 ; 
   reg __389860_389860;
   reg _389861_389861 ; 
   reg __389861_389861;
   reg _389862_389862 ; 
   reg __389862_389862;
   reg _389863_389863 ; 
   reg __389863_389863;
   reg _389864_389864 ; 
   reg __389864_389864;
   reg _389865_389865 ; 
   reg __389865_389865;
   reg _389866_389866 ; 
   reg __389866_389866;
   reg _389867_389867 ; 
   reg __389867_389867;
   reg _389868_389868 ; 
   reg __389868_389868;
   reg _389869_389869 ; 
   reg __389869_389869;
   reg _389870_389870 ; 
   reg __389870_389870;
   reg _389871_389871 ; 
   reg __389871_389871;
   reg _389872_389872 ; 
   reg __389872_389872;
   reg _389873_389873 ; 
   reg __389873_389873;
   reg _389874_389874 ; 
   reg __389874_389874;
   reg _389875_389875 ; 
   reg __389875_389875;
   reg _389876_389876 ; 
   reg __389876_389876;
   reg _389877_389877 ; 
   reg __389877_389877;
   reg _389878_389878 ; 
   reg __389878_389878;
   reg _389879_389879 ; 
   reg __389879_389879;
   reg _389880_389880 ; 
   reg __389880_389880;
   reg _389881_389881 ; 
   reg __389881_389881;
   reg _389882_389882 ; 
   reg __389882_389882;
   reg _389883_389883 ; 
   reg __389883_389883;
   reg _389884_389884 ; 
   reg __389884_389884;
   reg _389885_389885 ; 
   reg __389885_389885;
   reg _389886_389886 ; 
   reg __389886_389886;
   reg _389887_389887 ; 
   reg __389887_389887;
   reg _389888_389888 ; 
   reg __389888_389888;
   reg _389889_389889 ; 
   reg __389889_389889;
   reg _389890_389890 ; 
   reg __389890_389890;
   reg _389891_389891 ; 
   reg __389891_389891;
   reg _389892_389892 ; 
   reg __389892_389892;
   reg _389893_389893 ; 
   reg __389893_389893;
   reg _389894_389894 ; 
   reg __389894_389894;
   reg _389895_389895 ; 
   reg __389895_389895;
   reg _389896_389896 ; 
   reg __389896_389896;
   reg _389897_389897 ; 
   reg __389897_389897;
   reg _389898_389898 ; 
   reg __389898_389898;
   reg _389899_389899 ; 
   reg __389899_389899;
   reg _389900_389900 ; 
   reg __389900_389900;
   reg _389901_389901 ; 
   reg __389901_389901;
   reg _389902_389902 ; 
   reg __389902_389902;
   reg _389903_389903 ; 
   reg __389903_389903;
   reg _389904_389904 ; 
   reg __389904_389904;
   reg _389905_389905 ; 
   reg __389905_389905;
   reg _389906_389906 ; 
   reg __389906_389906;
   reg _389907_389907 ; 
   reg __389907_389907;
   reg _389908_389908 ; 
   reg __389908_389908;
   reg _389909_389909 ; 
   reg __389909_389909;
   reg _389910_389910 ; 
   reg __389910_389910;
   reg _389911_389911 ; 
   reg __389911_389911;
   reg _389912_389912 ; 
   reg __389912_389912;
   reg _389913_389913 ; 
   reg __389913_389913;
   reg _389914_389914 ; 
   reg __389914_389914;
   reg _389915_389915 ; 
   reg __389915_389915;
   reg _389916_389916 ; 
   reg __389916_389916;
   reg _389917_389917 ; 
   reg __389917_389917;
   reg _389918_389918 ; 
   reg __389918_389918;
   reg _389919_389919 ; 
   reg __389919_389919;
   reg _389920_389920 ; 
   reg __389920_389920;
   reg _389921_389921 ; 
   reg __389921_389921;
   reg _389922_389922 ; 
   reg __389922_389922;
   reg _389923_389923 ; 
   reg __389923_389923;
   reg _389924_389924 ; 
   reg __389924_389924;
   reg _389925_389925 ; 
   reg __389925_389925;
   reg _389926_389926 ; 
   reg __389926_389926;
   reg _389927_389927 ; 
   reg __389927_389927;
   reg _389928_389928 ; 
   reg __389928_389928;
   reg _389929_389929 ; 
   reg __389929_389929;
   reg _389930_389930 ; 
   reg __389930_389930;
   reg _389931_389931 ; 
   reg __389931_389931;
   reg _389932_389932 ; 
   reg __389932_389932;
   reg _389933_389933 ; 
   reg __389933_389933;
   reg _389934_389934 ; 
   reg __389934_389934;
   reg _389935_389935 ; 
   reg __389935_389935;
   reg _389936_389936 ; 
   reg __389936_389936;
   reg _389937_389937 ; 
   reg __389937_389937;
   reg _389938_389938 ; 
   reg __389938_389938;
   reg _389939_389939 ; 
   reg __389939_389939;
   reg _389940_389940 ; 
   reg __389940_389940;
   reg _389941_389941 ; 
   reg __389941_389941;
   reg _389942_389942 ; 
   reg __389942_389942;
   reg _389943_389943 ; 
   reg __389943_389943;
   reg _389944_389944 ; 
   reg __389944_389944;
   reg _389945_389945 ; 
   reg __389945_389945;
   reg _389946_389946 ; 
   reg __389946_389946;
   reg _389947_389947 ; 
   reg __389947_389947;
   reg _389948_389948 ; 
   reg __389948_389948;
   reg _389949_389949 ; 
   reg __389949_389949;
   reg _389950_389950 ; 
   reg __389950_389950;
   reg _389951_389951 ; 
   reg __389951_389951;
   reg _389952_389952 ; 
   reg __389952_389952;
   reg _389953_389953 ; 
   reg __389953_389953;
   reg _389954_389954 ; 
   reg __389954_389954;
   reg _389955_389955 ; 
   reg __389955_389955;
   reg _389956_389956 ; 
   reg __389956_389956;
   reg _389957_389957 ; 
   reg __389957_389957;
   reg _389958_389958 ; 
   reg __389958_389958;
   reg _389959_389959 ; 
   reg __389959_389959;
   reg _389960_389960 ; 
   reg __389960_389960;
   reg _389961_389961 ; 
   reg __389961_389961;
   reg _389962_389962 ; 
   reg __389962_389962;
   reg _389963_389963 ; 
   reg __389963_389963;
   reg _389964_389964 ; 
   reg __389964_389964;
   reg _389965_389965 ; 
   reg __389965_389965;
   reg _389966_389966 ; 
   reg __389966_389966;
   reg _389967_389967 ; 
   reg __389967_389967;
   reg _389968_389968 ; 
   reg __389968_389968;
   reg _389969_389969 ; 
   reg __389969_389969;
   reg _389970_389970 ; 
   reg __389970_389970;
   reg _389971_389971 ; 
   reg __389971_389971;
   reg _389972_389972 ; 
   reg __389972_389972;
   reg _389973_389973 ; 
   reg __389973_389973;
   reg _389974_389974 ; 
   reg __389974_389974;
   reg _389975_389975 ; 
   reg __389975_389975;
   reg _389976_389976 ; 
   reg __389976_389976;
   reg _389977_389977 ; 
   reg __389977_389977;
   reg _389978_389978 ; 
   reg __389978_389978;
   reg _389979_389979 ; 
   reg __389979_389979;
   reg _389980_389980 ; 
   reg __389980_389980;
   reg _389981_389981 ; 
   reg __389981_389981;
   reg _389982_389982 ; 
   reg __389982_389982;
   reg _389983_389983 ; 
   reg __389983_389983;
   reg _389984_389984 ; 
   reg __389984_389984;
   reg _389985_389985 ; 
   reg __389985_389985;
   reg _389986_389986 ; 
   reg __389986_389986;
   reg _389987_389987 ; 
   reg __389987_389987;
   reg _389988_389988 ; 
   reg __389988_389988;
   reg _389989_389989 ; 
   reg __389989_389989;
   reg _389990_389990 ; 
   reg __389990_389990;
   reg _389991_389991 ; 
   reg __389991_389991;
   reg _389992_389992 ; 
   reg __389992_389992;
   reg _389993_389993 ; 
   reg __389993_389993;
   reg _389994_389994 ; 
   reg __389994_389994;
   reg _389995_389995 ; 
   reg __389995_389995;
   reg _389996_389996 ; 
   reg __389996_389996;
   reg _389997_389997 ; 
   reg __389997_389997;
   reg _389998_389998 ; 
   reg __389998_389998;
   reg _389999_389999 ; 
   reg __389999_389999;
   reg _390000_390000 ; 
   reg __390000_390000;
   reg _390001_390001 ; 
   reg __390001_390001;
   reg _390002_390002 ; 
   reg __390002_390002;
   reg _390003_390003 ; 
   reg __390003_390003;
   reg _390004_390004 ; 
   reg __390004_390004;
   reg _390005_390005 ; 
   reg __390005_390005;
   reg _390006_390006 ; 
   reg __390006_390006;
   reg _390007_390007 ; 
   reg __390007_390007;
   reg _390008_390008 ; 
   reg __390008_390008;
   reg _390009_390009 ; 
   reg __390009_390009;
   reg _390010_390010 ; 
   reg __390010_390010;
   reg _390011_390011 ; 
   reg __390011_390011;
   reg _390012_390012 ; 
   reg __390012_390012;
   reg _390013_390013 ; 
   reg __390013_390013;
   reg _390014_390014 ; 
   reg __390014_390014;
   reg _390015_390015 ; 
   reg __390015_390015;
   reg _390016_390016 ; 
   reg __390016_390016;
   reg _390017_390017 ; 
   reg __390017_390017;
   reg _390018_390018 ; 
   reg __390018_390018;
   reg _390019_390019 ; 
   reg __390019_390019;
   reg _390020_390020 ; 
   reg __390020_390020;
   reg _390021_390021 ; 
   reg __390021_390021;
   reg _390022_390022 ; 
   reg __390022_390022;
   reg _390023_390023 ; 
   reg __390023_390023;
   reg _390024_390024 ; 
   reg __390024_390024;
   reg _390025_390025 ; 
   reg __390025_390025;
   reg _390026_390026 ; 
   reg __390026_390026;
   reg _390027_390027 ; 
   reg __390027_390027;
   reg _390028_390028 ; 
   reg __390028_390028;
   reg _390029_390029 ; 
   reg __390029_390029;
   reg _390030_390030 ; 
   reg __390030_390030;
   reg _390031_390031 ; 
   reg __390031_390031;
   reg _390032_390032 ; 
   reg __390032_390032;
   reg _390033_390033 ; 
   reg __390033_390033;
   reg _390034_390034 ; 
   reg __390034_390034;
   reg _390035_390035 ; 
   reg __390035_390035;
   reg _390036_390036 ; 
   reg __390036_390036;
   reg _390037_390037 ; 
   reg __390037_390037;
   reg _390038_390038 ; 
   reg __390038_390038;
   reg _390039_390039 ; 
   reg __390039_390039;
   reg _390040_390040 ; 
   reg __390040_390040;
   reg _390041_390041 ; 
   reg __390041_390041;
   reg _390042_390042 ; 
   reg __390042_390042;
   reg _390043_390043 ; 
   reg __390043_390043;
   reg _390044_390044 ; 
   reg __390044_390044;
   reg _390045_390045 ; 
   reg __390045_390045;
   reg _390046_390046 ; 
   reg __390046_390046;
   reg _390047_390047 ; 
   reg __390047_390047;
   reg _390048_390048 ; 
   reg __390048_390048;
   reg _390049_390049 ; 
   reg __390049_390049;
   reg _390050_390050 ; 
   reg __390050_390050;
   reg _390051_390051 ; 
   reg __390051_390051;
   reg _390052_390052 ; 
   reg __390052_390052;
   reg _390053_390053 ; 
   reg __390053_390053;
   reg _390054_390054 ; 
   reg __390054_390054;
   reg _390055_390055 ; 
   reg __390055_390055;
   reg _390056_390056 ; 
   reg __390056_390056;
   reg _390057_390057 ; 
   reg __390057_390057;
   reg _390058_390058 ; 
   reg __390058_390058;
   reg _390059_390059 ; 
   reg __390059_390059;
   reg _390060_390060 ; 
   reg __390060_390060;
   reg _390061_390061 ; 
   reg __390061_390061;
   reg _390062_390062 ; 
   reg __390062_390062;
   reg _390063_390063 ; 
   reg __390063_390063;
   reg _390064_390064 ; 
   reg __390064_390064;
   reg _390065_390065 ; 
   reg __390065_390065;
   reg _390066_390066 ; 
   reg __390066_390066;
   reg _390067_390067 ; 
   reg __390067_390067;
   reg _390068_390068 ; 
   reg __390068_390068;
   reg _390069_390069 ; 
   reg __390069_390069;
   reg _390070_390070 ; 
   reg __390070_390070;
   reg _390071_390071 ; 
   reg __390071_390071;
   reg _390072_390072 ; 
   reg __390072_390072;
   reg _390073_390073 ; 
   reg __390073_390073;
   reg _390074_390074 ; 
   reg __390074_390074;
   reg _390075_390075 ; 
   reg __390075_390075;
   reg _390076_390076 ; 
   reg __390076_390076;
   reg _390077_390077 ; 
   reg __390077_390077;
   reg _390078_390078 ; 
   reg __390078_390078;
   reg _390079_390079 ; 
   reg __390079_390079;
   reg _390080_390080 ; 
   reg __390080_390080;
   reg _390081_390081 ; 
   reg __390081_390081;
   reg _390082_390082 ; 
   reg __390082_390082;
   reg _390083_390083 ; 
   reg __390083_390083;
   reg _390084_390084 ; 
   reg __390084_390084;
   reg _390085_390085 ; 
   reg __390085_390085;
   reg _390086_390086 ; 
   reg __390086_390086;
   reg _390087_390087 ; 
   reg __390087_390087;
   reg _390088_390088 ; 
   reg __390088_390088;
   reg _390089_390089 ; 
   reg __390089_390089;
   reg _390090_390090 ; 
   reg __390090_390090;
   reg _390091_390091 ; 
   reg __390091_390091;
   reg _390092_390092 ; 
   reg __390092_390092;
   reg _390093_390093 ; 
   reg __390093_390093;
   reg _390094_390094 ; 
   reg __390094_390094;
   reg _390095_390095 ; 
   reg __390095_390095;
   reg _390096_390096 ; 
   reg __390096_390096;
   reg _390097_390097 ; 
   reg __390097_390097;
   reg _390098_390098 ; 
   reg __390098_390098;
   reg _390099_390099 ; 
   reg __390099_390099;
   reg _390100_390100 ; 
   reg __390100_390100;
   reg _390101_390101 ; 
   reg __390101_390101;
   reg _390102_390102 ; 
   reg __390102_390102;
   reg _390103_390103 ; 
   reg __390103_390103;
   reg _390104_390104 ; 
   reg __390104_390104;
   reg _390105_390105 ; 
   reg __390105_390105;
   reg _390106_390106 ; 
   reg __390106_390106;
   reg _390107_390107 ; 
   reg __390107_390107;
   reg _390108_390108 ; 
   reg __390108_390108;
   reg _390109_390109 ; 
   reg __390109_390109;
   reg _390110_390110 ; 
   reg __390110_390110;
   reg _390111_390111 ; 
   reg __390111_390111;
   reg _390112_390112 ; 
   reg __390112_390112;
   reg _390113_390113 ; 
   reg __390113_390113;
   reg _390114_390114 ; 
   reg __390114_390114;
   reg _390115_390115 ; 
   reg __390115_390115;
   reg _390116_390116 ; 
   reg __390116_390116;
   reg _390117_390117 ; 
   reg __390117_390117;
   reg _390118_390118 ; 
   reg __390118_390118;
   reg _390119_390119 ; 
   reg __390119_390119;
   reg _390120_390120 ; 
   reg __390120_390120;
   reg _390121_390121 ; 
   reg __390121_390121;
   reg _390122_390122 ; 
   reg __390122_390122;
   reg _390123_390123 ; 
   reg __390123_390123;
   reg _390124_390124 ; 
   reg __390124_390124;
   reg _390125_390125 ; 
   reg __390125_390125;
   reg _390126_390126 ; 
   reg __390126_390126;
   reg _390127_390127 ; 
   reg __390127_390127;
   reg _390128_390128 ; 
   reg __390128_390128;
   reg _390129_390129 ; 
   reg __390129_390129;
   reg _390130_390130 ; 
   reg __390130_390130;
   reg _390131_390131 ; 
   reg __390131_390131;
   reg _390132_390132 ; 
   reg __390132_390132;
   reg _390133_390133 ; 
   reg __390133_390133;
   reg _390134_390134 ; 
   reg __390134_390134;
   reg _390135_390135 ; 
   reg __390135_390135;
   reg _390136_390136 ; 
   reg __390136_390136;
   reg _390137_390137 ; 
   reg __390137_390137;
   reg _390138_390138 ; 
   reg __390138_390138;
   reg _390139_390139 ; 
   reg __390139_390139;
   reg _390140_390140 ; 
   reg __390140_390140;
   reg _390141_390141 ; 
   reg __390141_390141;
   reg _390142_390142 ; 
   reg __390142_390142;
   reg _390143_390143 ; 
   reg __390143_390143;
   reg _390144_390144 ; 
   reg __390144_390144;
   reg _390145_390145 ; 
   reg __390145_390145;
   reg _390146_390146 ; 
   reg __390146_390146;
   reg _390147_390147 ; 
   reg __390147_390147;
   reg _390148_390148 ; 
   reg __390148_390148;
   reg _390149_390149 ; 
   reg __390149_390149;
   reg _390150_390150 ; 
   reg __390150_390150;
   reg _390151_390151 ; 
   reg __390151_390151;
   reg _390152_390152 ; 
   reg __390152_390152;
   reg _390153_390153 ; 
   reg __390153_390153;
   reg _390154_390154 ; 
   reg __390154_390154;
   reg _390155_390155 ; 
   reg __390155_390155;
   reg _390156_390156 ; 
   reg __390156_390156;
   reg _390157_390157 ; 
   reg __390157_390157;
   reg _390158_390158 ; 
   reg __390158_390158;
   reg _390159_390159 ; 
   reg __390159_390159;
   reg _390160_390160 ; 
   reg __390160_390160;
   reg _390161_390161 ; 
   reg __390161_390161;
   reg _390162_390162 ; 
   reg __390162_390162;
   reg _390163_390163 ; 
   reg __390163_390163;
   reg _390164_390164 ; 
   reg __390164_390164;
   reg _390165_390165 ; 
   reg __390165_390165;
   reg _390166_390166 ; 
   reg __390166_390166;
   reg _390167_390167 ; 
   reg __390167_390167;
   reg _390168_390168 ; 
   reg __390168_390168;
   reg _390169_390169 ; 
   reg __390169_390169;
   reg _390170_390170 ; 
   reg __390170_390170;
   reg _390171_390171 ; 
   reg __390171_390171;
   reg _390172_390172 ; 
   reg __390172_390172;
   reg _390173_390173 ; 
   reg __390173_390173;
   reg _390174_390174 ; 
   reg __390174_390174;
   reg _390175_390175 ; 
   reg __390175_390175;
   reg _390176_390176 ; 
   reg __390176_390176;
   reg _390177_390177 ; 
   reg __390177_390177;
   reg _390178_390178 ; 
   reg __390178_390178;
   reg _390179_390179 ; 
   reg __390179_390179;
   reg _390180_390180 ; 
   reg __390180_390180;
   reg _390181_390181 ; 
   reg __390181_390181;
   reg _390182_390182 ; 
   reg __390182_390182;
   reg _390183_390183 ; 
   reg __390183_390183;
   reg _390184_390184 ; 
   reg __390184_390184;
   reg _390185_390185 ; 
   reg __390185_390185;
   reg _390186_390186 ; 
   reg __390186_390186;
   reg _390187_390187 ; 
   reg __390187_390187;
   reg _390188_390188 ; 
   reg __390188_390188;
   reg _390189_390189 ; 
   reg __390189_390189;
   reg _390190_390190 ; 
   reg __390190_390190;
   reg _390191_390191 ; 
   reg __390191_390191;
   reg _390192_390192 ; 
   reg __390192_390192;
   reg _390193_390193 ; 
   reg __390193_390193;
   reg _390194_390194 ; 
   reg __390194_390194;
   reg _390195_390195 ; 
   reg __390195_390195;
   reg _390196_390196 ; 
   reg __390196_390196;
   reg _390197_390197 ; 
   reg __390197_390197;
   reg _390198_390198 ; 
   reg __390198_390198;
   reg _390199_390199 ; 
   reg __390199_390199;
   reg _390200_390200 ; 
   reg __390200_390200;
   reg _390201_390201 ; 
   reg __390201_390201;
   reg _390202_390202 ; 
   reg __390202_390202;
   reg _390203_390203 ; 
   reg __390203_390203;
   reg _390204_390204 ; 
   reg __390204_390204;
   reg _390205_390205 ; 
   reg __390205_390205;
   reg _390206_390206 ; 
   reg __390206_390206;
   reg _390207_390207 ; 
   reg __390207_390207;
   reg _390208_390208 ; 
   reg __390208_390208;
   reg _390209_390209 ; 
   reg __390209_390209;
   reg _390210_390210 ; 
   reg __390210_390210;
   reg _390211_390211 ; 
   reg __390211_390211;
   reg _390212_390212 ; 
   reg __390212_390212;
   reg _390213_390213 ; 
   reg __390213_390213;
   reg _390214_390214 ; 
   reg __390214_390214;
   reg _390215_390215 ; 
   reg __390215_390215;
   reg _390216_390216 ; 
   reg __390216_390216;
   reg _390217_390217 ; 
   reg __390217_390217;
   reg _390218_390218 ; 
   reg __390218_390218;
   reg _390219_390219 ; 
   reg __390219_390219;
   reg _390220_390220 ; 
   reg __390220_390220;
   reg _390221_390221 ; 
   reg __390221_390221;
   reg _390222_390222 ; 
   reg __390222_390222;
   reg _390223_390223 ; 
   reg __390223_390223;
   reg _390224_390224 ; 
   reg __390224_390224;
   reg _390225_390225 ; 
   reg __390225_390225;
   reg _390226_390226 ; 
   reg __390226_390226;
   reg _390227_390227 ; 
   reg __390227_390227;
   reg _390228_390228 ; 
   reg __390228_390228;
   reg _390229_390229 ; 
   reg __390229_390229;
   reg _390230_390230 ; 
   reg __390230_390230;
   reg _390231_390231 ; 
   reg __390231_390231;
   reg _390232_390232 ; 
   reg __390232_390232;
   reg _390233_390233 ; 
   reg __390233_390233;
   reg _390234_390234 ; 
   reg __390234_390234;
   reg _390235_390235 ; 
   reg __390235_390235;
   reg _390236_390236 ; 
   reg __390236_390236;
   reg _390237_390237 ; 
   reg __390237_390237;
   reg _390238_390238 ; 
   reg __390238_390238;
   reg _390239_390239 ; 
   reg __390239_390239;
   reg _390240_390240 ; 
   reg __390240_390240;
   reg _390241_390241 ; 
   reg __390241_390241;
   reg _390242_390242 ; 
   reg __390242_390242;
   reg _390243_390243 ; 
   reg __390243_390243;
   reg _390244_390244 ; 
   reg __390244_390244;
   reg _390245_390245 ; 
   reg __390245_390245;
   reg _390246_390246 ; 
   reg __390246_390246;
   reg _390247_390247 ; 
   reg __390247_390247;
   reg _390248_390248 ; 
   reg __390248_390248;
   reg _390249_390249 ; 
   reg __390249_390249;
   reg _390250_390250 ; 
   reg __390250_390250;
   reg _390251_390251 ; 
   reg __390251_390251;
   reg _390252_390252 ; 
   reg __390252_390252;
   reg _390253_390253 ; 
   reg __390253_390253;
   reg _390254_390254 ; 
   reg __390254_390254;
   reg _390255_390255 ; 
   reg __390255_390255;
   reg _390256_390256 ; 
   reg __390256_390256;
   reg _390257_390257 ; 
   reg __390257_390257;
   reg _390258_390258 ; 
   reg __390258_390258;
   reg _390259_390259 ; 
   reg __390259_390259;
   reg _390260_390260 ; 
   reg __390260_390260;
   reg _390261_390261 ; 
   reg __390261_390261;
   reg _390262_390262 ; 
   reg __390262_390262;
   reg _390263_390263 ; 
   reg __390263_390263;
   reg _390264_390264 ; 
   reg __390264_390264;
   reg _390265_390265 ; 
   reg __390265_390265;
   reg _390266_390266 ; 
   reg __390266_390266;
   reg _390267_390267 ; 
   reg __390267_390267;
   reg _390268_390268 ; 
   reg __390268_390268;
   reg _390269_390269 ; 
   reg __390269_390269;
   reg _390270_390270 ; 
   reg __390270_390270;
   reg _390271_390271 ; 
   reg __390271_390271;
   reg _390272_390272 ; 
   reg __390272_390272;
   reg _390273_390273 ; 
   reg __390273_390273;
   reg _390274_390274 ; 
   reg __390274_390274;
   reg _390275_390275 ; 
   reg __390275_390275;
   reg _390276_390276 ; 
   reg __390276_390276;
   reg _390277_390277 ; 
   reg __390277_390277;
   reg _390278_390278 ; 
   reg __390278_390278;
   reg _390279_390279 ; 
   reg __390279_390279;
   reg _390280_390280 ; 
   reg __390280_390280;
   reg _390281_390281 ; 
   reg __390281_390281;
   reg _390282_390282 ; 
   reg __390282_390282;
   reg _390283_390283 ; 
   reg __390283_390283;
   reg _390284_390284 ; 
   reg __390284_390284;
   reg _390285_390285 ; 
   reg __390285_390285;
   reg _390286_390286 ; 
   reg __390286_390286;
   reg _390287_390287 ; 
   reg __390287_390287;
   reg _390288_390288 ; 
   reg __390288_390288;
   reg _390289_390289 ; 
   reg __390289_390289;
   reg _390290_390290 ; 
   reg __390290_390290;
   reg _390291_390291 ; 
   reg __390291_390291;
   reg _390292_390292 ; 
   reg __390292_390292;
   reg _390293_390293 ; 
   reg __390293_390293;
   reg _390294_390294 ; 
   reg __390294_390294;
   reg _390295_390295 ; 
   reg __390295_390295;
   reg _390296_390296 ; 
   reg __390296_390296;
   reg _390297_390297 ; 
   reg __390297_390297;
   reg _390298_390298 ; 
   reg __390298_390298;
   reg _390299_390299 ; 
   reg __390299_390299;
   reg _390300_390300 ; 
   reg __390300_390300;
   reg _390301_390301 ; 
   reg __390301_390301;
   reg _390302_390302 ; 
   reg __390302_390302;
   reg _390303_390303 ; 
   reg __390303_390303;
   reg _390304_390304 ; 
   reg __390304_390304;
   reg _390305_390305 ; 
   reg __390305_390305;
   reg _390306_390306 ; 
   reg __390306_390306;
   reg _390307_390307 ; 
   reg __390307_390307;
   reg _390308_390308 ; 
   reg __390308_390308;
   reg _390309_390309 ; 
   reg __390309_390309;
   reg _390310_390310 ; 
   reg __390310_390310;
   reg _390311_390311 ; 
   reg __390311_390311;
   reg _390312_390312 ; 
   reg __390312_390312;
   reg _390313_390313 ; 
   reg __390313_390313;
   reg _390314_390314 ; 
   reg __390314_390314;
   reg _390315_390315 ; 
   reg __390315_390315;
   reg _390316_390316 ; 
   reg __390316_390316;
   reg _390317_390317 ; 
   reg __390317_390317;
   reg _390318_390318 ; 
   reg __390318_390318;
   reg _390319_390319 ; 
   reg __390319_390319;
   reg _390320_390320 ; 
   reg __390320_390320;
   reg _390321_390321 ; 
   reg __390321_390321;
   reg _390322_390322 ; 
   reg __390322_390322;
   reg _390323_390323 ; 
   reg __390323_390323;
   reg _390324_390324 ; 
   reg __390324_390324;
   reg _390325_390325 ; 
   reg __390325_390325;
   reg _390326_390326 ; 
   reg __390326_390326;
   reg _390327_390327 ; 
   reg __390327_390327;
   reg _390328_390328 ; 
   reg __390328_390328;
   reg _390329_390329 ; 
   reg __390329_390329;
   reg _390330_390330 ; 
   reg __390330_390330;
   reg _390331_390331 ; 
   reg __390331_390331;
   reg _390332_390332 ; 
   reg __390332_390332;
   reg _390333_390333 ; 
   reg __390333_390333;
   reg _390334_390334 ; 
   reg __390334_390334;
   reg _390335_390335 ; 
   reg __390335_390335;
   reg _390336_390336 ; 
   reg __390336_390336;
   reg _390337_390337 ; 
   reg __390337_390337;
   reg _390338_390338 ; 
   reg __390338_390338;
   reg _390339_390339 ; 
   reg __390339_390339;
   reg _390340_390340 ; 
   reg __390340_390340;
   reg _390341_390341 ; 
   reg __390341_390341;
   reg _390342_390342 ; 
   reg __390342_390342;
   reg _390343_390343 ; 
   reg __390343_390343;
   reg _390344_390344 ; 
   reg __390344_390344;
   reg _390345_390345 ; 
   reg __390345_390345;
   reg _390346_390346 ; 
   reg __390346_390346;
   reg _390347_390347 ; 
   reg __390347_390347;
   reg _390348_390348 ; 
   reg __390348_390348;
   reg _390349_390349 ; 
   reg __390349_390349;
   reg _390350_390350 ; 
   reg __390350_390350;
   reg _390351_390351 ; 
   reg __390351_390351;
   reg _390352_390352 ; 
   reg __390352_390352;
   reg _390353_390353 ; 
   reg __390353_390353;
   reg _390354_390354 ; 
   reg __390354_390354;
   reg _390355_390355 ; 
   reg __390355_390355;
   reg _390356_390356 ; 
   reg __390356_390356;
   reg _390357_390357 ; 
   reg __390357_390357;
   reg _390358_390358 ; 
   reg __390358_390358;
   reg _390359_390359 ; 
   reg __390359_390359;
   reg _390360_390360 ; 
   reg __390360_390360;
   reg _390361_390361 ; 
   reg __390361_390361;
   reg _390362_390362 ; 
   reg __390362_390362;
   reg _390363_390363 ; 
   reg __390363_390363;
   reg _390364_390364 ; 
   reg __390364_390364;
   reg _390365_390365 ; 
   reg __390365_390365;
   reg _390366_390366 ; 
   reg __390366_390366;
   reg _390367_390367 ; 
   reg __390367_390367;
   reg _390368_390368 ; 
   reg __390368_390368;
   reg _390369_390369 ; 
   reg __390369_390369;
   reg _390370_390370 ; 
   reg __390370_390370;
   reg _390371_390371 ; 
   reg __390371_390371;
   reg _390372_390372 ; 
   reg __390372_390372;
   reg _390373_390373 ; 
   reg __390373_390373;
   reg _390374_390374 ; 
   reg __390374_390374;
   reg _390375_390375 ; 
   reg __390375_390375;
   reg _390376_390376 ; 
   reg __390376_390376;
   reg _390377_390377 ; 
   reg __390377_390377;
   reg _390378_390378 ; 
   reg __390378_390378;
   reg _390379_390379 ; 
   reg __390379_390379;
   reg _390380_390380 ; 
   reg __390380_390380;
   reg _390381_390381 ; 
   reg __390381_390381;
   reg _390382_390382 ; 
   reg __390382_390382;
   reg _390383_390383 ; 
   reg __390383_390383;
   reg _390384_390384 ; 
   reg __390384_390384;
   reg _390385_390385 ; 
   reg __390385_390385;
   reg _390386_390386 ; 
   reg __390386_390386;
   reg _390387_390387 ; 
   reg __390387_390387;
   reg _390388_390388 ; 
   reg __390388_390388;
   reg _390389_390389 ; 
   reg __390389_390389;
   reg _390390_390390 ; 
   reg __390390_390390;
   reg _390391_390391 ; 
   reg __390391_390391;
   reg _390392_390392 ; 
   reg __390392_390392;
   reg _390393_390393 ; 
   reg __390393_390393;
   reg _390394_390394 ; 
   reg __390394_390394;
   reg _390395_390395 ; 
   reg __390395_390395;
   reg _390396_390396 ; 
   reg __390396_390396;
   reg _390397_390397 ; 
   reg __390397_390397;
   reg _390398_390398 ; 
   reg __390398_390398;
   reg _390399_390399 ; 
   reg __390399_390399;
   reg _390400_390400 ; 
   reg __390400_390400;
   reg _390401_390401 ; 
   reg __390401_390401;
   reg _390402_390402 ; 
   reg __390402_390402;
   reg _390403_390403 ; 
   reg __390403_390403;
   reg _390404_390404 ; 
   reg __390404_390404;
   reg _390405_390405 ; 
   reg __390405_390405;
   reg _390406_390406 ; 
   reg __390406_390406;
   reg _390407_390407 ; 
   reg __390407_390407;
   reg _390408_390408 ; 
   reg __390408_390408;
   reg _390409_390409 ; 
   reg __390409_390409;
   reg _390410_390410 ; 
   reg __390410_390410;
   reg _390411_390411 ; 
   reg __390411_390411;
   reg _390412_390412 ; 
   reg __390412_390412;
   reg _390413_390413 ; 
   reg __390413_390413;
   reg _390414_390414 ; 
   reg __390414_390414;
   reg _390415_390415 ; 
   reg __390415_390415;
   reg _390416_390416 ; 
   reg __390416_390416;
   reg _390417_390417 ; 
   reg __390417_390417;
   reg _390418_390418 ; 
   reg __390418_390418;
   reg _390419_390419 ; 
   reg __390419_390419;
   reg _390420_390420 ; 
   reg __390420_390420;
   reg _390421_390421 ; 
   reg __390421_390421;
   reg _390422_390422 ; 
   reg __390422_390422;
   reg _390423_390423 ; 
   reg __390423_390423;
   reg _390424_390424 ; 
   reg __390424_390424;
   reg _390425_390425 ; 
   reg __390425_390425;
   reg _390426_390426 ; 
   reg __390426_390426;
   reg _390427_390427 ; 
   reg __390427_390427;
   reg _390428_390428 ; 
   reg __390428_390428;
   reg _390429_390429 ; 
   reg __390429_390429;
   reg _390430_390430 ; 
   reg __390430_390430;
   reg _390431_390431 ; 
   reg __390431_390431;
   reg _390432_390432 ; 
   reg __390432_390432;
   reg _390433_390433 ; 
   reg __390433_390433;
   reg _390434_390434 ; 
   reg __390434_390434;
   reg _390435_390435 ; 
   reg __390435_390435;
   reg _390436_390436 ; 
   reg __390436_390436;
   reg _390437_390437 ; 
   reg __390437_390437;
   reg _390438_390438 ; 
   reg __390438_390438;
   reg _390439_390439 ; 
   reg __390439_390439;
   reg _390440_390440 ; 
   reg __390440_390440;
   reg _390441_390441 ; 
   reg __390441_390441;
   reg _390442_390442 ; 
   reg __390442_390442;
   reg _390443_390443 ; 
   reg __390443_390443;
   reg _390444_390444 ; 
   reg __390444_390444;
   reg _390445_390445 ; 
   reg __390445_390445;
   reg _390446_390446 ; 
   reg __390446_390446;
   reg _390447_390447 ; 
   reg __390447_390447;
   reg _390448_390448 ; 
   reg __390448_390448;
   reg _390449_390449 ; 
   reg __390449_390449;
   reg _390450_390450 ; 
   reg __390450_390450;
   reg _390451_390451 ; 
   reg __390451_390451;
   reg _390452_390452 ; 
   reg __390452_390452;
   reg _390453_390453 ; 
   reg __390453_390453;
   reg _390454_390454 ; 
   reg __390454_390454;
   reg _390455_390455 ; 
   reg __390455_390455;
   reg _390456_390456 ; 
   reg __390456_390456;
   reg _390457_390457 ; 
   reg __390457_390457;
   reg _390458_390458 ; 
   reg __390458_390458;
   reg _390459_390459 ; 
   reg __390459_390459;
   reg _390460_390460 ; 
   reg __390460_390460;
   reg _390461_390461 ; 
   reg __390461_390461;
   reg _390462_390462 ; 
   reg __390462_390462;
   reg _390463_390463 ; 
   reg __390463_390463;
   reg _390464_390464 ; 
   reg __390464_390464;
   reg _390465_390465 ; 
   reg __390465_390465;
   reg _390466_390466 ; 
   reg __390466_390466;
   reg _390467_390467 ; 
   reg __390467_390467;
   reg _390468_390468 ; 
   reg __390468_390468;
   reg _390469_390469 ; 
   reg __390469_390469;
   reg _390470_390470 ; 
   reg __390470_390470;
   reg _390471_390471 ; 
   reg __390471_390471;
   reg _390472_390472 ; 
   reg __390472_390472;
   reg _390473_390473 ; 
   reg __390473_390473;
   reg _390474_390474 ; 
   reg __390474_390474;
   reg _390475_390475 ; 
   reg __390475_390475;
   reg _390476_390476 ; 
   reg __390476_390476;
   reg _390477_390477 ; 
   reg __390477_390477;
   reg _390478_390478 ; 
   reg __390478_390478;
   reg _390479_390479 ; 
   reg __390479_390479;
   reg _390480_390480 ; 
   reg __390480_390480;
   reg _390481_390481 ; 
   reg __390481_390481;
   reg _390482_390482 ; 
   reg __390482_390482;
   reg _390483_390483 ; 
   reg __390483_390483;
   reg _390484_390484 ; 
   reg __390484_390484;
   reg _390485_390485 ; 
   reg __390485_390485;
   reg _390486_390486 ; 
   reg __390486_390486;
   reg _390487_390487 ; 
   reg __390487_390487;
   reg _390488_390488 ; 
   reg __390488_390488;
   reg _390489_390489 ; 
   reg __390489_390489;
   reg _390490_390490 ; 
   reg __390490_390490;
   reg _390491_390491 ; 
   reg __390491_390491;
   reg _390492_390492 ; 
   reg __390492_390492;
   reg _390493_390493 ; 
   reg __390493_390493;
   reg _390494_390494 ; 
   reg __390494_390494;
   reg _390495_390495 ; 
   reg __390495_390495;
   reg _390496_390496 ; 
   reg __390496_390496;
   reg _390497_390497 ; 
   reg __390497_390497;
   reg _390498_390498 ; 
   reg __390498_390498;
   reg _390499_390499 ; 
   reg __390499_390499;
   reg _390500_390500 ; 
   reg __390500_390500;
   reg _390501_390501 ; 
   reg __390501_390501;
   reg _390502_390502 ; 
   reg __390502_390502;
   reg _390503_390503 ; 
   reg __390503_390503;
   reg _390504_390504 ; 
   reg __390504_390504;
   reg _390505_390505 ; 
   reg __390505_390505;
   reg _390506_390506 ; 
   reg __390506_390506;
   reg _390507_390507 ; 
   reg __390507_390507;
   reg _390508_390508 ; 
   reg __390508_390508;
   reg _390509_390509 ; 
   reg __390509_390509;
   reg _390510_390510 ; 
   reg __390510_390510;
   reg _390511_390511 ; 
   reg __390511_390511;
   reg _390512_390512 ; 
   reg __390512_390512;
   reg _390513_390513 ; 
   reg __390513_390513;
   reg _390514_390514 ; 
   reg __390514_390514;
   reg _390515_390515 ; 
   reg __390515_390515;
   reg _390516_390516 ; 
   reg __390516_390516;
   reg _390517_390517 ; 
   reg __390517_390517;
   reg _390518_390518 ; 
   reg __390518_390518;
   reg _390519_390519 ; 
   reg __390519_390519;
   reg _390520_390520 ; 
   reg __390520_390520;
   reg _390521_390521 ; 
   reg __390521_390521;
   reg _390522_390522 ; 
   reg __390522_390522;
   reg _390523_390523 ; 
   reg __390523_390523;
   reg _390524_390524 ; 
   reg __390524_390524;
   reg _390525_390525 ; 
   reg __390525_390525;
   reg _390526_390526 ; 
   reg __390526_390526;
   reg _390527_390527 ; 
   reg __390527_390527;
   reg _390528_390528 ; 
   reg __390528_390528;
   reg _390529_390529 ; 
   reg __390529_390529;
   reg _390530_390530 ; 
   reg __390530_390530;
   reg _390531_390531 ; 
   reg __390531_390531;
   reg _390532_390532 ; 
   reg __390532_390532;
   reg _390533_390533 ; 
   reg __390533_390533;
   reg _390534_390534 ; 
   reg __390534_390534;
   reg _390535_390535 ; 
   reg __390535_390535;
   reg _390536_390536 ; 
   reg __390536_390536;
   reg _390537_390537 ; 
   reg __390537_390537;
   reg _390538_390538 ; 
   reg __390538_390538;
   reg _390539_390539 ; 
   reg __390539_390539;
   reg _390540_390540 ; 
   reg __390540_390540;
   reg _390541_390541 ; 
   reg __390541_390541;
   reg _390542_390542 ; 
   reg __390542_390542;
   reg _390543_390543 ; 
   reg __390543_390543;
   reg _390544_390544 ; 
   reg __390544_390544;
   reg _390545_390545 ; 
   reg __390545_390545;
   reg _390546_390546 ; 
   reg __390546_390546;
   reg _390547_390547 ; 
   reg __390547_390547;
   reg _390548_390548 ; 
   reg __390548_390548;
   reg _390549_390549 ; 
   reg __390549_390549;
   reg _390550_390550 ; 
   reg __390550_390550;
   reg _390551_390551 ; 
   reg __390551_390551;
   reg _390552_390552 ; 
   reg __390552_390552;
   reg _390553_390553 ; 
   reg __390553_390553;
   reg _390554_390554 ; 
   reg __390554_390554;
   reg _390555_390555 ; 
   reg __390555_390555;
   reg _390556_390556 ; 
   reg __390556_390556;
   reg _390557_390557 ; 
   reg __390557_390557;
   reg _390558_390558 ; 
   reg __390558_390558;
   reg _390559_390559 ; 
   reg __390559_390559;
   reg _390560_390560 ; 
   reg __390560_390560;
   reg _390561_390561 ; 
   reg __390561_390561;
   reg _390562_390562 ; 
   reg __390562_390562;
   reg _390563_390563 ; 
   reg __390563_390563;
   reg _390564_390564 ; 
   reg __390564_390564;
   reg _390565_390565 ; 
   reg __390565_390565;
   reg _390566_390566 ; 
   reg __390566_390566;
   reg _390567_390567 ; 
   reg __390567_390567;
   reg _390568_390568 ; 
   reg __390568_390568;
   reg _390569_390569 ; 
   reg __390569_390569;
   reg _390570_390570 ; 
   reg __390570_390570;
   reg _390571_390571 ; 
   reg __390571_390571;
   reg _390572_390572 ; 
   reg __390572_390572;
   reg _390573_390573 ; 
   reg __390573_390573;
   reg _390574_390574 ; 
   reg __390574_390574;
   reg _390575_390575 ; 
   reg __390575_390575;
   reg _390576_390576 ; 
   reg __390576_390576;
   reg _390577_390577 ; 
   reg __390577_390577;
   reg _390578_390578 ; 
   reg __390578_390578;
   reg _390579_390579 ; 
   reg __390579_390579;
   reg _390580_390580 ; 
   reg __390580_390580;
   reg _390581_390581 ; 
   reg __390581_390581;
   reg _390582_390582 ; 
   reg __390582_390582;
   reg _390583_390583 ; 
   reg __390583_390583;
   reg _390584_390584 ; 
   reg __390584_390584;
   reg _390585_390585 ; 
   reg __390585_390585;
   reg _390586_390586 ; 
   reg __390586_390586;
   reg _390587_390587 ; 
   reg __390587_390587;
   reg _390588_390588 ; 
   reg __390588_390588;
   reg _390589_390589 ; 
   reg __390589_390589;
   reg _390590_390590 ; 
   reg __390590_390590;
   reg _390591_390591 ; 
   reg __390591_390591;
   reg _390592_390592 ; 
   reg __390592_390592;
   reg _390593_390593 ; 
   reg __390593_390593;
   reg _390594_390594 ; 
   reg __390594_390594;
   reg _390595_390595 ; 
   reg __390595_390595;
   reg _390596_390596 ; 
   reg __390596_390596;
   reg _390597_390597 ; 
   reg __390597_390597;
   reg _390598_390598 ; 
   reg __390598_390598;
   reg _390599_390599 ; 
   reg __390599_390599;
   reg _390600_390600 ; 
   reg __390600_390600;
   reg _390601_390601 ; 
   reg __390601_390601;
   reg _390602_390602 ; 
   reg __390602_390602;
   reg _390603_390603 ; 
   reg __390603_390603;
   reg _390604_390604 ; 
   reg __390604_390604;
   reg _390605_390605 ; 
   reg __390605_390605;
   reg _390606_390606 ; 
   reg __390606_390606;
   reg _390607_390607 ; 
   reg __390607_390607;
   reg _390608_390608 ; 
   reg __390608_390608;
   reg _390609_390609 ; 
   reg __390609_390609;
   reg _390610_390610 ; 
   reg __390610_390610;
   reg _390611_390611 ; 
   reg __390611_390611;
   reg _390612_390612 ; 
   reg __390612_390612;
   reg _390613_390613 ; 
   reg __390613_390613;
   reg _390614_390614 ; 
   reg __390614_390614;
   reg _390615_390615 ; 
   reg __390615_390615;
   reg _390616_390616 ; 
   reg __390616_390616;
   reg _390617_390617 ; 
   reg __390617_390617;
   reg _390618_390618 ; 
   reg __390618_390618;
   reg _390619_390619 ; 
   reg __390619_390619;
   reg _390620_390620 ; 
   reg __390620_390620;
   reg _390621_390621 ; 
   reg __390621_390621;
   reg _390622_390622 ; 
   reg __390622_390622;
   reg _390623_390623 ; 
   reg __390623_390623;
   reg _390624_390624 ; 
   reg __390624_390624;
   reg _390625_390625 ; 
   reg __390625_390625;
   reg _390626_390626 ; 
   reg __390626_390626;
   reg _390627_390627 ; 
   reg __390627_390627;
   reg _390628_390628 ; 
   reg __390628_390628;
   reg _390629_390629 ; 
   reg __390629_390629;
   reg _390630_390630 ; 
   reg __390630_390630;
   reg _390631_390631 ; 
   reg __390631_390631;
   reg _390632_390632 ; 
   reg __390632_390632;
   reg _390633_390633 ; 
   reg __390633_390633;
   reg _390634_390634 ; 
   reg __390634_390634;
   reg _390635_390635 ; 
   reg __390635_390635;
   reg _390636_390636 ; 
   reg __390636_390636;
   reg _390637_390637 ; 
   reg __390637_390637;
   reg _390638_390638 ; 
   reg __390638_390638;
   reg _390639_390639 ; 
   reg __390639_390639;
   reg _390640_390640 ; 
   reg __390640_390640;
   reg _390641_390641 ; 
   reg __390641_390641;
   reg _390642_390642 ; 
   reg __390642_390642;
   reg _390643_390643 ; 
   reg __390643_390643;
   reg _390644_390644 ; 
   reg __390644_390644;
   reg _390645_390645 ; 
   reg __390645_390645;
   reg _390646_390646 ; 
   reg __390646_390646;
   reg _390647_390647 ; 
   reg __390647_390647;
   reg _390648_390648 ; 
   reg __390648_390648;
   reg _390649_390649 ; 
   reg __390649_390649;
   reg _390650_390650 ; 
   reg __390650_390650;
   reg _390651_390651 ; 
   reg __390651_390651;
   reg _390652_390652 ; 
   reg __390652_390652;
   reg _390653_390653 ; 
   reg __390653_390653;
   reg _390654_390654 ; 
   reg __390654_390654;
   reg _390655_390655 ; 
   reg __390655_390655;
   reg _390656_390656 ; 
   reg __390656_390656;
   reg _390657_390657 ; 
   reg __390657_390657;
   reg _390658_390658 ; 
   reg __390658_390658;
   reg _390659_390659 ; 
   reg __390659_390659;
   reg _390660_390660 ; 
   reg __390660_390660;
   reg _390661_390661 ; 
   reg __390661_390661;
   reg _390662_390662 ; 
   reg __390662_390662;
   reg _390663_390663 ; 
   reg __390663_390663;
   reg _390664_390664 ; 
   reg __390664_390664;
   reg _390665_390665 ; 
   reg __390665_390665;
   reg _390666_390666 ; 
   reg __390666_390666;
   reg _390667_390667 ; 
   reg __390667_390667;
   reg _390668_390668 ; 
   reg __390668_390668;
   reg _390669_390669 ; 
   reg __390669_390669;
   reg _390670_390670 ; 
   reg __390670_390670;
   reg _390671_390671 ; 
   reg __390671_390671;
   reg _390672_390672 ; 
   reg __390672_390672;
   reg _390673_390673 ; 
   reg __390673_390673;
   reg _390674_390674 ; 
   reg __390674_390674;
   reg _390675_390675 ; 
   reg __390675_390675;
   reg _390676_390676 ; 
   reg __390676_390676;
   reg _390677_390677 ; 
   reg __390677_390677;
   reg _390678_390678 ; 
   reg __390678_390678;
   reg _390679_390679 ; 
   reg __390679_390679;
   reg _390680_390680 ; 
   reg __390680_390680;
   reg _390681_390681 ; 
   reg __390681_390681;
   reg _390682_390682 ; 
   reg __390682_390682;
   reg _390683_390683 ; 
   reg __390683_390683;
   reg _390684_390684 ; 
   reg __390684_390684;
   reg _390685_390685 ; 
   reg __390685_390685;
   reg _390686_390686 ; 
   reg __390686_390686;
   reg _390687_390687 ; 
   reg __390687_390687;
   reg _390688_390688 ; 
   reg __390688_390688;
   reg _390689_390689 ; 
   reg __390689_390689;
   reg _390690_390690 ; 
   reg __390690_390690;
   reg _390691_390691 ; 
   reg __390691_390691;
   reg _390692_390692 ; 
   reg __390692_390692;
   reg _390693_390693 ; 
   reg __390693_390693;
   reg _390694_390694 ; 
   reg __390694_390694;
   reg _390695_390695 ; 
   reg __390695_390695;
   reg _390696_390696 ; 
   reg __390696_390696;
   reg _390697_390697 ; 
   reg __390697_390697;
   reg _390698_390698 ; 
   reg __390698_390698;
   reg _390699_390699 ; 
   reg __390699_390699;
   reg _390700_390700 ; 
   reg __390700_390700;
   reg _390701_390701 ; 
   reg __390701_390701;
   reg _390702_390702 ; 
   reg __390702_390702;
   reg _390703_390703 ; 
   reg __390703_390703;
   reg _390704_390704 ; 
   reg __390704_390704;
   reg _390705_390705 ; 
   reg __390705_390705;
   reg _390706_390706 ; 
   reg __390706_390706;
   reg _390707_390707 ; 
   reg __390707_390707;
   reg _390708_390708 ; 
   reg __390708_390708;
   reg _390709_390709 ; 
   reg __390709_390709;
   reg _390710_390710 ; 
   reg __390710_390710;
   reg _390711_390711 ; 
   reg __390711_390711;
   reg _390712_390712 ; 
   reg __390712_390712;
   reg _390713_390713 ; 
   reg __390713_390713;
   reg _390714_390714 ; 
   reg __390714_390714;
   reg _390715_390715 ; 
   reg __390715_390715;
   reg _390716_390716 ; 
   reg __390716_390716;
   reg _390717_390717 ; 
   reg __390717_390717;
   reg _390718_390718 ; 
   reg __390718_390718;
   reg _390719_390719 ; 
   reg __390719_390719;
   reg _390720_390720 ; 
   reg __390720_390720;
   reg _390721_390721 ; 
   reg __390721_390721;
   reg _390722_390722 ; 
   reg __390722_390722;
   reg _390723_390723 ; 
   reg __390723_390723;
   reg _390724_390724 ; 
   reg __390724_390724;
   reg _390725_390725 ; 
   reg __390725_390725;
   reg _390726_390726 ; 
   reg __390726_390726;
   reg _390727_390727 ; 
   reg __390727_390727;
   reg _390728_390728 ; 
   reg __390728_390728;
   reg _390729_390729 ; 
   reg __390729_390729;
   reg _390730_390730 ; 
   reg __390730_390730;
   reg _390731_390731 ; 
   reg __390731_390731;
   reg _390732_390732 ; 
   reg __390732_390732;
   reg _390733_390733 ; 
   reg __390733_390733;
   reg _390734_390734 ; 
   reg __390734_390734;
   reg _390735_390735 ; 
   reg __390735_390735;
   reg _390736_390736 ; 
   reg __390736_390736;
   reg _390737_390737 ; 
   reg __390737_390737;
   reg _390738_390738 ; 
   reg __390738_390738;
   reg _390739_390739 ; 
   reg __390739_390739;
   reg _390740_390740 ; 
   reg __390740_390740;
   reg _390741_390741 ; 
   reg __390741_390741;
   reg _390742_390742 ; 
   reg __390742_390742;
   reg _390743_390743 ; 
   reg __390743_390743;
   reg _390744_390744 ; 
   reg __390744_390744;
   reg _390745_390745 ; 
   reg __390745_390745;
   reg _390746_390746 ; 
   reg __390746_390746;
   reg _390747_390747 ; 
   reg __390747_390747;
   reg _390748_390748 ; 
   reg __390748_390748;
   reg _390749_390749 ; 
   reg __390749_390749;
   reg _390750_390750 ; 
   reg __390750_390750;
   reg _390751_390751 ; 
   reg __390751_390751;
   reg _390752_390752 ; 
   reg __390752_390752;
   reg _390753_390753 ; 
   reg __390753_390753;
   reg _390754_390754 ; 
   reg __390754_390754;
   reg _390755_390755 ; 
   reg __390755_390755;
   reg _390756_390756 ; 
   reg __390756_390756;
   reg _390757_390757 ; 
   reg __390757_390757;
   reg _390758_390758 ; 
   reg __390758_390758;
   reg _390759_390759 ; 
   reg __390759_390759;
   reg _390760_390760 ; 
   reg __390760_390760;
   reg _390761_390761 ; 
   reg __390761_390761;
   reg _390762_390762 ; 
   reg __390762_390762;
   reg _390763_390763 ; 
   reg __390763_390763;
   reg _390764_390764 ; 
   reg __390764_390764;
   reg _390765_390765 ; 
   reg __390765_390765;
   reg _390766_390766 ; 
   reg __390766_390766;
   reg _390767_390767 ; 
   reg __390767_390767;
   reg _390768_390768 ; 
   reg __390768_390768;
   reg _390769_390769 ; 
   reg __390769_390769;
   reg _390770_390770 ; 
   reg __390770_390770;
   reg _390771_390771 ; 
   reg __390771_390771;
   reg _390772_390772 ; 
   reg __390772_390772;
   reg _390773_390773 ; 
   reg __390773_390773;
   reg _390774_390774 ; 
   reg __390774_390774;
   reg _390775_390775 ; 
   reg __390775_390775;
   reg _390776_390776 ; 
   reg __390776_390776;
   reg _390777_390777 ; 
   reg __390777_390777;
   reg _390778_390778 ; 
   reg __390778_390778;
   reg _390779_390779 ; 
   reg __390779_390779;
   reg _390780_390780 ; 
   reg __390780_390780;
   reg _390781_390781 ; 
   reg __390781_390781;
   reg _390782_390782 ; 
   reg __390782_390782;
   reg _390783_390783 ; 
   reg __390783_390783;
   reg _390784_390784 ; 
   reg __390784_390784;
   reg _390785_390785 ; 
   reg __390785_390785;
   reg _390786_390786 ; 
   reg __390786_390786;
   reg _390787_390787 ; 
   reg __390787_390787;
   reg _390788_390788 ; 
   reg __390788_390788;
   reg _390789_390789 ; 
   reg __390789_390789;
   reg _390790_390790 ; 
   reg __390790_390790;
   reg _390791_390791 ; 
   reg __390791_390791;
   reg _390792_390792 ; 
   reg __390792_390792;
   reg _390793_390793 ; 
   reg __390793_390793;
   reg _390794_390794 ; 
   reg __390794_390794;
   reg _390795_390795 ; 
   reg __390795_390795;
   reg _390796_390796 ; 
   reg __390796_390796;
   reg _390797_390797 ; 
   reg __390797_390797;
   reg _390798_390798 ; 
   reg __390798_390798;
   reg _390799_390799 ; 
   reg __390799_390799;
   reg _390800_390800 ; 
   reg __390800_390800;
   reg _390801_390801 ; 
   reg __390801_390801;
   reg _390802_390802 ; 
   reg __390802_390802;
   reg _390803_390803 ; 
   reg __390803_390803;
   reg _390804_390804 ; 
   reg __390804_390804;
   reg _390805_390805 ; 
   reg __390805_390805;
   reg _390806_390806 ; 
   reg __390806_390806;
   reg _390807_390807 ; 
   reg __390807_390807;
   reg _390808_390808 ; 
   reg __390808_390808;
   reg _390809_390809 ; 
   reg __390809_390809;
   reg _390810_390810 ; 
   reg __390810_390810;
   reg _390811_390811 ; 
   reg __390811_390811;
   reg _390812_390812 ; 
   reg __390812_390812;
   reg _390813_390813 ; 
   reg __390813_390813;
   reg _390814_390814 ; 
   reg __390814_390814;
   reg _390815_390815 ; 
   reg __390815_390815;
   reg _390816_390816 ; 
   reg __390816_390816;
   reg _390817_390817 ; 
   reg __390817_390817;
   reg _390818_390818 ; 
   reg __390818_390818;
   reg _390819_390819 ; 
   reg __390819_390819;
   reg _390820_390820 ; 
   reg __390820_390820;
   reg _390821_390821 ; 
   reg __390821_390821;
   reg _390822_390822 ; 
   reg __390822_390822;
   reg _390823_390823 ; 
   reg __390823_390823;
   reg _390824_390824 ; 
   reg __390824_390824;
   reg _390825_390825 ; 
   reg __390825_390825;
   reg _390826_390826 ; 
   reg __390826_390826;
   reg _390827_390827 ; 
   reg __390827_390827;
   reg _390828_390828 ; 
   reg __390828_390828;
   reg _390829_390829 ; 
   reg __390829_390829;
   reg _390830_390830 ; 
   reg __390830_390830;
   reg _390831_390831 ; 
   reg __390831_390831;
   reg _390832_390832 ; 
   reg __390832_390832;
   reg _390833_390833 ; 
   reg __390833_390833;
   reg _390834_390834 ; 
   reg __390834_390834;
   reg _390835_390835 ; 
   reg __390835_390835;
   reg _390836_390836 ; 
   reg __390836_390836;
   reg _390837_390837 ; 
   reg __390837_390837;
   reg _390838_390838 ; 
   reg __390838_390838;
   reg _390839_390839 ; 
   reg __390839_390839;
   reg _390840_390840 ; 
   reg __390840_390840;
   reg _390841_390841 ; 
   reg __390841_390841;
   reg _390842_390842 ; 
   reg __390842_390842;
   reg _390843_390843 ; 
   reg __390843_390843;
   reg _390844_390844 ; 
   reg __390844_390844;
   reg _390845_390845 ; 
   reg __390845_390845;
   reg _390846_390846 ; 
   reg __390846_390846;
   reg _390847_390847 ; 
   reg __390847_390847;
   reg _390848_390848 ; 
   reg __390848_390848;
   reg _390849_390849 ; 
   reg __390849_390849;
   reg _390850_390850 ; 
   reg __390850_390850;
   reg _390851_390851 ; 
   reg __390851_390851;
   reg _390852_390852 ; 
   reg __390852_390852;
   reg _390853_390853 ; 
   reg __390853_390853;
   reg _390854_390854 ; 
   reg __390854_390854;
   reg _390855_390855 ; 
   reg __390855_390855;
   reg _390856_390856 ; 
   reg __390856_390856;
   reg _390857_390857 ; 
   reg __390857_390857;
   reg _390858_390858 ; 
   reg __390858_390858;
   reg _390859_390859 ; 
   reg __390859_390859;
   reg _390860_390860 ; 
   reg __390860_390860;
   reg _390861_390861 ; 
   reg __390861_390861;
   reg _390862_390862 ; 
   reg __390862_390862;
   reg _390863_390863 ; 
   reg __390863_390863;
   reg _390864_390864 ; 
   reg __390864_390864;
   reg _390865_390865 ; 
   reg __390865_390865;
   reg _390866_390866 ; 
   reg __390866_390866;
   reg _390867_390867 ; 
   reg __390867_390867;
   reg _390868_390868 ; 
   reg __390868_390868;
   reg _390869_390869 ; 
   reg __390869_390869;
   reg _390870_390870 ; 
   reg __390870_390870;
   reg _390871_390871 ; 
   reg __390871_390871;
   reg _390872_390872 ; 
   reg __390872_390872;
   reg _390873_390873 ; 
   reg __390873_390873;
   reg _390874_390874 ; 
   reg __390874_390874;
   reg _390875_390875 ; 
   reg __390875_390875;
   reg _390876_390876 ; 
   reg __390876_390876;
   reg _390877_390877 ; 
   reg __390877_390877;
   reg _390878_390878 ; 
   reg __390878_390878;
   reg _390879_390879 ; 
   reg __390879_390879;
   reg _390880_390880 ; 
   reg __390880_390880;
   reg _390881_390881 ; 
   reg __390881_390881;
   reg _390882_390882 ; 
   reg __390882_390882;
   reg _390883_390883 ; 
   reg __390883_390883;
   reg _390884_390884 ; 
   reg __390884_390884;
   reg _390885_390885 ; 
   reg __390885_390885;
   reg _390886_390886 ; 
   reg __390886_390886;
   reg _390887_390887 ; 
   reg __390887_390887;
   reg _390888_390888 ; 
   reg __390888_390888;
   reg _390889_390889 ; 
   reg __390889_390889;
   reg _390890_390890 ; 
   reg __390890_390890;
   reg _390891_390891 ; 
   reg __390891_390891;
   reg _390892_390892 ; 
   reg __390892_390892;
   reg _390893_390893 ; 
   reg __390893_390893;
   reg _390894_390894 ; 
   reg __390894_390894;
   reg _390895_390895 ; 
   reg __390895_390895;
   reg _390896_390896 ; 
   reg __390896_390896;
   reg _390897_390897 ; 
   reg __390897_390897;
   reg _390898_390898 ; 
   reg __390898_390898;
   reg _390899_390899 ; 
   reg __390899_390899;
   reg _390900_390900 ; 
   reg __390900_390900;
   reg _390901_390901 ; 
   reg __390901_390901;
   reg _390902_390902 ; 
   reg __390902_390902;
   reg _390903_390903 ; 
   reg __390903_390903;
   reg _390904_390904 ; 
   reg __390904_390904;
   reg _390905_390905 ; 
   reg __390905_390905;
   reg _390906_390906 ; 
   reg __390906_390906;
   reg _390907_390907 ; 
   reg __390907_390907;
   reg _390908_390908 ; 
   reg __390908_390908;
   reg _390909_390909 ; 
   reg __390909_390909;
   reg _390910_390910 ; 
   reg __390910_390910;
   reg _390911_390911 ; 
   reg __390911_390911;
   reg _390912_390912 ; 
   reg __390912_390912;
   reg _390913_390913 ; 
   reg __390913_390913;
   reg _390914_390914 ; 
   reg __390914_390914;
   reg _390915_390915 ; 
   reg __390915_390915;
   reg _390916_390916 ; 
   reg __390916_390916;
   reg _390917_390917 ; 
   reg __390917_390917;
   reg _390918_390918 ; 
   reg __390918_390918;
   reg _390919_390919 ; 
   reg __390919_390919;
   reg _390920_390920 ; 
   reg __390920_390920;
   reg _390921_390921 ; 
   reg __390921_390921;
   reg _390922_390922 ; 
   reg __390922_390922;
   reg _390923_390923 ; 
   reg __390923_390923;
   reg _390924_390924 ; 
   reg __390924_390924;
   reg _390925_390925 ; 
   reg __390925_390925;
   reg _390926_390926 ; 
   reg __390926_390926;
   reg _390927_390927 ; 
   reg __390927_390927;
   reg _390928_390928 ; 
   reg __390928_390928;
   reg _390929_390929 ; 
   reg __390929_390929;
   reg _390930_390930 ; 
   reg __390930_390930;
   reg _390931_390931 ; 
   reg __390931_390931;
   reg _390932_390932 ; 
   reg __390932_390932;
   reg _390933_390933 ; 
   reg __390933_390933;
   reg _390934_390934 ; 
   reg __390934_390934;
   reg _390935_390935 ; 
   reg __390935_390935;
   reg _390936_390936 ; 
   reg __390936_390936;
   reg _390937_390937 ; 
   reg __390937_390937;
   reg _390938_390938 ; 
   reg __390938_390938;
   reg _390939_390939 ; 
   reg __390939_390939;
   reg _390940_390940 ; 
   reg __390940_390940;
   reg _390941_390941 ; 
   reg __390941_390941;
   reg _390942_390942 ; 
   reg __390942_390942;
   reg _390943_390943 ; 
   reg __390943_390943;
   reg _390944_390944 ; 
   reg __390944_390944;
   reg _390945_390945 ; 
   reg __390945_390945;
   reg _390946_390946 ; 
   reg __390946_390946;
   reg _390947_390947 ; 
   reg __390947_390947;
   reg _390948_390948 ; 
   reg __390948_390948;
   reg _390949_390949 ; 
   reg __390949_390949;
   reg _390950_390950 ; 
   reg __390950_390950;
   reg _390951_390951 ; 
   reg __390951_390951;
   reg _390952_390952 ; 
   reg __390952_390952;
   reg _390953_390953 ; 
   reg __390953_390953;
   reg _390954_390954 ; 
   reg __390954_390954;
   reg _390955_390955 ; 
   reg __390955_390955;
   reg _390956_390956 ; 
   reg __390956_390956;
   reg _390957_390957 ; 
   reg __390957_390957;
   reg _390958_390958 ; 
   reg __390958_390958;
   reg _390959_390959 ; 
   reg __390959_390959;
   reg _390960_390960 ; 
   reg __390960_390960;
   reg _390961_390961 ; 
   reg __390961_390961;
   reg _390962_390962 ; 
   reg __390962_390962;
   reg _390963_390963 ; 
   reg __390963_390963;
   reg _390964_390964 ; 
   reg __390964_390964;
   reg _390965_390965 ; 
   reg __390965_390965;
   reg _390966_390966 ; 
   reg __390966_390966;
   reg _390967_390967 ; 
   reg __390967_390967;
   reg _390968_390968 ; 
   reg __390968_390968;
   reg _390969_390969 ; 
   reg __390969_390969;
   reg _390970_390970 ; 
   reg __390970_390970;
   reg _390971_390971 ; 
   reg __390971_390971;
   reg _390972_390972 ; 
   reg __390972_390972;
   reg _390973_390973 ; 
   reg __390973_390973;
   reg _390974_390974 ; 
   reg __390974_390974;
   reg _390975_390975 ; 
   reg __390975_390975;
   reg _390976_390976 ; 
   reg __390976_390976;
   reg _390977_390977 ; 
   reg __390977_390977;
   reg _390978_390978 ; 
   reg __390978_390978;
   reg _390979_390979 ; 
   reg __390979_390979;
   reg _390980_390980 ; 
   reg __390980_390980;
   reg _390981_390981 ; 
   reg __390981_390981;
   reg _390982_390982 ; 
   reg __390982_390982;
   reg _390983_390983 ; 
   reg __390983_390983;
   reg _390984_390984 ; 
   reg __390984_390984;
   reg _390985_390985 ; 
   reg __390985_390985;
   reg _390986_390986 ; 
   reg __390986_390986;
   reg _390987_390987 ; 
   reg __390987_390987;
   reg _390988_390988 ; 
   reg __390988_390988;
   reg _390989_390989 ; 
   reg __390989_390989;
   reg _390990_390990 ; 
   reg __390990_390990;
   reg _390991_390991 ; 
   reg __390991_390991;
   reg _390992_390992 ; 
   reg __390992_390992;
   reg _390993_390993 ; 
   reg __390993_390993;
   reg _390994_390994 ; 
   reg __390994_390994;
   reg _390995_390995 ; 
   reg __390995_390995;
   reg _390996_390996 ; 
   reg __390996_390996;
   reg _390997_390997 ; 
   reg __390997_390997;
   reg _390998_390998 ; 
   reg __390998_390998;
   reg _390999_390999 ; 
   reg __390999_390999;
   reg _391000_391000 ; 
   reg __391000_391000;
   reg _391001_391001 ; 
   reg __391001_391001;
   reg _391002_391002 ; 
   reg __391002_391002;
   reg _391003_391003 ; 
   reg __391003_391003;
   reg _391004_391004 ; 
   reg __391004_391004;
   reg _391005_391005 ; 
   reg __391005_391005;
   reg _391006_391006 ; 
   reg __391006_391006;
   reg _391007_391007 ; 
   reg __391007_391007;
   reg _391008_391008 ; 
   reg __391008_391008;
   reg _391009_391009 ; 
   reg __391009_391009;
   reg _391010_391010 ; 
   reg __391010_391010;
   reg _391011_391011 ; 
   reg __391011_391011;
   reg _391012_391012 ; 
   reg __391012_391012;
   reg _391013_391013 ; 
   reg __391013_391013;
   reg _391014_391014 ; 
   reg __391014_391014;
   reg _391015_391015 ; 
   reg __391015_391015;
   reg _391016_391016 ; 
   reg __391016_391016;
   reg _391017_391017 ; 
   reg __391017_391017;
   reg _391018_391018 ; 
   reg __391018_391018;
   reg _391019_391019 ; 
   reg __391019_391019;
   reg _391020_391020 ; 
   reg __391020_391020;
   reg _391021_391021 ; 
   reg __391021_391021;
   reg _391022_391022 ; 
   reg __391022_391022;
   reg _391023_391023 ; 
   reg __391023_391023;
   reg _391024_391024 ; 
   reg __391024_391024;
   reg _391025_391025 ; 
   reg __391025_391025;
   reg _391026_391026 ; 
   reg __391026_391026;
   reg _391027_391027 ; 
   reg __391027_391027;
   reg _391028_391028 ; 
   reg __391028_391028;
   reg _391029_391029 ; 
   reg __391029_391029;
   reg _391030_391030 ; 
   reg __391030_391030;
   reg _391031_391031 ; 
   reg __391031_391031;
   reg _391032_391032 ; 
   reg __391032_391032;
   reg _391033_391033 ; 
   reg __391033_391033;
   reg _391034_391034 ; 
   reg __391034_391034;
   reg _391035_391035 ; 
   reg __391035_391035;
   reg _391036_391036 ; 
   reg __391036_391036;
   reg _391037_391037 ; 
   reg __391037_391037;
   reg _391038_391038 ; 
   reg __391038_391038;
   reg _391039_391039 ; 
   reg __391039_391039;
   reg _391040_391040 ; 
   reg __391040_391040;
   reg _391041_391041 ; 
   reg __391041_391041;
   reg _391042_391042 ; 
   reg __391042_391042;
   reg _391043_391043 ; 
   reg __391043_391043;
   reg _391044_391044 ; 
   reg __391044_391044;
   reg _391045_391045 ; 
   reg __391045_391045;
   reg _391046_391046 ; 
   reg __391046_391046;
   reg _391047_391047 ; 
   reg __391047_391047;
   reg _391048_391048 ; 
   reg __391048_391048;
   reg _391049_391049 ; 
   reg __391049_391049;
   reg _391050_391050 ; 
   reg __391050_391050;
   reg _391051_391051 ; 
   reg __391051_391051;
   reg _391052_391052 ; 
   reg __391052_391052;
   reg _391053_391053 ; 
   reg __391053_391053;
   reg _391054_391054 ; 
   reg __391054_391054;
   reg _391055_391055 ; 
   reg __391055_391055;
   reg _391056_391056 ; 
   reg __391056_391056;
   reg _391057_391057 ; 
   reg __391057_391057;
   reg _391058_391058 ; 
   reg __391058_391058;
   reg _391059_391059 ; 
   reg __391059_391059;
   reg _391060_391060 ; 
   reg __391060_391060;
   reg _391061_391061 ; 
   reg __391061_391061;
   reg _391062_391062 ; 
   reg __391062_391062;
   reg _391063_391063 ; 
   reg __391063_391063;
   reg _391064_391064 ; 
   reg __391064_391064;
   reg _391065_391065 ; 
   reg __391065_391065;
   reg _391066_391066 ; 
   reg __391066_391066;
   reg _391067_391067 ; 
   reg __391067_391067;
   reg _391068_391068 ; 
   reg __391068_391068;
   reg _391069_391069 ; 
   reg __391069_391069;
   reg _391070_391070 ; 
   reg __391070_391070;
   reg _391071_391071 ; 
   reg __391071_391071;
   reg _391072_391072 ; 
   reg __391072_391072;
   reg _391073_391073 ; 
   reg __391073_391073;
   reg _391074_391074 ; 
   reg __391074_391074;
   reg _391075_391075 ; 
   reg __391075_391075;
   reg _391076_391076 ; 
   reg __391076_391076;
   reg _391077_391077 ; 
   reg __391077_391077;
   reg _391078_391078 ; 
   reg __391078_391078;
   reg _391079_391079 ; 
   reg __391079_391079;
   reg _391080_391080 ; 
   reg __391080_391080;
   reg _391081_391081 ; 
   reg __391081_391081;
   reg _391082_391082 ; 
   reg __391082_391082;
   reg _391083_391083 ; 
   reg __391083_391083;
   reg _391084_391084 ; 
   reg __391084_391084;
   reg _391085_391085 ; 
   reg __391085_391085;
   reg _391086_391086 ; 
   reg __391086_391086;
   reg _391087_391087 ; 
   reg __391087_391087;
   reg _391088_391088 ; 
   reg __391088_391088;
   reg _391089_391089 ; 
   reg __391089_391089;
   reg _391090_391090 ; 
   reg __391090_391090;
   reg _391091_391091 ; 
   reg __391091_391091;
   reg _391092_391092 ; 
   reg __391092_391092;
   reg _391093_391093 ; 
   reg __391093_391093;
   reg _391094_391094 ; 
   reg __391094_391094;
   reg _391095_391095 ; 
   reg __391095_391095;
   reg _391096_391096 ; 
   reg __391096_391096;
   reg _391097_391097 ; 
   reg __391097_391097;
   reg _391098_391098 ; 
   reg __391098_391098;
   reg _391099_391099 ; 
   reg __391099_391099;
   reg _391100_391100 ; 
   reg __391100_391100;
   reg _391101_391101 ; 
   reg __391101_391101;
   reg _391102_391102 ; 
   reg __391102_391102;
   reg _391103_391103 ; 
   reg __391103_391103;
   reg _391104_391104 ; 
   reg __391104_391104;
   reg _391105_391105 ; 
   reg __391105_391105;
   reg _391106_391106 ; 
   reg __391106_391106;
   reg _391107_391107 ; 
   reg __391107_391107;
   reg _391108_391108 ; 
   reg __391108_391108;
   reg _391109_391109 ; 
   reg __391109_391109;
   reg _391110_391110 ; 
   reg __391110_391110;
   reg _391111_391111 ; 
   reg __391111_391111;
   reg _391112_391112 ; 
   reg __391112_391112;
   reg _391113_391113 ; 
   reg __391113_391113;
   reg _391114_391114 ; 
   reg __391114_391114;
   reg _391115_391115 ; 
   reg __391115_391115;
   reg _391116_391116 ; 
   reg __391116_391116;
   reg _391117_391117 ; 
   reg __391117_391117;
   reg _391118_391118 ; 
   reg __391118_391118;
   reg _391119_391119 ; 
   reg __391119_391119;
   reg _391120_391120 ; 
   reg __391120_391120;
   reg _391121_391121 ; 
   reg __391121_391121;
   reg _391122_391122 ; 
   reg __391122_391122;
   reg _391123_391123 ; 
   reg __391123_391123;
   reg _391124_391124 ; 
   reg __391124_391124;
   reg _391125_391125 ; 
   reg __391125_391125;
   reg _391126_391126 ; 
   reg __391126_391126;
   reg _391127_391127 ; 
   reg __391127_391127;
   reg _391128_391128 ; 
   reg __391128_391128;
   reg _391129_391129 ; 
   reg __391129_391129;
   reg _391130_391130 ; 
   reg __391130_391130;
   reg _391131_391131 ; 
   reg __391131_391131;
   reg _391132_391132 ; 
   reg __391132_391132;
   reg _391133_391133 ; 
   reg __391133_391133;
   reg _391134_391134 ; 
   reg __391134_391134;
   reg _391135_391135 ; 
   reg __391135_391135;
   reg _391136_391136 ; 
   reg __391136_391136;
   reg _391137_391137 ; 
   reg __391137_391137;
   reg _391138_391138 ; 
   reg __391138_391138;
   reg _391139_391139 ; 
   reg __391139_391139;
   reg _391140_391140 ; 
   reg __391140_391140;
   reg _391141_391141 ; 
   reg __391141_391141;
   reg _391142_391142 ; 
   reg __391142_391142;
   reg _391143_391143 ; 
   reg __391143_391143;
   reg _391144_391144 ; 
   reg __391144_391144;
   reg _391145_391145 ; 
   reg __391145_391145;
   reg _391146_391146 ; 
   reg __391146_391146;
   reg _391147_391147 ; 
   reg __391147_391147;
   reg _391148_391148 ; 
   reg __391148_391148;
   reg _391149_391149 ; 
   reg __391149_391149;
   reg _391150_391150 ; 
   reg __391150_391150;
   reg _391151_391151 ; 
   reg __391151_391151;
   reg _391152_391152 ; 
   reg __391152_391152;
   reg _391153_391153 ; 
   reg __391153_391153;
   reg _391154_391154 ; 
   reg __391154_391154;
   reg _391155_391155 ; 
   reg __391155_391155;
   reg _391156_391156 ; 
   reg __391156_391156;
   reg _391157_391157 ; 
   reg __391157_391157;
   reg _391158_391158 ; 
   reg __391158_391158;
   reg _391159_391159 ; 
   reg __391159_391159;
   reg _391160_391160 ; 
   reg __391160_391160;
   reg _391161_391161 ; 
   reg __391161_391161;
   reg _391162_391162 ; 
   reg __391162_391162;
   reg _391163_391163 ; 
   reg __391163_391163;
   reg _391164_391164 ; 
   reg __391164_391164;
   reg _391165_391165 ; 
   reg __391165_391165;
   reg _391166_391166 ; 
   reg __391166_391166;
   reg _391167_391167 ; 
   reg __391167_391167;
   reg _391168_391168 ; 
   reg __391168_391168;
   reg _391169_391169 ; 
   reg __391169_391169;
   reg _391170_391170 ; 
   reg __391170_391170;
   reg _391171_391171 ; 
   reg __391171_391171;
   reg _391172_391172 ; 
   reg __391172_391172;
   reg _391173_391173 ; 
   reg __391173_391173;
   reg _391174_391174 ; 
   reg __391174_391174;
   reg _391175_391175 ; 
   reg __391175_391175;
   reg _391176_391176 ; 
   reg __391176_391176;
   reg _391177_391177 ; 
   reg __391177_391177;
   reg _391178_391178 ; 
   reg __391178_391178;
   reg _391179_391179 ; 
   reg __391179_391179;
   reg _391180_391180 ; 
   reg __391180_391180;
   reg _391181_391181 ; 
   reg __391181_391181;
   reg _391182_391182 ; 
   reg __391182_391182;
   reg _391183_391183 ; 
   reg __391183_391183;
   reg _391184_391184 ; 
   reg __391184_391184;
   reg _391185_391185 ; 
   reg __391185_391185;
   reg _391186_391186 ; 
   reg __391186_391186;
   reg _391187_391187 ; 
   reg __391187_391187;
   reg _391188_391188 ; 
   reg __391188_391188;
   reg _391189_391189 ; 
   reg __391189_391189;
   reg _391190_391190 ; 
   reg __391190_391190;
   reg _391191_391191 ; 
   reg __391191_391191;
   reg _391192_391192 ; 
   reg __391192_391192;
   reg _391193_391193 ; 
   reg __391193_391193;
   reg _391194_391194 ; 
   reg __391194_391194;
   reg _391195_391195 ; 
   reg __391195_391195;
   reg _391196_391196 ; 
   reg __391196_391196;
   reg _391197_391197 ; 
   reg __391197_391197;
   reg _391198_391198 ; 
   reg __391198_391198;
   reg _391199_391199 ; 
   reg __391199_391199;
   reg _391200_391200 ; 
   reg __391200_391200;
   reg _391201_391201 ; 
   reg __391201_391201;
   reg _391202_391202 ; 
   reg __391202_391202;
   reg _391203_391203 ; 
   reg __391203_391203;
   reg _391204_391204 ; 
   reg __391204_391204;
   reg _391205_391205 ; 
   reg __391205_391205;
   reg _391206_391206 ; 
   reg __391206_391206;
   reg _391207_391207 ; 
   reg __391207_391207;
   reg _391208_391208 ; 
   reg __391208_391208;
   reg _391209_391209 ; 
   reg __391209_391209;
   reg _391210_391210 ; 
   reg __391210_391210;
   reg _391211_391211 ; 
   reg __391211_391211;
   reg _391212_391212 ; 
   reg __391212_391212;
   reg _391213_391213 ; 
   reg __391213_391213;
   reg _391214_391214 ; 
   reg __391214_391214;
   reg _391215_391215 ; 
   reg __391215_391215;
   reg _391216_391216 ; 
   reg __391216_391216;
   reg _391217_391217 ; 
   reg __391217_391217;
   reg _391218_391218 ; 
   reg __391218_391218;
   reg _391219_391219 ; 
   reg __391219_391219;
   reg _391220_391220 ; 
   reg __391220_391220;
   reg _391221_391221 ; 
   reg __391221_391221;
   reg _391222_391222 ; 
   reg __391222_391222;
   reg _391223_391223 ; 
   reg __391223_391223;
   reg _391224_391224 ; 
   reg __391224_391224;
   reg _391225_391225 ; 
   reg __391225_391225;
   reg _391226_391226 ; 
   reg __391226_391226;
   reg _391227_391227 ; 
   reg __391227_391227;
   reg _391228_391228 ; 
   reg __391228_391228;
   reg _391229_391229 ; 
   reg __391229_391229;
   reg _391230_391230 ; 
   reg __391230_391230;
   reg _391231_391231 ; 
   reg __391231_391231;
   reg _391232_391232 ; 
   reg __391232_391232;
   reg _391233_391233 ; 
   reg __391233_391233;
   reg _391234_391234 ; 
   reg __391234_391234;
   reg _391235_391235 ; 
   reg __391235_391235;
   reg _391236_391236 ; 
   reg __391236_391236;
   reg _391237_391237 ; 
   reg __391237_391237;
   reg _391238_391238 ; 
   reg __391238_391238;
   reg _391239_391239 ; 
   reg __391239_391239;
   reg _391240_391240 ; 
   reg __391240_391240;
   reg _391241_391241 ; 
   reg __391241_391241;
   reg _391242_391242 ; 
   reg __391242_391242;
   reg _391243_391243 ; 
   reg __391243_391243;
   reg _391244_391244 ; 
   reg __391244_391244;
   reg _391245_391245 ; 
   reg __391245_391245;
   reg _391246_391246 ; 
   reg __391246_391246;
   reg _391247_391247 ; 
   reg __391247_391247;
   reg _391248_391248 ; 
   reg __391248_391248;
   reg _391249_391249 ; 
   reg __391249_391249;
   reg _391250_391250 ; 
   reg __391250_391250;
   reg _391251_391251 ; 
   reg __391251_391251;
   reg _391252_391252 ; 
   reg __391252_391252;
   reg _391253_391253 ; 
   reg __391253_391253;
   reg _391254_391254 ; 
   reg __391254_391254;
   reg _391255_391255 ; 
   reg __391255_391255;
   reg _391256_391256 ; 
   reg __391256_391256;
   reg _391257_391257 ; 
   reg __391257_391257;
   reg _391258_391258 ; 
   reg __391258_391258;
   reg _391259_391259 ; 
   reg __391259_391259;
   reg _391260_391260 ; 
   reg __391260_391260;
   reg _391261_391261 ; 
   reg __391261_391261;
   reg _391262_391262 ; 
   reg __391262_391262;
   reg _391263_391263 ; 
   reg __391263_391263;
   reg _391264_391264 ; 
   reg __391264_391264;
   reg _391265_391265 ; 
   reg __391265_391265;
   reg _391266_391266 ; 
   reg __391266_391266;
   reg _391267_391267 ; 
   reg __391267_391267;
   reg _391268_391268 ; 
   reg __391268_391268;
   reg _391269_391269 ; 
   reg __391269_391269;
   reg _391270_391270 ; 
   reg __391270_391270;
   reg _391271_391271 ; 
   reg __391271_391271;
   reg _391272_391272 ; 
   reg __391272_391272;
   reg _391273_391273 ; 
   reg __391273_391273;
   reg _391274_391274 ; 
   reg __391274_391274;
   reg _391275_391275 ; 
   reg __391275_391275;
   reg _391276_391276 ; 
   reg __391276_391276;
   reg _391277_391277 ; 
   reg __391277_391277;
   reg _391278_391278 ; 
   reg __391278_391278;
   reg _391279_391279 ; 
   reg __391279_391279;
   reg _391280_391280 ; 
   reg __391280_391280;
   reg _391281_391281 ; 
   reg __391281_391281;
   reg _391282_391282 ; 
   reg __391282_391282;
   reg _391283_391283 ; 
   reg __391283_391283;
   reg _391284_391284 ; 
   reg __391284_391284;
   reg _391285_391285 ; 
   reg __391285_391285;
   reg _391286_391286 ; 
   reg __391286_391286;
   reg _391287_391287 ; 
   reg __391287_391287;
   reg _391288_391288 ; 
   reg __391288_391288;
   reg _391289_391289 ; 
   reg __391289_391289;
   reg _391290_391290 ; 
   reg __391290_391290;
   reg _391291_391291 ; 
   reg __391291_391291;
   reg _391292_391292 ; 
   reg __391292_391292;
   reg _391293_391293 ; 
   reg __391293_391293;
   reg _391294_391294 ; 
   reg __391294_391294;
   reg _391295_391295 ; 
   reg __391295_391295;
   reg _391296_391296 ; 
   reg __391296_391296;
   reg _391297_391297 ; 
   reg __391297_391297;
   reg _391298_391298 ; 
   reg __391298_391298;
   reg _391299_391299 ; 
   reg __391299_391299;
   reg _391300_391300 ; 
   reg __391300_391300;
   reg _391301_391301 ; 
   reg __391301_391301;
   reg _391302_391302 ; 
   reg __391302_391302;
   reg _391303_391303 ; 
   reg __391303_391303;
   reg _391304_391304 ; 
   reg __391304_391304;
   reg _391305_391305 ; 
   reg __391305_391305;
   reg _391306_391306 ; 
   reg __391306_391306;
   reg _391307_391307 ; 
   reg __391307_391307;
   reg _391308_391308 ; 
   reg __391308_391308;
   reg _391309_391309 ; 
   reg __391309_391309;
   reg _391310_391310 ; 
   reg __391310_391310;
   reg _391311_391311 ; 
   reg __391311_391311;
   reg _391312_391312 ; 
   reg __391312_391312;
   reg _391313_391313 ; 
   reg __391313_391313;
   reg _391314_391314 ; 
   reg __391314_391314;
   reg _391315_391315 ; 
   reg __391315_391315;
   reg _391316_391316 ; 
   reg __391316_391316;
   reg _391317_391317 ; 
   reg __391317_391317;
   reg _391318_391318 ; 
   reg __391318_391318;
   reg _391319_391319 ; 
   reg __391319_391319;
   reg _391320_391320 ; 
   reg __391320_391320;
   reg _391321_391321 ; 
   reg __391321_391321;
   reg _391322_391322 ; 
   reg __391322_391322;
   reg _391323_391323 ; 
   reg __391323_391323;
   reg _391324_391324 ; 
   reg __391324_391324;
   reg _391325_391325 ; 
   reg __391325_391325;
   reg _391326_391326 ; 
   reg __391326_391326;
   reg _391327_391327 ; 
   reg __391327_391327;
   reg _391328_391328 ; 
   reg __391328_391328;
   reg _391329_391329 ; 
   reg __391329_391329;
   reg _391330_391330 ; 
   reg __391330_391330;
   reg _391331_391331 ; 
   reg __391331_391331;
   reg _391332_391332 ; 
   reg __391332_391332;
   reg _391333_391333 ; 
   reg __391333_391333;
   reg _391334_391334 ; 
   reg __391334_391334;
   reg _391335_391335 ; 
   reg __391335_391335;
   reg _391336_391336 ; 
   reg __391336_391336;
   reg _391337_391337 ; 
   reg __391337_391337;
   reg _391338_391338 ; 
   reg __391338_391338;
   reg _391339_391339 ; 
   reg __391339_391339;
   reg _391340_391340 ; 
   reg __391340_391340;
   reg _391341_391341 ; 
   reg __391341_391341;
   reg _391342_391342 ; 
   reg __391342_391342;
   reg _391343_391343 ; 
   reg __391343_391343;
   reg _391344_391344 ; 
   reg __391344_391344;
   reg _391345_391345 ; 
   reg __391345_391345;
   reg _391346_391346 ; 
   reg __391346_391346;
   reg _391347_391347 ; 
   reg __391347_391347;
   reg _391348_391348 ; 
   reg __391348_391348;
   reg _391349_391349 ; 
   reg __391349_391349;
   reg _391350_391350 ; 
   reg __391350_391350;
   reg _391351_391351 ; 
   reg __391351_391351;
   reg _391352_391352 ; 
   reg __391352_391352;
   reg _391353_391353 ; 
   reg __391353_391353;
   reg _391354_391354 ; 
   reg __391354_391354;
   reg _391355_391355 ; 
   reg __391355_391355;
   reg _391356_391356 ; 
   reg __391356_391356;
   reg _391357_391357 ; 
   reg __391357_391357;
   reg _391358_391358 ; 
   reg __391358_391358;
   reg _391359_391359 ; 
   reg __391359_391359;
   reg _391360_391360 ; 
   reg __391360_391360;
   reg _391361_391361 ; 
   reg __391361_391361;
   reg _391362_391362 ; 
   reg __391362_391362;
   reg _391363_391363 ; 
   reg __391363_391363;
   reg _391364_391364 ; 
   reg __391364_391364;
   reg _391365_391365 ; 
   reg __391365_391365;
   reg _391366_391366 ; 
   reg __391366_391366;
   reg _391367_391367 ; 
   reg __391367_391367;
   reg _391368_391368 ; 
   reg __391368_391368;
   reg _391369_391369 ; 
   reg __391369_391369;
   reg _391370_391370 ; 
   reg __391370_391370;
   reg _391371_391371 ; 
   reg __391371_391371;
   reg _391372_391372 ; 
   reg __391372_391372;
   reg _391373_391373 ; 
   reg __391373_391373;
   reg _391374_391374 ; 
   reg __391374_391374;
   reg _391375_391375 ; 
   reg __391375_391375;
   reg _391376_391376 ; 
   reg __391376_391376;
   reg _391377_391377 ; 
   reg __391377_391377;
   reg _391378_391378 ; 
   reg __391378_391378;
   reg _391379_391379 ; 
   reg __391379_391379;
   reg _391380_391380 ; 
   reg __391380_391380;
   reg _391381_391381 ; 
   reg __391381_391381;
   reg _391382_391382 ; 
   reg __391382_391382;
   reg _391383_391383 ; 
   reg __391383_391383;
   reg _391384_391384 ; 
   reg __391384_391384;
   reg _391385_391385 ; 
   reg __391385_391385;
   reg _391386_391386 ; 
   reg __391386_391386;
   reg _391387_391387 ; 
   reg __391387_391387;
   reg _391388_391388 ; 
   reg __391388_391388;
   reg _391389_391389 ; 
   reg __391389_391389;
   reg _391390_391390 ; 
   reg __391390_391390;
   reg _391391_391391 ; 
   reg __391391_391391;
   reg _391392_391392 ; 
   reg __391392_391392;
   reg _391393_391393 ; 
   reg __391393_391393;
   reg _391394_391394 ; 
   reg __391394_391394;
   reg _391395_391395 ; 
   reg __391395_391395;
   reg _391396_391396 ; 
   reg __391396_391396;
   reg _391397_391397 ; 
   reg __391397_391397;
   reg _391398_391398 ; 
   reg __391398_391398;
   reg _391399_391399 ; 
   reg __391399_391399;
   reg _391400_391400 ; 
   reg __391400_391400;
   reg _391401_391401 ; 
   reg __391401_391401;
   reg _391402_391402 ; 
   reg __391402_391402;
   reg _391403_391403 ; 
   reg __391403_391403;
   reg _391404_391404 ; 
   reg __391404_391404;
   reg _391405_391405 ; 
   reg __391405_391405;
   reg _391406_391406 ; 
   reg __391406_391406;
   reg _391407_391407 ; 
   reg __391407_391407;
   reg _391408_391408 ; 
   reg __391408_391408;
   reg _391409_391409 ; 
   reg __391409_391409;
   reg _391410_391410 ; 
   reg __391410_391410;
   reg _391411_391411 ; 
   reg __391411_391411;
   reg _391412_391412 ; 
   reg __391412_391412;
   reg _391413_391413 ; 
   reg __391413_391413;
   reg _391414_391414 ; 
   reg __391414_391414;
   reg _391415_391415 ; 
   reg __391415_391415;
   reg _391416_391416 ; 
   reg __391416_391416;
   reg _391417_391417 ; 
   reg __391417_391417;
   reg _391418_391418 ; 
   reg __391418_391418;
   reg _391419_391419 ; 
   reg __391419_391419;
   reg _391420_391420 ; 
   reg __391420_391420;
   reg _391421_391421 ; 
   reg __391421_391421;
   reg _391422_391422 ; 
   reg __391422_391422;
   reg _391423_391423 ; 
   reg __391423_391423;
   reg _391424_391424 ; 
   reg __391424_391424;
   reg _391425_391425 ; 
   reg __391425_391425;
   reg _391426_391426 ; 
   reg __391426_391426;
   reg _391427_391427 ; 
   reg __391427_391427;
   reg _391428_391428 ; 
   reg __391428_391428;
   reg _391429_391429 ; 
   reg __391429_391429;
   reg _391430_391430 ; 
   reg __391430_391430;
   reg _391431_391431 ; 
   reg __391431_391431;
   reg _391432_391432 ; 
   reg __391432_391432;
   reg _391433_391433 ; 
   reg __391433_391433;
   reg _391434_391434 ; 
   reg __391434_391434;
   reg _391435_391435 ; 
   reg __391435_391435;
   reg _391436_391436 ; 
   reg __391436_391436;
   reg _391437_391437 ; 
   reg __391437_391437;
   reg _391438_391438 ; 
   reg __391438_391438;
   reg _391439_391439 ; 
   reg __391439_391439;
   reg _391440_391440 ; 
   reg __391440_391440;
   reg _391441_391441 ; 
   reg __391441_391441;
   reg _391442_391442 ; 
   reg __391442_391442;
   reg _391443_391443 ; 
   reg __391443_391443;
   reg _391444_391444 ; 
   reg __391444_391444;
   reg _391445_391445 ; 
   reg __391445_391445;
   reg _391446_391446 ; 
   reg __391446_391446;
   reg _391447_391447 ; 
   reg __391447_391447;
   reg _391448_391448 ; 
   reg __391448_391448;
   reg _391449_391449 ; 
   reg __391449_391449;
   reg _391450_391450 ; 
   reg __391450_391450;
   reg _391451_391451 ; 
   reg __391451_391451;
   reg _391452_391452 ; 
   reg __391452_391452;
   reg _391453_391453 ; 
   reg __391453_391453;
   reg _391454_391454 ; 
   reg __391454_391454;
   reg _391455_391455 ; 
   reg __391455_391455;
   reg _391456_391456 ; 
   reg __391456_391456;
   reg _391457_391457 ; 
   reg __391457_391457;
   reg _391458_391458 ; 
   reg __391458_391458;
   reg _391459_391459 ; 
   reg __391459_391459;
   reg _391460_391460 ; 
   reg __391460_391460;
   reg _391461_391461 ; 
   reg __391461_391461;
   reg _391462_391462 ; 
   reg __391462_391462;
   reg _391463_391463 ; 
   reg __391463_391463;
   reg _391464_391464 ; 
   reg __391464_391464;
   reg _391465_391465 ; 
   reg __391465_391465;
   reg _391466_391466 ; 
   reg __391466_391466;
   reg _391467_391467 ; 
   reg __391467_391467;
   reg _391468_391468 ; 
   reg __391468_391468;
   reg _391469_391469 ; 
   reg __391469_391469;
   reg _391470_391470 ; 
   reg __391470_391470;
   reg _391471_391471 ; 
   reg __391471_391471;
   reg _391472_391472 ; 
   reg __391472_391472;
   reg _391473_391473 ; 
   reg __391473_391473;
   reg _391474_391474 ; 
   reg __391474_391474;
   reg _391475_391475 ; 
   reg __391475_391475;
   reg _391476_391476 ; 
   reg __391476_391476;
   reg _391477_391477 ; 
   reg __391477_391477;
   reg _391478_391478 ; 
   reg __391478_391478;
   reg _391479_391479 ; 
   reg __391479_391479;
   reg _391480_391480 ; 
   reg __391480_391480;
   reg _391481_391481 ; 
   reg __391481_391481;
   reg _391482_391482 ; 
   reg __391482_391482;
   reg _391483_391483 ; 
   reg __391483_391483;
   reg _391484_391484 ; 
   reg __391484_391484;
   reg _391485_391485 ; 
   reg __391485_391485;
   reg _391486_391486 ; 
   reg __391486_391486;
   reg _391487_391487 ; 
   reg __391487_391487;
   reg _391488_391488 ; 
   reg __391488_391488;
   reg _391489_391489 ; 
   reg __391489_391489;
   reg _391490_391490 ; 
   reg __391490_391490;
   reg _391491_391491 ; 
   reg __391491_391491;
   reg _391492_391492 ; 
   reg __391492_391492;
   reg _391493_391493 ; 
   reg __391493_391493;
   reg _391494_391494 ; 
   reg __391494_391494;
   reg _391495_391495 ; 
   reg __391495_391495;
   reg _391496_391496 ; 
   reg __391496_391496;
   reg _391497_391497 ; 
   reg __391497_391497;
   reg _391498_391498 ; 
   reg __391498_391498;
   reg _391499_391499 ; 
   reg __391499_391499;
   reg _391500_391500 ; 
   reg __391500_391500;
   reg _391501_391501 ; 
   reg __391501_391501;
   reg _391502_391502 ; 
   reg __391502_391502;
   reg _391503_391503 ; 
   reg __391503_391503;
   reg _391504_391504 ; 
   reg __391504_391504;
   reg _391505_391505 ; 
   reg __391505_391505;
   reg _391506_391506 ; 
   reg __391506_391506;
   reg _391507_391507 ; 
   reg __391507_391507;
   reg _391508_391508 ; 
   reg __391508_391508;
   reg _391509_391509 ; 
   reg __391509_391509;
   reg _391510_391510 ; 
   reg __391510_391510;
   reg _391511_391511 ; 
   reg __391511_391511;
   reg _391512_391512 ; 
   reg __391512_391512;
   reg _391513_391513 ; 
   reg __391513_391513;
   reg _391514_391514 ; 
   reg __391514_391514;
   reg _391515_391515 ; 
   reg __391515_391515;
   reg _391516_391516 ; 
   reg __391516_391516;
   reg _391517_391517 ; 
   reg __391517_391517;
   reg _391518_391518 ; 
   reg __391518_391518;
   reg _391519_391519 ; 
   reg __391519_391519;
   reg _391520_391520 ; 
   reg __391520_391520;
   reg _391521_391521 ; 
   reg __391521_391521;
   reg _391522_391522 ; 
   reg __391522_391522;
   reg _391523_391523 ; 
   reg __391523_391523;
   reg _391524_391524 ; 
   reg __391524_391524;
   reg _391525_391525 ; 
   reg __391525_391525;
   reg _391526_391526 ; 
   reg __391526_391526;
   reg _391527_391527 ; 
   reg __391527_391527;
   reg _391528_391528 ; 
   reg __391528_391528;
   reg _391529_391529 ; 
   reg __391529_391529;
   reg _391530_391530 ; 
   reg __391530_391530;
   reg _391531_391531 ; 
   reg __391531_391531;
   reg _391532_391532 ; 
   reg __391532_391532;
   reg _391533_391533 ; 
   reg __391533_391533;
   reg _391534_391534 ; 
   reg __391534_391534;
   reg _391535_391535 ; 
   reg __391535_391535;
   reg _391536_391536 ; 
   reg __391536_391536;
   reg _391537_391537 ; 
   reg __391537_391537;
   reg _391538_391538 ; 
   reg __391538_391538;
   reg _391539_391539 ; 
   reg __391539_391539;
   reg _391540_391540 ; 
   reg __391540_391540;
   reg _391541_391541 ; 
   reg __391541_391541;
   reg _391542_391542 ; 
   reg __391542_391542;
   reg _391543_391543 ; 
   reg __391543_391543;
   reg _391544_391544 ; 
   reg __391544_391544;
   reg _391545_391545 ; 
   reg __391545_391545;
   reg _391546_391546 ; 
   reg __391546_391546;
   reg _391547_391547 ; 
   reg __391547_391547;
   reg _391548_391548 ; 
   reg __391548_391548;
   reg _391549_391549 ; 
   reg __391549_391549;
   reg _391550_391550 ; 
   reg __391550_391550;
   reg _391551_391551 ; 
   reg __391551_391551;
   reg _391552_391552 ; 
   reg __391552_391552;
   reg _391553_391553 ; 
   reg __391553_391553;
   reg _391554_391554 ; 
   reg __391554_391554;
   reg _391555_391555 ; 
   reg __391555_391555;
   reg _391556_391556 ; 
   reg __391556_391556;
   reg _391557_391557 ; 
   reg __391557_391557;
   reg _391558_391558 ; 
   reg __391558_391558;
   reg _391559_391559 ; 
   reg __391559_391559;
   reg _391560_391560 ; 
   reg __391560_391560;
   reg _391561_391561 ; 
   reg __391561_391561;
   reg _391562_391562 ; 
   reg __391562_391562;
   reg _391563_391563 ; 
   reg __391563_391563;
   reg _391564_391564 ; 
   reg __391564_391564;
   reg _391565_391565 ; 
   reg __391565_391565;
   reg _391566_391566 ; 
   reg __391566_391566;
   reg _391567_391567 ; 
   reg __391567_391567;
   reg _391568_391568 ; 
   reg __391568_391568;
   reg _391569_391569 ; 
   reg __391569_391569;
   reg _391570_391570 ; 
   reg __391570_391570;
   reg _391571_391571 ; 
   reg __391571_391571;
   reg _391572_391572 ; 
   reg __391572_391572;
   reg _391573_391573 ; 
   reg __391573_391573;
   reg _391574_391574 ; 
   reg __391574_391574;
   reg _391575_391575 ; 
   reg __391575_391575;
   reg _391576_391576 ; 
   reg __391576_391576;
   reg _391577_391577 ; 
   reg __391577_391577;
   reg _391578_391578 ; 
   reg __391578_391578;
   reg _391579_391579 ; 
   reg __391579_391579;
   reg _391580_391580 ; 
   reg __391580_391580;
   reg _391581_391581 ; 
   reg __391581_391581;
   reg _391582_391582 ; 
   reg __391582_391582;
   reg _391583_391583 ; 
   reg __391583_391583;
   reg _391584_391584 ; 
   reg __391584_391584;
   reg _391585_391585 ; 
   reg __391585_391585;
   reg _391586_391586 ; 
   reg __391586_391586;
   reg _391587_391587 ; 
   reg __391587_391587;
   reg _391588_391588 ; 
   reg __391588_391588;
   reg _391589_391589 ; 
   reg __391589_391589;
   reg _391590_391590 ; 
   reg __391590_391590;
   reg _391591_391591 ; 
   reg __391591_391591;
   reg _391592_391592 ; 
   reg __391592_391592;
   reg _391593_391593 ; 
   reg __391593_391593;
   reg _391594_391594 ; 
   reg __391594_391594;
   reg _391595_391595 ; 
   reg __391595_391595;
   reg _391596_391596 ; 
   reg __391596_391596;
   reg _391597_391597 ; 
   reg __391597_391597;
   reg _391598_391598 ; 
   reg __391598_391598;
   reg _391599_391599 ; 
   reg __391599_391599;
   reg _391600_391600 ; 
   reg __391600_391600;
   reg _391601_391601 ; 
   reg __391601_391601;
   reg _391602_391602 ; 
   reg __391602_391602;
   reg _391603_391603 ; 
   reg __391603_391603;
   reg _391604_391604 ; 
   reg __391604_391604;
   reg _391605_391605 ; 
   reg __391605_391605;
   reg _391606_391606 ; 
   reg __391606_391606;
   reg _391607_391607 ; 
   reg __391607_391607;
   reg _391608_391608 ; 
   reg __391608_391608;
   reg _391609_391609 ; 
   reg __391609_391609;
   reg _391610_391610 ; 
   reg __391610_391610;
   reg _391611_391611 ; 
   reg __391611_391611;
   reg _391612_391612 ; 
   reg __391612_391612;
   reg _391613_391613 ; 
   reg __391613_391613;
   reg _391614_391614 ; 
   reg __391614_391614;
   reg _391615_391615 ; 
   reg __391615_391615;
   reg _391616_391616 ; 
   reg __391616_391616;
   reg _391617_391617 ; 
   reg __391617_391617;
   reg _391618_391618 ; 
   reg __391618_391618;
   reg _391619_391619 ; 
   reg __391619_391619;
   reg _391620_391620 ; 
   reg __391620_391620;
   reg _391621_391621 ; 
   reg __391621_391621;
   reg _391622_391622 ; 
   reg __391622_391622;
   reg _391623_391623 ; 
   reg __391623_391623;
   reg _391624_391624 ; 
   reg __391624_391624;
   reg _391625_391625 ; 
   reg __391625_391625;
   reg _391626_391626 ; 
   reg __391626_391626;
   reg _391627_391627 ; 
   reg __391627_391627;
   reg _391628_391628 ; 
   reg __391628_391628;
   reg _391629_391629 ; 
   reg __391629_391629;
   reg _391630_391630 ; 
   reg __391630_391630;
   reg _391631_391631 ; 
   reg __391631_391631;
   reg _391632_391632 ; 
   reg __391632_391632;
   reg _391633_391633 ; 
   reg __391633_391633;
   reg _391634_391634 ; 
   reg __391634_391634;
   reg _391635_391635 ; 
   reg __391635_391635;
   reg _391636_391636 ; 
   reg __391636_391636;
   reg _391637_391637 ; 
   reg __391637_391637;
   reg _391638_391638 ; 
   reg __391638_391638;
   reg _391639_391639 ; 
   reg __391639_391639;
   reg _391640_391640 ; 
   reg __391640_391640;
   reg _391641_391641 ; 
   reg __391641_391641;
   reg _391642_391642 ; 
   reg __391642_391642;
   reg _391643_391643 ; 
   reg __391643_391643;
   reg _391644_391644 ; 
   reg __391644_391644;
   reg _391645_391645 ; 
   reg __391645_391645;
   reg _391646_391646 ; 
   reg __391646_391646;
   reg _391647_391647 ; 
   reg __391647_391647;
   reg _391648_391648 ; 
   reg __391648_391648;
   reg _391649_391649 ; 
   reg __391649_391649;
   reg _391650_391650 ; 
   reg __391650_391650;
   reg _391651_391651 ; 
   reg __391651_391651;
   reg _391652_391652 ; 
   reg __391652_391652;
   reg _391653_391653 ; 
   reg __391653_391653;
   reg _391654_391654 ; 
   reg __391654_391654;
   reg _391655_391655 ; 
   reg __391655_391655;
   reg _391656_391656 ; 
   reg __391656_391656;
   reg _391657_391657 ; 
   reg __391657_391657;
   reg _391658_391658 ; 
   reg __391658_391658;
   reg _391659_391659 ; 
   reg __391659_391659;
   reg _391660_391660 ; 
   reg __391660_391660;
   reg _391661_391661 ; 
   reg __391661_391661;
   reg _391662_391662 ; 
   reg __391662_391662;
   reg _391663_391663 ; 
   reg __391663_391663;
   reg _391664_391664 ; 
   reg __391664_391664;
   reg _391665_391665 ; 
   reg __391665_391665;
   reg _391666_391666 ; 
   reg __391666_391666;
   reg _391667_391667 ; 
   reg __391667_391667;
   reg _391668_391668 ; 
   reg __391668_391668;
   reg _391669_391669 ; 
   reg __391669_391669;
   reg _391670_391670 ; 
   reg __391670_391670;
   reg _391671_391671 ; 
   reg __391671_391671;
   reg _391672_391672 ; 
   reg __391672_391672;
   reg _391673_391673 ; 
   reg __391673_391673;
   reg _391674_391674 ; 
   reg __391674_391674;
   reg _391675_391675 ; 
   reg __391675_391675;
   reg _391676_391676 ; 
   reg __391676_391676;
   reg _391677_391677 ; 
   reg __391677_391677;
   reg _391678_391678 ; 
   reg __391678_391678;
   reg _391679_391679 ; 
   reg __391679_391679;
   reg _391680_391680 ; 
   reg __391680_391680;
   reg _391681_391681 ; 
   reg __391681_391681;
   reg _391682_391682 ; 
   reg __391682_391682;
   reg _391683_391683 ; 
   reg __391683_391683;
   reg _391684_391684 ; 
   reg __391684_391684;
   reg _391685_391685 ; 
   reg __391685_391685;
   reg _391686_391686 ; 
   reg __391686_391686;
   reg _391687_391687 ; 
   reg __391687_391687;
   reg _391688_391688 ; 
   reg __391688_391688;
   reg _391689_391689 ; 
   reg __391689_391689;
   reg _391690_391690 ; 
   reg __391690_391690;
   reg _391691_391691 ; 
   reg __391691_391691;
   reg _391692_391692 ; 
   reg __391692_391692;
   reg _391693_391693 ; 
   reg __391693_391693;
   reg _391694_391694 ; 
   reg __391694_391694;
   reg _391695_391695 ; 
   reg __391695_391695;
   reg _391696_391696 ; 
   reg __391696_391696;
   reg _391697_391697 ; 
   reg __391697_391697;
   reg _391698_391698 ; 
   reg __391698_391698;
   reg _391699_391699 ; 
   reg __391699_391699;
   reg _391700_391700 ; 
   reg __391700_391700;
   reg _391701_391701 ; 
   reg __391701_391701;
   reg _391702_391702 ; 
   reg __391702_391702;
   reg _391703_391703 ; 
   reg __391703_391703;
   reg _391704_391704 ; 
   reg __391704_391704;
   reg _391705_391705 ; 
   reg __391705_391705;
   reg _391706_391706 ; 
   reg __391706_391706;
   reg _391707_391707 ; 
   reg __391707_391707;
   reg _391708_391708 ; 
   reg __391708_391708;
   reg _391709_391709 ; 
   reg __391709_391709;
   reg _391710_391710 ; 
   reg __391710_391710;
   reg _391711_391711 ; 
   reg __391711_391711;
   reg _391712_391712 ; 
   reg __391712_391712;
   reg _391713_391713 ; 
   reg __391713_391713;
   reg _391714_391714 ; 
   reg __391714_391714;
   reg _391715_391715 ; 
   reg __391715_391715;
   reg _391716_391716 ; 
   reg __391716_391716;
   reg _391717_391717 ; 
   reg __391717_391717;
   reg _391718_391718 ; 
   reg __391718_391718;
   reg _391719_391719 ; 
   reg __391719_391719;
   reg _391720_391720 ; 
   reg __391720_391720;
   reg _391721_391721 ; 
   reg __391721_391721;
   reg _391722_391722 ; 
   reg __391722_391722;
   reg _391723_391723 ; 
   reg __391723_391723;
   reg _391724_391724 ; 
   reg __391724_391724;
   reg _391725_391725 ; 
   reg __391725_391725;
   reg _391726_391726 ; 
   reg __391726_391726;
   reg _391727_391727 ; 
   reg __391727_391727;
   reg _391728_391728 ; 
   reg __391728_391728;
   reg _391729_391729 ; 
   reg __391729_391729;
   reg _391730_391730 ; 
   reg __391730_391730;
   reg _391731_391731 ; 
   reg __391731_391731;
   reg _391732_391732 ; 
   reg __391732_391732;
   reg _391733_391733 ; 
   reg __391733_391733;
   reg _391734_391734 ; 
   reg __391734_391734;
   reg _391735_391735 ; 
   reg __391735_391735;
   reg _391736_391736 ; 
   reg __391736_391736;
   reg _391737_391737 ; 
   reg __391737_391737;
   reg _391738_391738 ; 
   reg __391738_391738;
   reg _391739_391739 ; 
   reg __391739_391739;
   reg _391740_391740 ; 
   reg __391740_391740;
   reg _391741_391741 ; 
   reg __391741_391741;
   reg _391742_391742 ; 
   reg __391742_391742;
   reg _391743_391743 ; 
   reg __391743_391743;
   reg _391744_391744 ; 
   reg __391744_391744;
   reg _391745_391745 ; 
   reg __391745_391745;
   reg _391746_391746 ; 
   reg __391746_391746;
   reg _391747_391747 ; 
   reg __391747_391747;
   reg _391748_391748 ; 
   reg __391748_391748;
   reg _391749_391749 ; 
   reg __391749_391749;
   reg _391750_391750 ; 
   reg __391750_391750;
   reg _391751_391751 ; 
   reg __391751_391751;
   reg _391752_391752 ; 
   reg __391752_391752;
   reg _391753_391753 ; 
   reg __391753_391753;
   reg _391754_391754 ; 
   reg __391754_391754;
   reg _391755_391755 ; 
   reg __391755_391755;
   reg _391756_391756 ; 
   reg __391756_391756;
   reg _391757_391757 ; 
   reg __391757_391757;
   reg _391758_391758 ; 
   reg __391758_391758;
   reg _391759_391759 ; 
   reg __391759_391759;
   reg _391760_391760 ; 
   reg __391760_391760;
   reg _391761_391761 ; 
   reg __391761_391761;
   reg _391762_391762 ; 
   reg __391762_391762;
   reg _391763_391763 ; 
   reg __391763_391763;
   reg _391764_391764 ; 
   reg __391764_391764;
   reg _391765_391765 ; 
   reg __391765_391765;
   reg _391766_391766 ; 
   reg __391766_391766;
   reg _391767_391767 ; 
   reg __391767_391767;
   reg _391768_391768 ; 
   reg __391768_391768;
   reg _391769_391769 ; 
   reg __391769_391769;
   reg _391770_391770 ; 
   reg __391770_391770;
   reg _391771_391771 ; 
   reg __391771_391771;
   reg _391772_391772 ; 
   reg __391772_391772;
   reg _391773_391773 ; 
   reg __391773_391773;
   reg _391774_391774 ; 
   reg __391774_391774;
   reg _391775_391775 ; 
   reg __391775_391775;
   reg _391776_391776 ; 
   reg __391776_391776;
   reg _391777_391777 ; 
   reg __391777_391777;
   reg _391778_391778 ; 
   reg __391778_391778;
   reg _391779_391779 ; 
   reg __391779_391779;
   reg _391780_391780 ; 
   reg __391780_391780;
   reg _391781_391781 ; 
   reg __391781_391781;
   reg _391782_391782 ; 
   reg __391782_391782;
   reg _391783_391783 ; 
   reg __391783_391783;
   reg _391784_391784 ; 
   reg __391784_391784;
   reg _391785_391785 ; 
   reg __391785_391785;
   reg _391786_391786 ; 
   reg __391786_391786;
   reg _391787_391787 ; 
   reg __391787_391787;
   reg _391788_391788 ; 
   reg __391788_391788;
   reg _391789_391789 ; 
   reg __391789_391789;
   reg _391790_391790 ; 
   reg __391790_391790;
   reg _391791_391791 ; 
   reg __391791_391791;
   reg _391792_391792 ; 
   reg __391792_391792;
   reg _391793_391793 ; 
   reg __391793_391793;
   reg _391794_391794 ; 
   reg __391794_391794;
   reg _391795_391795 ; 
   reg __391795_391795;
   reg _391796_391796 ; 
   reg __391796_391796;
   reg _391797_391797 ; 
   reg __391797_391797;
   reg _391798_391798 ; 
   reg __391798_391798;
   reg _391799_391799 ; 
   reg __391799_391799;
   reg _391800_391800 ; 
   reg __391800_391800;
   reg _391801_391801 ; 
   reg __391801_391801;
   reg _391802_391802 ; 
   reg __391802_391802;
   reg _391803_391803 ; 
   reg __391803_391803;
   reg _391804_391804 ; 
   reg __391804_391804;
   reg _391805_391805 ; 
   reg __391805_391805;
   reg _391806_391806 ; 
   reg __391806_391806;
   reg _391807_391807 ; 
   reg __391807_391807;
   reg _391808_391808 ; 
   reg __391808_391808;
   reg _391809_391809 ; 
   reg __391809_391809;
   reg _391810_391810 ; 
   reg __391810_391810;
   reg _391811_391811 ; 
   reg __391811_391811;
   reg _391812_391812 ; 
   reg __391812_391812;
   reg _391813_391813 ; 
   reg __391813_391813;
   reg _391814_391814 ; 
   reg __391814_391814;
   reg _391815_391815 ; 
   reg __391815_391815;
   reg _391816_391816 ; 
   reg __391816_391816;
   reg _391817_391817 ; 
   reg __391817_391817;
   reg _391818_391818 ; 
   reg __391818_391818;
   reg _391819_391819 ; 
   reg __391819_391819;
   reg _391820_391820 ; 
   reg __391820_391820;
   reg _391821_391821 ; 
   reg __391821_391821;
   reg _391822_391822 ; 
   reg __391822_391822;
   reg _391823_391823 ; 
   reg __391823_391823;
   reg _391824_391824 ; 
   reg __391824_391824;
   reg _391825_391825 ; 
   reg __391825_391825;
   reg _391826_391826 ; 
   reg __391826_391826;
   reg _391827_391827 ; 
   reg __391827_391827;
   reg _391828_391828 ; 
   reg __391828_391828;
   reg _391829_391829 ; 
   reg __391829_391829;
   reg _391830_391830 ; 
   reg __391830_391830;
   reg _391831_391831 ; 
   reg __391831_391831;
   reg _391832_391832 ; 
   reg __391832_391832;
   reg _391833_391833 ; 
   reg __391833_391833;
   reg _391834_391834 ; 
   reg __391834_391834;
   reg _391835_391835 ; 
   reg __391835_391835;
   reg _391836_391836 ; 
   reg __391836_391836;
   reg _391837_391837 ; 
   reg __391837_391837;
   reg _391838_391838 ; 
   reg __391838_391838;
   reg _391839_391839 ; 
   reg __391839_391839;
   reg _391840_391840 ; 
   reg __391840_391840;
   reg _391841_391841 ; 
   reg __391841_391841;
   reg _391842_391842 ; 
   reg __391842_391842;
   reg _391843_391843 ; 
   reg __391843_391843;
   reg _391844_391844 ; 
   reg __391844_391844;
   reg _391845_391845 ; 
   reg __391845_391845;
   reg _391846_391846 ; 
   reg __391846_391846;
   reg _391847_391847 ; 
   reg __391847_391847;
   reg _391848_391848 ; 
   reg __391848_391848;
   reg _391849_391849 ; 
   reg __391849_391849;
   reg _391850_391850 ; 
   reg __391850_391850;
   reg _391851_391851 ; 
   reg __391851_391851;
   reg _391852_391852 ; 
   reg __391852_391852;
   reg _391853_391853 ; 
   reg __391853_391853;
   reg _391854_391854 ; 
   reg __391854_391854;
   reg _391855_391855 ; 
   reg __391855_391855;
   reg _391856_391856 ; 
   reg __391856_391856;
   reg _391857_391857 ; 
   reg __391857_391857;
   reg _391858_391858 ; 
   reg __391858_391858;
   reg _391859_391859 ; 
   reg __391859_391859;
   reg _391860_391860 ; 
   reg __391860_391860;
   reg _391861_391861 ; 
   reg __391861_391861;
   reg _391862_391862 ; 
   reg __391862_391862;
   reg _391863_391863 ; 
   reg __391863_391863;
   reg _391864_391864 ; 
   reg __391864_391864;
   reg _391865_391865 ; 
   reg __391865_391865;
   reg _391866_391866 ; 
   reg __391866_391866;
   reg _391867_391867 ; 
   reg __391867_391867;
   reg _391868_391868 ; 
   reg __391868_391868;
   reg _391869_391869 ; 
   reg __391869_391869;
   reg _391870_391870 ; 
   reg __391870_391870;
   reg _391871_391871 ; 
   reg __391871_391871;
   reg _391872_391872 ; 
   reg __391872_391872;
   reg _391873_391873 ; 
   reg __391873_391873;
   reg _391874_391874 ; 
   reg __391874_391874;
   reg _391875_391875 ; 
   reg __391875_391875;
   reg _391876_391876 ; 
   reg __391876_391876;
   reg _391877_391877 ; 
   reg __391877_391877;
   reg _391878_391878 ; 
   reg __391878_391878;
   reg _391879_391879 ; 
   reg __391879_391879;
   reg _391880_391880 ; 
   reg __391880_391880;
   reg _391881_391881 ; 
   reg __391881_391881;
   reg _391882_391882 ; 
   reg __391882_391882;
   reg _391883_391883 ; 
   reg __391883_391883;
   reg _391884_391884 ; 
   reg __391884_391884;
   reg _391885_391885 ; 
   reg __391885_391885;
   reg _391886_391886 ; 
   reg __391886_391886;
   reg _391887_391887 ; 
   reg __391887_391887;
   reg _391888_391888 ; 
   reg __391888_391888;
   reg _391889_391889 ; 
   reg __391889_391889;
   reg _391890_391890 ; 
   reg __391890_391890;
   reg _391891_391891 ; 
   reg __391891_391891;
   reg _391892_391892 ; 
   reg __391892_391892;
   reg _391893_391893 ; 
   reg __391893_391893;
   reg _391894_391894 ; 
   reg __391894_391894;
   reg _391895_391895 ; 
   reg __391895_391895;
   reg _391896_391896 ; 
   reg __391896_391896;
   reg _391897_391897 ; 
   reg __391897_391897;
   reg _391898_391898 ; 
   reg __391898_391898;
   reg _391899_391899 ; 
   reg __391899_391899;
   reg _391900_391900 ; 
   reg __391900_391900;
   reg _391901_391901 ; 
   reg __391901_391901;
   reg _391902_391902 ; 
   reg __391902_391902;
   reg _391903_391903 ; 
   reg __391903_391903;
   reg _391904_391904 ; 
   reg __391904_391904;
   reg _391905_391905 ; 
   reg __391905_391905;
   reg _391906_391906 ; 
   reg __391906_391906;
   reg _391907_391907 ; 
   reg __391907_391907;
   reg _391908_391908 ; 
   reg __391908_391908;
   reg _391909_391909 ; 
   reg __391909_391909;
   reg _391910_391910 ; 
   reg __391910_391910;
   reg _391911_391911 ; 
   reg __391911_391911;
   reg _391912_391912 ; 
   reg __391912_391912;
   reg _391913_391913 ; 
   reg __391913_391913;
   reg _391914_391914 ; 
   reg __391914_391914;
   reg _391915_391915 ; 
   reg __391915_391915;
   reg _391916_391916 ; 
   reg __391916_391916;
   reg _391917_391917 ; 
   reg __391917_391917;
   reg _391918_391918 ; 
   reg __391918_391918;
   reg _391919_391919 ; 
   reg __391919_391919;
   reg _391920_391920 ; 
   reg __391920_391920;
   reg _391921_391921 ; 
   reg __391921_391921;
   reg _391922_391922 ; 
   reg __391922_391922;
   reg _391923_391923 ; 
   reg __391923_391923;
   reg _391924_391924 ; 
   reg __391924_391924;
   reg _391925_391925 ; 
   reg __391925_391925;
   reg _391926_391926 ; 
   reg __391926_391926;
   reg _391927_391927 ; 
   reg __391927_391927;
   reg _391928_391928 ; 
   reg __391928_391928;
   reg _391929_391929 ; 
   reg __391929_391929;
   reg _391930_391930 ; 
   reg __391930_391930;
   reg _391931_391931 ; 
   reg __391931_391931;
   reg _391932_391932 ; 
   reg __391932_391932;
   reg _391933_391933 ; 
   reg __391933_391933;
   reg _391934_391934 ; 
   reg __391934_391934;
   reg _391935_391935 ; 
   reg __391935_391935;
   reg _391936_391936 ; 
   reg __391936_391936;
   reg _391937_391937 ; 
   reg __391937_391937;
   reg _391938_391938 ; 
   reg __391938_391938;
   reg _391939_391939 ; 
   reg __391939_391939;
   reg _391940_391940 ; 
   reg __391940_391940;
   reg _391941_391941 ; 
   reg __391941_391941;
   reg _391942_391942 ; 
   reg __391942_391942;
   reg _391943_391943 ; 
   reg __391943_391943;
   reg _391944_391944 ; 
   reg __391944_391944;
   reg _391945_391945 ; 
   reg __391945_391945;
   reg _391946_391946 ; 
   reg __391946_391946;
   reg _391947_391947 ; 
   reg __391947_391947;
   reg _391948_391948 ; 
   reg __391948_391948;
   reg _391949_391949 ; 
   reg __391949_391949;
   reg _391950_391950 ; 
   reg __391950_391950;
   reg _391951_391951 ; 
   reg __391951_391951;
   reg _391952_391952 ; 
   reg __391952_391952;
   reg _391953_391953 ; 
   reg __391953_391953;
   reg _391954_391954 ; 
   reg __391954_391954;
   reg _391955_391955 ; 
   reg __391955_391955;
   reg _391956_391956 ; 
   reg __391956_391956;
   reg _391957_391957 ; 
   reg __391957_391957;
   reg _391958_391958 ; 
   reg __391958_391958;
   reg _391959_391959 ; 
   reg __391959_391959;
   reg _391960_391960 ; 
   reg __391960_391960;
   reg _391961_391961 ; 
   reg __391961_391961;
   reg _391962_391962 ; 
   reg __391962_391962;
   reg _391963_391963 ; 
   reg __391963_391963;
   reg _391964_391964 ; 
   reg __391964_391964;
   reg _391965_391965 ; 
   reg __391965_391965;
   reg _391966_391966 ; 
   reg __391966_391966;
   reg _391967_391967 ; 
   reg __391967_391967;
   reg _391968_391968 ; 
   reg __391968_391968;
   reg _391969_391969 ; 
   reg __391969_391969;
   reg _391970_391970 ; 
   reg __391970_391970;
   reg _391971_391971 ; 
   reg __391971_391971;
   reg _391972_391972 ; 
   reg __391972_391972;
   reg _391973_391973 ; 
   reg __391973_391973;
   reg _391974_391974 ; 
   reg __391974_391974;
   reg _391975_391975 ; 
   reg __391975_391975;
   reg _391976_391976 ; 
   reg __391976_391976;
   reg _391977_391977 ; 
   reg __391977_391977;
   reg _391978_391978 ; 
   reg __391978_391978;
   reg _391979_391979 ; 
   reg __391979_391979;
   reg _391980_391980 ; 
   reg __391980_391980;
   reg _391981_391981 ; 
   reg __391981_391981;
   reg _391982_391982 ; 
   reg __391982_391982;
   reg _391983_391983 ; 
   reg __391983_391983;
   reg _391984_391984 ; 
   reg __391984_391984;
   reg _391985_391985 ; 
   reg __391985_391985;
   reg _391986_391986 ; 
   reg __391986_391986;
   reg _391987_391987 ; 
   reg __391987_391987;
   reg _391988_391988 ; 
   reg __391988_391988;
   reg _391989_391989 ; 
   reg __391989_391989;
   reg _391990_391990 ; 
   reg __391990_391990;
   reg _391991_391991 ; 
   reg __391991_391991;
   reg _391992_391992 ; 
   reg __391992_391992;
   reg _391993_391993 ; 
   reg __391993_391993;
   reg _391994_391994 ; 
   reg __391994_391994;
   reg _391995_391995 ; 
   reg __391995_391995;
   reg _391996_391996 ; 
   reg __391996_391996;
   reg _391997_391997 ; 
   reg __391997_391997;
   reg _391998_391998 ; 
   reg __391998_391998;
   reg _391999_391999 ; 
   reg __391999_391999;
   reg _392000_392000 ; 
   reg __392000_392000;
   reg _392001_392001 ; 
   reg __392001_392001;
   reg _392002_392002 ; 
   reg __392002_392002;
   reg _392003_392003 ; 
   reg __392003_392003;
   reg _392004_392004 ; 
   reg __392004_392004;
   reg _392005_392005 ; 
   reg __392005_392005;
   reg _392006_392006 ; 
   reg __392006_392006;
   reg _392007_392007 ; 
   reg __392007_392007;
   reg _392008_392008 ; 
   reg __392008_392008;
   reg _392009_392009 ; 
   reg __392009_392009;
   reg _392010_392010 ; 
   reg __392010_392010;
   reg _392011_392011 ; 
   reg __392011_392011;
   reg _392012_392012 ; 
   reg __392012_392012;
   reg _392013_392013 ; 
   reg __392013_392013;
   reg _392014_392014 ; 
   reg __392014_392014;
   reg _392015_392015 ; 
   reg __392015_392015;
   reg _392016_392016 ; 
   reg __392016_392016;
   reg _392017_392017 ; 
   reg __392017_392017;
   reg _392018_392018 ; 
   reg __392018_392018;
   reg _392019_392019 ; 
   reg __392019_392019;
   reg _392020_392020 ; 
   reg __392020_392020;
   reg _392021_392021 ; 
   reg __392021_392021;
   reg _392022_392022 ; 
   reg __392022_392022;
   reg _392023_392023 ; 
   reg __392023_392023;
   reg _392024_392024 ; 
   reg __392024_392024;
   reg _392025_392025 ; 
   reg __392025_392025;
   reg _392026_392026 ; 
   reg __392026_392026;
   reg _392027_392027 ; 
   reg __392027_392027;
   reg _392028_392028 ; 
   reg __392028_392028;
   reg _392029_392029 ; 
   reg __392029_392029;
   reg _392030_392030 ; 
   reg __392030_392030;
   reg _392031_392031 ; 
   reg __392031_392031;
   reg _392032_392032 ; 
   reg __392032_392032;
   reg _392033_392033 ; 
   reg __392033_392033;
   reg _392034_392034 ; 
   reg __392034_392034;
   reg _392035_392035 ; 
   reg __392035_392035;
   reg _392036_392036 ; 
   reg __392036_392036;
   reg _392037_392037 ; 
   reg __392037_392037;
   reg _392038_392038 ; 
   reg __392038_392038;
   reg _392039_392039 ; 
   reg __392039_392039;
   reg _392040_392040 ; 
   reg __392040_392040;
   reg _392041_392041 ; 
   reg __392041_392041;
   reg _392042_392042 ; 
   reg __392042_392042;
   reg _392043_392043 ; 
   reg __392043_392043;
   reg _392044_392044 ; 
   reg __392044_392044;
   reg _392045_392045 ; 
   reg __392045_392045;
   reg _392046_392046 ; 
   reg __392046_392046;
   reg _392047_392047 ; 
   reg __392047_392047;
   reg _392048_392048 ; 
   reg __392048_392048;
   reg _392049_392049 ; 
   reg __392049_392049;
   reg _392050_392050 ; 
   reg __392050_392050;
   reg _392051_392051 ; 
   reg __392051_392051;
   reg _392052_392052 ; 
   reg __392052_392052;
   reg _392053_392053 ; 
   reg __392053_392053;
   reg _392054_392054 ; 
   reg __392054_392054;
   reg _392055_392055 ; 
   reg __392055_392055;
   reg _392056_392056 ; 
   reg __392056_392056;
   reg _392057_392057 ; 
   reg __392057_392057;
   reg _392058_392058 ; 
   reg __392058_392058;
   reg _392059_392059 ; 
   reg __392059_392059;
   reg _392060_392060 ; 
   reg __392060_392060;
   reg _392061_392061 ; 
   reg __392061_392061;
   reg _392062_392062 ; 
   reg __392062_392062;
   reg _392063_392063 ; 
   reg __392063_392063;
   reg _392064_392064 ; 
   reg __392064_392064;
   reg _392065_392065 ; 
   reg __392065_392065;
   reg _392066_392066 ; 
   reg __392066_392066;
   reg _392067_392067 ; 
   reg __392067_392067;
   reg _392068_392068 ; 
   reg __392068_392068;
   reg _392069_392069 ; 
   reg __392069_392069;
   reg _392070_392070 ; 
   reg __392070_392070;
   reg _392071_392071 ; 
   reg __392071_392071;
   reg _392072_392072 ; 
   reg __392072_392072;
   reg _392073_392073 ; 
   reg __392073_392073;
   reg _392074_392074 ; 
   reg __392074_392074;
   reg _392075_392075 ; 
   reg __392075_392075;
   reg _392076_392076 ; 
   reg __392076_392076;
   reg _392077_392077 ; 
   reg __392077_392077;
   reg _392078_392078 ; 
   reg __392078_392078;
   reg _392079_392079 ; 
   reg __392079_392079;
   reg _392080_392080 ; 
   reg __392080_392080;
   reg _392081_392081 ; 
   reg __392081_392081;
   reg _392082_392082 ; 
   reg __392082_392082;
   reg _392083_392083 ; 
   reg __392083_392083;
   reg _392084_392084 ; 
   reg __392084_392084;
   reg _392085_392085 ; 
   reg __392085_392085;
   reg _392086_392086 ; 
   reg __392086_392086;
   reg _392087_392087 ; 
   reg __392087_392087;
   reg _392088_392088 ; 
   reg __392088_392088;
   reg _392089_392089 ; 
   reg __392089_392089;
   reg _392090_392090 ; 
   reg __392090_392090;
   reg _392091_392091 ; 
   reg __392091_392091;
   reg _392092_392092 ; 
   reg __392092_392092;
   reg _392093_392093 ; 
   reg __392093_392093;
   reg _392094_392094 ; 
   reg __392094_392094;
   reg _392095_392095 ; 
   reg __392095_392095;
   reg _392096_392096 ; 
   reg __392096_392096;
   reg _392097_392097 ; 
   reg __392097_392097;
   reg _392098_392098 ; 
   reg __392098_392098;
   reg _392099_392099 ; 
   reg __392099_392099;
   reg _392100_392100 ; 
   reg __392100_392100;
   reg _392101_392101 ; 
   reg __392101_392101;
   reg _392102_392102 ; 
   reg __392102_392102;
   reg _392103_392103 ; 
   reg __392103_392103;
   reg _392104_392104 ; 
   reg __392104_392104;
   reg _392105_392105 ; 
   reg __392105_392105;
   reg _392106_392106 ; 
   reg __392106_392106;
   reg _392107_392107 ; 
   reg __392107_392107;
   reg _392108_392108 ; 
   reg __392108_392108;
   reg _392109_392109 ; 
   reg __392109_392109;
   reg _392110_392110 ; 
   reg __392110_392110;
   reg _392111_392111 ; 
   reg __392111_392111;
   reg _392112_392112 ; 
   reg __392112_392112;
   reg _392113_392113 ; 
   reg __392113_392113;
   reg _392114_392114 ; 
   reg __392114_392114;
   reg _392115_392115 ; 
   reg __392115_392115;
   reg _392116_392116 ; 
   reg __392116_392116;
   reg _392117_392117 ; 
   reg __392117_392117;
   reg _392118_392118 ; 
   reg __392118_392118;
   reg _392119_392119 ; 
   reg __392119_392119;
   reg _392120_392120 ; 
   reg __392120_392120;
   reg _392121_392121 ; 
   reg __392121_392121;
   reg _392122_392122 ; 
   reg __392122_392122;
   reg _392123_392123 ; 
   reg __392123_392123;
   reg _392124_392124 ; 
   reg __392124_392124;
   reg _392125_392125 ; 
   reg __392125_392125;
   reg _392126_392126 ; 
   reg __392126_392126;
   reg _392127_392127 ; 
   reg __392127_392127;
   reg _392128_392128 ; 
   reg __392128_392128;
   reg _392129_392129 ; 
   reg __392129_392129;
   reg _392130_392130 ; 
   reg __392130_392130;
   reg _392131_392131 ; 
   reg __392131_392131;
   reg _392132_392132 ; 
   reg __392132_392132;
   reg _392133_392133 ; 
   reg __392133_392133;
   reg _392134_392134 ; 
   reg __392134_392134;
   reg _392135_392135 ; 
   reg __392135_392135;
   reg _392136_392136 ; 
   reg __392136_392136;
   reg _392137_392137 ; 
   reg __392137_392137;
   reg _392138_392138 ; 
   reg __392138_392138;
   reg _392139_392139 ; 
   reg __392139_392139;
   reg _392140_392140 ; 
   reg __392140_392140;
   reg _392141_392141 ; 
   reg __392141_392141;
   reg _392142_392142 ; 
   reg __392142_392142;
   reg _392143_392143 ; 
   reg __392143_392143;
   reg _392144_392144 ; 
   reg __392144_392144;
   reg _392145_392145 ; 
   reg __392145_392145;
   reg _392146_392146 ; 
   reg __392146_392146;
   reg _392147_392147 ; 
   reg __392147_392147;
   reg _392148_392148 ; 
   reg __392148_392148;
   reg _392149_392149 ; 
   reg __392149_392149;
   reg _392150_392150 ; 
   reg __392150_392150;
   reg _392151_392151 ; 
   reg __392151_392151;
   reg _392152_392152 ; 
   reg __392152_392152;
   reg _392153_392153 ; 
   reg __392153_392153;
   reg _392154_392154 ; 
   reg __392154_392154;
   reg _392155_392155 ; 
   reg __392155_392155;
   reg _392156_392156 ; 
   reg __392156_392156;
   reg _392157_392157 ; 
   reg __392157_392157;
   reg _392158_392158 ; 
   reg __392158_392158;
   reg _392159_392159 ; 
   reg __392159_392159;
   reg _392160_392160 ; 
   reg __392160_392160;
   reg _392161_392161 ; 
   reg __392161_392161;
   reg _392162_392162 ; 
   reg __392162_392162;
   reg _392163_392163 ; 
   reg __392163_392163;
   reg _392164_392164 ; 
   reg __392164_392164;
   reg _392165_392165 ; 
   reg __392165_392165;
   reg _392166_392166 ; 
   reg __392166_392166;
   reg _392167_392167 ; 
   reg __392167_392167;
   reg _392168_392168 ; 
   reg __392168_392168;
   reg _392169_392169 ; 
   reg __392169_392169;
   reg _392170_392170 ; 
   reg __392170_392170;
   reg _392171_392171 ; 
   reg __392171_392171;
   reg _392172_392172 ; 
   reg __392172_392172;
   reg _392173_392173 ; 
   reg __392173_392173;
   reg _392174_392174 ; 
   reg __392174_392174;
   reg _392175_392175 ; 
   reg __392175_392175;
   reg _392176_392176 ; 
   reg __392176_392176;
   reg _392177_392177 ; 
   reg __392177_392177;
   reg _392178_392178 ; 
   reg __392178_392178;
   reg _392179_392179 ; 
   reg __392179_392179;
   reg _392180_392180 ; 
   reg __392180_392180;
   reg _392181_392181 ; 
   reg __392181_392181;
   reg _392182_392182 ; 
   reg __392182_392182;
   reg _392183_392183 ; 
   reg __392183_392183;
   reg _392184_392184 ; 
   reg __392184_392184;
   reg _392185_392185 ; 
   reg __392185_392185;
   reg _392186_392186 ; 
   reg __392186_392186;
   reg _392187_392187 ; 
   reg __392187_392187;
   reg _392188_392188 ; 
   reg __392188_392188;
   reg _392189_392189 ; 
   reg __392189_392189;
   reg _392190_392190 ; 
   reg __392190_392190;
   reg _392191_392191 ; 
   reg __392191_392191;
   reg _392192_392192 ; 
   reg __392192_392192;
   reg _392193_392193 ; 
   reg __392193_392193;
   reg _392194_392194 ; 
   reg __392194_392194;
   reg _392195_392195 ; 
   reg __392195_392195;
   reg _392196_392196 ; 
   reg __392196_392196;
   reg _392197_392197 ; 
   reg __392197_392197;
   reg _392198_392198 ; 
   reg __392198_392198;
   reg _392199_392199 ; 
   reg __392199_392199;
   reg _392200_392200 ; 
   reg __392200_392200;
   reg _392201_392201 ; 
   reg __392201_392201;
   reg _392202_392202 ; 
   reg __392202_392202;
   reg _392203_392203 ; 
   reg __392203_392203;
   reg _392204_392204 ; 
   reg __392204_392204;
   reg _392205_392205 ; 
   reg __392205_392205;
   reg _392206_392206 ; 
   reg __392206_392206;
   reg _392207_392207 ; 
   reg __392207_392207;
   reg _392208_392208 ; 
   reg __392208_392208;
   reg _392209_392209 ; 
   reg __392209_392209;
   reg _392210_392210 ; 
   reg __392210_392210;
   reg _392211_392211 ; 
   reg __392211_392211;
   reg _392212_392212 ; 
   reg __392212_392212;
   reg _392213_392213 ; 
   reg __392213_392213;
   reg _392214_392214 ; 
   reg __392214_392214;
   reg _392215_392215 ; 
   reg __392215_392215;
   reg _392216_392216 ; 
   reg __392216_392216;
   reg _392217_392217 ; 
   reg __392217_392217;
   reg _392218_392218 ; 
   reg __392218_392218;
   reg _392219_392219 ; 
   reg __392219_392219;
   reg _392220_392220 ; 
   reg __392220_392220;
   reg _392221_392221 ; 
   reg __392221_392221;
   reg _392222_392222 ; 
   reg __392222_392222;
   reg _392223_392223 ; 
   reg __392223_392223;
   reg _392224_392224 ; 
   reg __392224_392224;
   reg _392225_392225 ; 
   reg __392225_392225;
   reg _392226_392226 ; 
   reg __392226_392226;
   reg _392227_392227 ; 
   reg __392227_392227;
   reg _392228_392228 ; 
   reg __392228_392228;
   reg _392229_392229 ; 
   reg __392229_392229;
   reg _392230_392230 ; 
   reg __392230_392230;
   reg _392231_392231 ; 
   reg __392231_392231;
   reg _392232_392232 ; 
   reg __392232_392232;
   reg _392233_392233 ; 
   reg __392233_392233;
   reg _392234_392234 ; 
   reg __392234_392234;
   reg _392235_392235 ; 
   reg __392235_392235;
   reg _392236_392236 ; 
   reg __392236_392236;
   reg _392237_392237 ; 
   reg __392237_392237;
   reg _392238_392238 ; 
   reg __392238_392238;
   reg _392239_392239 ; 
   reg __392239_392239;
   reg _392240_392240 ; 
   reg __392240_392240;
   reg _392241_392241 ; 
   reg __392241_392241;
   reg _392242_392242 ; 
   reg __392242_392242;
   reg _392243_392243 ; 
   reg __392243_392243;
   reg _392244_392244 ; 
   reg __392244_392244;
   reg _392245_392245 ; 
   reg __392245_392245;
   reg _392246_392246 ; 
   reg __392246_392246;
   reg _392247_392247 ; 
   reg __392247_392247;
   reg _392248_392248 ; 
   reg __392248_392248;
   reg _392249_392249 ; 
   reg __392249_392249;
   reg _392250_392250 ; 
   reg __392250_392250;
   reg _392251_392251 ; 
   reg __392251_392251;
   reg _392252_392252 ; 
   reg __392252_392252;
   reg _392253_392253 ; 
   reg __392253_392253;
   reg _392254_392254 ; 
   reg __392254_392254;
   reg _392255_392255 ; 
   reg __392255_392255;
   reg _392256_392256 ; 
   reg __392256_392256;
   reg _392257_392257 ; 
   reg __392257_392257;
   reg _392258_392258 ; 
   reg __392258_392258;
   reg _392259_392259 ; 
   reg __392259_392259;
   reg _392260_392260 ; 
   reg __392260_392260;
   reg _392261_392261 ; 
   reg __392261_392261;
   reg _392262_392262 ; 
   reg __392262_392262;
   reg _392263_392263 ; 
   reg __392263_392263;
   reg _392264_392264 ; 
   reg __392264_392264;
   reg _392265_392265 ; 
   reg __392265_392265;
   reg _392266_392266 ; 
   reg __392266_392266;
   reg _392267_392267 ; 
   reg __392267_392267;
   reg _392268_392268 ; 
   reg __392268_392268;
   reg _392269_392269 ; 
   reg __392269_392269;
   reg _392270_392270 ; 
   reg __392270_392270;
   reg _392271_392271 ; 
   reg __392271_392271;
   reg _392272_392272 ; 
   reg __392272_392272;
   reg _392273_392273 ; 
   reg __392273_392273;
   reg _392274_392274 ; 
   reg __392274_392274;
   reg _392275_392275 ; 
   reg __392275_392275;
   reg _392276_392276 ; 
   reg __392276_392276;
   reg _392277_392277 ; 
   reg __392277_392277;
   reg _392278_392278 ; 
   reg __392278_392278;
   reg _392279_392279 ; 
   reg __392279_392279;
   reg _392280_392280 ; 
   reg __392280_392280;
   reg _392281_392281 ; 
   reg __392281_392281;
   reg _392282_392282 ; 
   reg __392282_392282;
   reg _392283_392283 ; 
   reg __392283_392283;
   reg _392284_392284 ; 
   reg __392284_392284;
   reg _392285_392285 ; 
   reg __392285_392285;
   reg _392286_392286 ; 
   reg __392286_392286;
   reg _392287_392287 ; 
   reg __392287_392287;
   reg _392288_392288 ; 
   reg __392288_392288;
   reg _392289_392289 ; 
   reg __392289_392289;
   reg _392290_392290 ; 
   reg __392290_392290;
   reg _392291_392291 ; 
   reg __392291_392291;
   reg _392292_392292 ; 
   reg __392292_392292;
   reg _392293_392293 ; 
   reg __392293_392293;
   reg _392294_392294 ; 
   reg __392294_392294;
   reg _392295_392295 ; 
   reg __392295_392295;
   reg _392296_392296 ; 
   reg __392296_392296;
   reg _392297_392297 ; 
   reg __392297_392297;
   reg _392298_392298 ; 
   reg __392298_392298;
   reg _392299_392299 ; 
   reg __392299_392299;
   reg _392300_392300 ; 
   reg __392300_392300;
   reg _392301_392301 ; 
   reg __392301_392301;
   reg _392302_392302 ; 
   reg __392302_392302;
   reg _392303_392303 ; 
   reg __392303_392303;
   reg _392304_392304 ; 
   reg __392304_392304;
   reg _392305_392305 ; 
   reg __392305_392305;
   reg _392306_392306 ; 
   reg __392306_392306;
   reg _392307_392307 ; 
   reg __392307_392307;
   reg _392308_392308 ; 
   reg __392308_392308;
   reg _392309_392309 ; 
   reg __392309_392309;
   reg _392310_392310 ; 
   reg __392310_392310;
   reg _392311_392311 ; 
   reg __392311_392311;
   reg _392312_392312 ; 
   reg __392312_392312;
   reg _392313_392313 ; 
   reg __392313_392313;
   reg _392314_392314 ; 
   reg __392314_392314;
   reg _392315_392315 ; 
   reg __392315_392315;
   reg _392316_392316 ; 
   reg __392316_392316;
   reg _392317_392317 ; 
   reg __392317_392317;
   reg _392318_392318 ; 
   reg __392318_392318;
   reg _392319_392319 ; 
   reg __392319_392319;
   reg _392320_392320 ; 
   reg __392320_392320;
   reg _392321_392321 ; 
   reg __392321_392321;
   reg _392322_392322 ; 
   reg __392322_392322;
   reg _392323_392323 ; 
   reg __392323_392323;
   reg _392324_392324 ; 
   reg __392324_392324;
   reg _392325_392325 ; 
   reg __392325_392325;
   reg _392326_392326 ; 
   reg __392326_392326;
   reg _392327_392327 ; 
   reg __392327_392327;
   reg _392328_392328 ; 
   reg __392328_392328;
   reg _392329_392329 ; 
   reg __392329_392329;
   reg _392330_392330 ; 
   reg __392330_392330;
   reg _392331_392331 ; 
   reg __392331_392331;
   reg _392332_392332 ; 
   reg __392332_392332;
   reg _392333_392333 ; 
   reg __392333_392333;
   reg _392334_392334 ; 
   reg __392334_392334;
   reg _392335_392335 ; 
   reg __392335_392335;
   reg _392336_392336 ; 
   reg __392336_392336;
   reg _392337_392337 ; 
   reg __392337_392337;
   reg _392338_392338 ; 
   reg __392338_392338;
   reg _392339_392339 ; 
   reg __392339_392339;
   reg _392340_392340 ; 
   reg __392340_392340;
   reg _392341_392341 ; 
   reg __392341_392341;
   reg _392342_392342 ; 
   reg __392342_392342;
   reg _392343_392343 ; 
   reg __392343_392343;
   reg _392344_392344 ; 
   reg __392344_392344;
   reg _392345_392345 ; 
   reg __392345_392345;
   reg _392346_392346 ; 
   reg __392346_392346;
   reg _392347_392347 ; 
   reg __392347_392347;
   reg _392348_392348 ; 
   reg __392348_392348;
   reg _392349_392349 ; 
   reg __392349_392349;
   reg _392350_392350 ; 
   reg __392350_392350;
   reg _392351_392351 ; 
   reg __392351_392351;
   reg _392352_392352 ; 
   reg __392352_392352;
   reg _392353_392353 ; 
   reg __392353_392353;
   reg _392354_392354 ; 
   reg __392354_392354;
   reg _392355_392355 ; 
   reg __392355_392355;
   reg _392356_392356 ; 
   reg __392356_392356;
   reg _392357_392357 ; 
   reg __392357_392357;
   reg _392358_392358 ; 
   reg __392358_392358;
   reg _392359_392359 ; 
   reg __392359_392359;
   reg _392360_392360 ; 
   reg __392360_392360;
   reg _392361_392361 ; 
   reg __392361_392361;
   reg _392362_392362 ; 
   reg __392362_392362;
   reg _392363_392363 ; 
   reg __392363_392363;
   reg _392364_392364 ; 
   reg __392364_392364;
   reg _392365_392365 ; 
   reg __392365_392365;
   reg _392366_392366 ; 
   reg __392366_392366;
   reg _392367_392367 ; 
   reg __392367_392367;
   reg _392368_392368 ; 
   reg __392368_392368;
   reg _392369_392369 ; 
   reg __392369_392369;
   reg _392370_392370 ; 
   reg __392370_392370;
   reg _392371_392371 ; 
   reg __392371_392371;
   reg _392372_392372 ; 
   reg __392372_392372;
   reg _392373_392373 ; 
   reg __392373_392373;
   reg _392374_392374 ; 
   reg __392374_392374;
   reg _392375_392375 ; 
   reg __392375_392375;
   reg _392376_392376 ; 
   reg __392376_392376;
   reg _392377_392377 ; 
   reg __392377_392377;
   reg _392378_392378 ; 
   reg __392378_392378;
   reg _392379_392379 ; 
   reg __392379_392379;
   reg _392380_392380 ; 
   reg __392380_392380;
   reg _392381_392381 ; 
   reg __392381_392381;
   reg _392382_392382 ; 
   reg __392382_392382;
   reg _392383_392383 ; 
   reg __392383_392383;
   reg _392384_392384 ; 
   reg __392384_392384;
   reg _392385_392385 ; 
   reg __392385_392385;
   reg _392386_392386 ; 
   reg __392386_392386;
   reg _392387_392387 ; 
   reg __392387_392387;
   reg _392388_392388 ; 
   reg __392388_392388;
   reg _392389_392389 ; 
   reg __392389_392389;
   reg _392390_392390 ; 
   reg __392390_392390;
   reg _392391_392391 ; 
   reg __392391_392391;
   reg _392392_392392 ; 
   reg __392392_392392;
   reg _392393_392393 ; 
   reg __392393_392393;
   reg _392394_392394 ; 
   reg __392394_392394;
   reg _392395_392395 ; 
   reg __392395_392395;
   reg _392396_392396 ; 
   reg __392396_392396;
   reg _392397_392397 ; 
   reg __392397_392397;
   reg _392398_392398 ; 
   reg __392398_392398;
   reg _392399_392399 ; 
   reg __392399_392399;
   reg _392400_392400 ; 
   reg __392400_392400;
   reg _392401_392401 ; 
   reg __392401_392401;
   reg _392402_392402 ; 
   reg __392402_392402;
   reg _392403_392403 ; 
   reg __392403_392403;
   reg _392404_392404 ; 
   reg __392404_392404;
   reg _392405_392405 ; 
   reg __392405_392405;
   reg _392406_392406 ; 
   reg __392406_392406;
   reg _392407_392407 ; 
   reg __392407_392407;
   reg _392408_392408 ; 
   reg __392408_392408;
   reg _392409_392409 ; 
   reg __392409_392409;
   reg _392410_392410 ; 
   reg __392410_392410;
   reg _392411_392411 ; 
   reg __392411_392411;
   reg _392412_392412 ; 
   reg __392412_392412;
   reg _392413_392413 ; 
   reg __392413_392413;
   reg _392414_392414 ; 
   reg __392414_392414;
   reg _392415_392415 ; 
   reg __392415_392415;
   reg _392416_392416 ; 
   reg __392416_392416;
   reg _392417_392417 ; 
   reg __392417_392417;
   reg _392418_392418 ; 
   reg __392418_392418;
   reg _392419_392419 ; 
   reg __392419_392419;
   reg _392420_392420 ; 
   reg __392420_392420;
   reg _392421_392421 ; 
   reg __392421_392421;
   reg _392422_392422 ; 
   reg __392422_392422;
   reg _392423_392423 ; 
   reg __392423_392423;
   reg _392424_392424 ; 
   reg __392424_392424;
   reg _392425_392425 ; 
   reg __392425_392425;
   reg _392426_392426 ; 
   reg __392426_392426;
   reg _392427_392427 ; 
   reg __392427_392427;
   reg _392428_392428 ; 
   reg __392428_392428;
   reg _392429_392429 ; 
   reg __392429_392429;
   reg _392430_392430 ; 
   reg __392430_392430;
   reg _392431_392431 ; 
   reg __392431_392431;
   reg _392432_392432 ; 
   reg __392432_392432;
   reg _392433_392433 ; 
   reg __392433_392433;
   reg _392434_392434 ; 
   reg __392434_392434;
   reg _392435_392435 ; 
   reg __392435_392435;
   reg _392436_392436 ; 
   reg __392436_392436;
   reg _392437_392437 ; 
   reg __392437_392437;
   reg _392438_392438 ; 
   reg __392438_392438;
   reg _392439_392439 ; 
   reg __392439_392439;
   reg _392440_392440 ; 
   reg __392440_392440;
   reg _392441_392441 ; 
   reg __392441_392441;
   reg _392442_392442 ; 
   reg __392442_392442;
   reg _392443_392443 ; 
   reg __392443_392443;
   reg _392444_392444 ; 
   reg __392444_392444;
   reg _392445_392445 ; 
   reg __392445_392445;
   reg _392446_392446 ; 
   reg __392446_392446;
   reg _392447_392447 ; 
   reg __392447_392447;
   reg _392448_392448 ; 
   reg __392448_392448;
   reg _392449_392449 ; 
   reg __392449_392449;
   reg _392450_392450 ; 
   reg __392450_392450;
   reg _392451_392451 ; 
   reg __392451_392451;
   reg _392452_392452 ; 
   reg __392452_392452;
   reg _392453_392453 ; 
   reg __392453_392453;
   reg _392454_392454 ; 
   reg __392454_392454;
   reg _392455_392455 ; 
   reg __392455_392455;
   reg _392456_392456 ; 
   reg __392456_392456;
   reg _392457_392457 ; 
   reg __392457_392457;
   reg _392458_392458 ; 
   reg __392458_392458;
   reg _392459_392459 ; 
   reg __392459_392459;
   reg _392460_392460 ; 
   reg __392460_392460;
   reg _392461_392461 ; 
   reg __392461_392461;
   reg _392462_392462 ; 
   reg __392462_392462;
   reg _392463_392463 ; 
   reg __392463_392463;
   reg _392464_392464 ; 
   reg __392464_392464;
   reg _392465_392465 ; 
   reg __392465_392465;
   reg _392466_392466 ; 
   reg __392466_392466;
   reg _392467_392467 ; 
   reg __392467_392467;
   reg _392468_392468 ; 
   reg __392468_392468;
   reg _392469_392469 ; 
   reg __392469_392469;
   reg _392470_392470 ; 
   reg __392470_392470;
   reg _392471_392471 ; 
   reg __392471_392471;
   reg _392472_392472 ; 
   reg __392472_392472;
   reg _392473_392473 ; 
   reg __392473_392473;
   reg _392474_392474 ; 
   reg __392474_392474;
   reg _392475_392475 ; 
   reg __392475_392475;
   reg _392476_392476 ; 
   reg __392476_392476;
   reg _392477_392477 ; 
   reg __392477_392477;
   reg _392478_392478 ; 
   reg __392478_392478;
   reg _392479_392479 ; 
   reg __392479_392479;
   reg _392480_392480 ; 
   reg __392480_392480;
   reg _392481_392481 ; 
   reg __392481_392481;
   reg _392482_392482 ; 
   reg __392482_392482;
   reg _392483_392483 ; 
   reg __392483_392483;
   reg _392484_392484 ; 
   reg __392484_392484;
   reg _392485_392485 ; 
   reg __392485_392485;
   reg _392486_392486 ; 
   reg __392486_392486;
   reg _392487_392487 ; 
   reg __392487_392487;
   reg _392488_392488 ; 
   reg __392488_392488;
   reg _392489_392489 ; 
   reg __392489_392489;
   reg _392490_392490 ; 
   reg __392490_392490;
   reg _392491_392491 ; 
   reg __392491_392491;
   reg _392492_392492 ; 
   reg __392492_392492;
   reg _392493_392493 ; 
   reg __392493_392493;
   reg _392494_392494 ; 
   reg __392494_392494;
   reg _392495_392495 ; 
   reg __392495_392495;
   reg _392496_392496 ; 
   reg __392496_392496;
   reg _392497_392497 ; 
   reg __392497_392497;
   reg _392498_392498 ; 
   reg __392498_392498;
   reg _392499_392499 ; 
   reg __392499_392499;
   reg _392500_392500 ; 
   reg __392500_392500;
   reg _392501_392501 ; 
   reg __392501_392501;
   reg _392502_392502 ; 
   reg __392502_392502;
   reg _392503_392503 ; 
   reg __392503_392503;
   reg _392504_392504 ; 
   reg __392504_392504;
   reg _392505_392505 ; 
   reg __392505_392505;
   reg _392506_392506 ; 
   reg __392506_392506;
   reg _392507_392507 ; 
   reg __392507_392507;
   reg _392508_392508 ; 
   reg __392508_392508;
   reg _392509_392509 ; 
   reg __392509_392509;
   reg _392510_392510 ; 
   reg __392510_392510;
   reg _392511_392511 ; 
   reg __392511_392511;
   reg _392512_392512 ; 
   reg __392512_392512;
   reg _392513_392513 ; 
   reg __392513_392513;
   reg _392514_392514 ; 
   reg __392514_392514;
   reg _392515_392515 ; 
   reg __392515_392515;
   reg _392516_392516 ; 
   reg __392516_392516;
   reg _392517_392517 ; 
   reg __392517_392517;
   reg _392518_392518 ; 
   reg __392518_392518;
   reg _392519_392519 ; 
   reg __392519_392519;
   reg _392520_392520 ; 
   reg __392520_392520;
   reg _392521_392521 ; 
   reg __392521_392521;
   reg _392522_392522 ; 
   reg __392522_392522;
   reg _392523_392523 ; 
   reg __392523_392523;
   reg _392524_392524 ; 
   reg __392524_392524;
   reg _392525_392525 ; 
   reg __392525_392525;
   reg _392526_392526 ; 
   reg __392526_392526;
   reg _392527_392527 ; 
   reg __392527_392527;
   reg _392528_392528 ; 
   reg __392528_392528;
   reg _392529_392529 ; 
   reg __392529_392529;
   reg _392530_392530 ; 
   reg __392530_392530;
   reg _392531_392531 ; 
   reg __392531_392531;
   reg _392532_392532 ; 
   reg __392532_392532;
   reg _392533_392533 ; 
   reg __392533_392533;
   reg _392534_392534 ; 
   reg __392534_392534;
   reg _392535_392535 ; 
   reg __392535_392535;
   reg _392536_392536 ; 
   reg __392536_392536;
   reg _392537_392537 ; 
   reg __392537_392537;
   reg _392538_392538 ; 
   reg __392538_392538;
   reg _392539_392539 ; 
   reg __392539_392539;
   reg _392540_392540 ; 
   reg __392540_392540;
   reg _392541_392541 ; 
   reg __392541_392541;
   reg _392542_392542 ; 
   reg __392542_392542;
   reg _392543_392543 ; 
   reg __392543_392543;
   reg _392544_392544 ; 
   reg __392544_392544;
   reg _392545_392545 ; 
   reg __392545_392545;
   reg _392546_392546 ; 
   reg __392546_392546;
   reg _392547_392547 ; 
   reg __392547_392547;
   reg _392548_392548 ; 
   reg __392548_392548;
   reg _392549_392549 ; 
   reg __392549_392549;
   reg _392550_392550 ; 
   reg __392550_392550;
   reg _392551_392551 ; 
   reg __392551_392551;
   reg _392552_392552 ; 
   reg __392552_392552;
   reg _392553_392553 ; 
   reg __392553_392553;
   reg _392554_392554 ; 
   reg __392554_392554;
   reg _392555_392555 ; 
   reg __392555_392555;
   reg _392556_392556 ; 
   reg __392556_392556;
   reg _392557_392557 ; 
   reg __392557_392557;
   reg _392558_392558 ; 
   reg __392558_392558;
   reg _392559_392559 ; 
   reg __392559_392559;
   reg _392560_392560 ; 
   reg __392560_392560;
   reg _392561_392561 ; 
   reg __392561_392561;
   reg _392562_392562 ; 
   reg __392562_392562;
   reg _392563_392563 ; 
   reg __392563_392563;
   reg _392564_392564 ; 
   reg __392564_392564;
   reg _392565_392565 ; 
   reg __392565_392565;
   reg _392566_392566 ; 
   reg __392566_392566;
   reg _392567_392567 ; 
   reg __392567_392567;
   reg _392568_392568 ; 
   reg __392568_392568;
   reg _392569_392569 ; 
   reg __392569_392569;
   reg _392570_392570 ; 
   reg __392570_392570;
   reg _392571_392571 ; 
   reg __392571_392571;
   reg _392572_392572 ; 
   reg __392572_392572;
   reg _392573_392573 ; 
   reg __392573_392573;
   reg _392574_392574 ; 
   reg __392574_392574;
   reg _392575_392575 ; 
   reg __392575_392575;
   reg _392576_392576 ; 
   reg __392576_392576;
   reg _392577_392577 ; 
   reg __392577_392577;
   reg _392578_392578 ; 
   reg __392578_392578;
   reg _392579_392579 ; 
   reg __392579_392579;
   reg _392580_392580 ; 
   reg __392580_392580;
   reg _392581_392581 ; 
   reg __392581_392581;
   reg _392582_392582 ; 
   reg __392582_392582;
   reg _392583_392583 ; 
   reg __392583_392583;
   reg _392584_392584 ; 
   reg __392584_392584;
   reg _392585_392585 ; 
   reg __392585_392585;
   reg _392586_392586 ; 
   reg __392586_392586;
   reg _392587_392587 ; 
   reg __392587_392587;
   reg _392588_392588 ; 
   reg __392588_392588;
   reg _392589_392589 ; 
   reg __392589_392589;
   reg _392590_392590 ; 
   reg __392590_392590;
   reg _392591_392591 ; 
   reg __392591_392591;
   reg _392592_392592 ; 
   reg __392592_392592;
   reg _392593_392593 ; 
   reg __392593_392593;
   reg _392594_392594 ; 
   reg __392594_392594;
   reg _392595_392595 ; 
   reg __392595_392595;
   reg _392596_392596 ; 
   reg __392596_392596;
   reg _392597_392597 ; 
   reg __392597_392597;
   reg _392598_392598 ; 
   reg __392598_392598;
   reg _392599_392599 ; 
   reg __392599_392599;
   reg _392600_392600 ; 
   reg __392600_392600;
   reg _392601_392601 ; 
   reg __392601_392601;
   reg _392602_392602 ; 
   reg __392602_392602;
   reg _392603_392603 ; 
   reg __392603_392603;
   reg _392604_392604 ; 
   reg __392604_392604;
   reg _392605_392605 ; 
   reg __392605_392605;
   reg _392606_392606 ; 
   reg __392606_392606;
   reg _392607_392607 ; 
   reg __392607_392607;
   reg _392608_392608 ; 
   reg __392608_392608;
   reg _392609_392609 ; 
   reg __392609_392609;
   reg _392610_392610 ; 
   reg __392610_392610;
   reg _392611_392611 ; 
   reg __392611_392611;
   reg _392612_392612 ; 
   reg __392612_392612;
   reg _392613_392613 ; 
   reg __392613_392613;
   reg _392614_392614 ; 
   reg __392614_392614;
   reg _392615_392615 ; 
   reg __392615_392615;
   reg _392616_392616 ; 
   reg __392616_392616;
   reg _392617_392617 ; 
   reg __392617_392617;
   reg _392618_392618 ; 
   reg __392618_392618;
   reg _392619_392619 ; 
   reg __392619_392619;
   reg _392620_392620 ; 
   reg __392620_392620;
   reg _392621_392621 ; 
   reg __392621_392621;
   reg _392622_392622 ; 
   reg __392622_392622;
   reg _392623_392623 ; 
   reg __392623_392623;
   reg _392624_392624 ; 
   reg __392624_392624;
   reg _392625_392625 ; 
   reg __392625_392625;
   reg _392626_392626 ; 
   reg __392626_392626;
   reg _392627_392627 ; 
   reg __392627_392627;
   reg _392628_392628 ; 
   reg __392628_392628;
   reg _392629_392629 ; 
   reg __392629_392629;
   reg _392630_392630 ; 
   reg __392630_392630;
   reg _392631_392631 ; 
   reg __392631_392631;
   reg _392632_392632 ; 
   reg __392632_392632;
   reg _392633_392633 ; 
   reg __392633_392633;
   reg _392634_392634 ; 
   reg __392634_392634;
   reg _392635_392635 ; 
   reg __392635_392635;
   reg _392636_392636 ; 
   reg __392636_392636;
   reg _392637_392637 ; 
   reg __392637_392637;
   reg _392638_392638 ; 
   reg __392638_392638;
   reg _392639_392639 ; 
   reg __392639_392639;
   reg _392640_392640 ; 
   reg __392640_392640;
   reg _392641_392641 ; 
   reg __392641_392641;
   reg _392642_392642 ; 
   reg __392642_392642;
   reg _392643_392643 ; 
   reg __392643_392643;
   reg _392644_392644 ; 
   reg __392644_392644;
   reg _392645_392645 ; 
   reg __392645_392645;
   reg _392646_392646 ; 
   reg __392646_392646;
   reg _392647_392647 ; 
   reg __392647_392647;
   reg _392648_392648 ; 
   reg __392648_392648;
   reg _392649_392649 ; 
   reg __392649_392649;
   reg _392650_392650 ; 
   reg __392650_392650;
   reg _392651_392651 ; 
   reg __392651_392651;
   reg _392652_392652 ; 
   reg __392652_392652;
   reg _392653_392653 ; 
   reg __392653_392653;
   reg _392654_392654 ; 
   reg __392654_392654;
   reg _392655_392655 ; 
   reg __392655_392655;
   reg _392656_392656 ; 
   reg __392656_392656;
   reg _392657_392657 ; 
   reg __392657_392657;
   reg _392658_392658 ; 
   reg __392658_392658;
   reg _392659_392659 ; 
   reg __392659_392659;
   reg _392660_392660 ; 
   reg __392660_392660;
   reg _392661_392661 ; 
   reg __392661_392661;
   reg _392662_392662 ; 
   reg __392662_392662;
   reg _392663_392663 ; 
   reg __392663_392663;
   reg _392664_392664 ; 
   reg __392664_392664;
   reg _392665_392665 ; 
   reg __392665_392665;
   reg _392666_392666 ; 
   reg __392666_392666;
   reg _392667_392667 ; 
   reg __392667_392667;
   reg _392668_392668 ; 
   reg __392668_392668;
   reg _392669_392669 ; 
   reg __392669_392669;
   reg _392670_392670 ; 
   reg __392670_392670;
   reg _392671_392671 ; 
   reg __392671_392671;
   reg _392672_392672 ; 
   reg __392672_392672;
   reg _392673_392673 ; 
   reg __392673_392673;
   reg _392674_392674 ; 
   reg __392674_392674;
   reg _392675_392675 ; 
   reg __392675_392675;
   reg _392676_392676 ; 
   reg __392676_392676;
   reg _392677_392677 ; 
   reg __392677_392677;
   reg _392678_392678 ; 
   reg __392678_392678;
   reg _392679_392679 ; 
   reg __392679_392679;
   reg _392680_392680 ; 
   reg __392680_392680;
   reg _392681_392681 ; 
   reg __392681_392681;
   reg _392682_392682 ; 
   reg __392682_392682;
   reg _392683_392683 ; 
   reg __392683_392683;
   reg _392684_392684 ; 
   reg __392684_392684;
   reg _392685_392685 ; 
   reg __392685_392685;
   reg _392686_392686 ; 
   reg __392686_392686;
   reg _392687_392687 ; 
   reg __392687_392687;
   reg _392688_392688 ; 
   reg __392688_392688;
   reg _392689_392689 ; 
   reg __392689_392689;
   reg _392690_392690 ; 
   reg __392690_392690;
   reg _392691_392691 ; 
   reg __392691_392691;
   reg _392692_392692 ; 
   reg __392692_392692;
   reg _392693_392693 ; 
   reg __392693_392693;
   reg _392694_392694 ; 
   reg __392694_392694;
   reg _392695_392695 ; 
   reg __392695_392695;
   reg _392696_392696 ; 
   reg __392696_392696;
   reg _392697_392697 ; 
   reg __392697_392697;
   reg _392698_392698 ; 
   reg __392698_392698;
   reg _392699_392699 ; 
   reg __392699_392699;
   reg _392700_392700 ; 
   reg __392700_392700;
   reg _392701_392701 ; 
   reg __392701_392701;
   reg _392702_392702 ; 
   reg __392702_392702;
   reg _392703_392703 ; 
   reg __392703_392703;
   reg _392704_392704 ; 
   reg __392704_392704;
   reg _392705_392705 ; 
   reg __392705_392705;
   reg _392706_392706 ; 
   reg __392706_392706;
   reg _392707_392707 ; 
   reg __392707_392707;
   reg _392708_392708 ; 
   reg __392708_392708;
   reg _392709_392709 ; 
   reg __392709_392709;
   reg _392710_392710 ; 
   reg __392710_392710;
   reg _392711_392711 ; 
   reg __392711_392711;
   reg _392712_392712 ; 
   reg __392712_392712;
   reg _392713_392713 ; 
   reg __392713_392713;
   reg _392714_392714 ; 
   reg __392714_392714;
   reg _392715_392715 ; 
   reg __392715_392715;
   reg _392716_392716 ; 
   reg __392716_392716;
   reg _392717_392717 ; 
   reg __392717_392717;
   reg _392718_392718 ; 
   reg __392718_392718;
   reg _392719_392719 ; 
   reg __392719_392719;
   reg _392720_392720 ; 
   reg __392720_392720;
   reg _392721_392721 ; 
   reg __392721_392721;
   reg _392722_392722 ; 
   reg __392722_392722;
   reg _392723_392723 ; 
   reg __392723_392723;
   reg _392724_392724 ; 
   reg __392724_392724;
   reg _392725_392725 ; 
   reg __392725_392725;
   reg _392726_392726 ; 
   reg __392726_392726;
   reg _392727_392727 ; 
   reg __392727_392727;
   reg _392728_392728 ; 
   reg __392728_392728;
   reg _392729_392729 ; 
   reg __392729_392729;
   reg _392730_392730 ; 
   reg __392730_392730;
   reg _392731_392731 ; 
   reg __392731_392731;
   reg _392732_392732 ; 
   reg __392732_392732;
   reg _392733_392733 ; 
   reg __392733_392733;
   reg _392734_392734 ; 
   reg __392734_392734;
   reg _392735_392735 ; 
   reg __392735_392735;
   reg _392736_392736 ; 
   reg __392736_392736;
   reg _392737_392737 ; 
   reg __392737_392737;
   reg _392738_392738 ; 
   reg __392738_392738;
   reg _392739_392739 ; 
   reg __392739_392739;
   reg _392740_392740 ; 
   reg __392740_392740;
   reg _392741_392741 ; 
   reg __392741_392741;
   reg _392742_392742 ; 
   reg __392742_392742;
   reg _392743_392743 ; 
   reg __392743_392743;
   reg _392744_392744 ; 
   reg __392744_392744;
   reg _392745_392745 ; 
   reg __392745_392745;
   reg _392746_392746 ; 
   reg __392746_392746;
   reg _392747_392747 ; 
   reg __392747_392747;
   reg _392748_392748 ; 
   reg __392748_392748;
   reg _392749_392749 ; 
   reg __392749_392749;
   reg _392750_392750 ; 
   reg __392750_392750;
   reg _392751_392751 ; 
   reg __392751_392751;
   reg _392752_392752 ; 
   reg __392752_392752;
   reg _392753_392753 ; 
   reg __392753_392753;
   reg _392754_392754 ; 
   reg __392754_392754;
   reg _392755_392755 ; 
   reg __392755_392755;
   reg _392756_392756 ; 
   reg __392756_392756;
   reg _392757_392757 ; 
   reg __392757_392757;
   reg _392758_392758 ; 
   reg __392758_392758;
   reg _392759_392759 ; 
   reg __392759_392759;
   reg _392760_392760 ; 
   reg __392760_392760;
   reg _392761_392761 ; 
   reg __392761_392761;
   reg _392762_392762 ; 
   reg __392762_392762;
   reg _392763_392763 ; 
   reg __392763_392763;
   reg _392764_392764 ; 
   reg __392764_392764;
   reg _392765_392765 ; 
   reg __392765_392765;
   reg _392766_392766 ; 
   reg __392766_392766;
   reg _392767_392767 ; 
   reg __392767_392767;
   reg _392768_392768 ; 
   reg __392768_392768;
   reg _392769_392769 ; 
   reg __392769_392769;
   reg _392770_392770 ; 
   reg __392770_392770;
   reg _392771_392771 ; 
   reg __392771_392771;
   reg _392772_392772 ; 
   reg __392772_392772;
   reg _392773_392773 ; 
   reg __392773_392773;
   reg _392774_392774 ; 
   reg __392774_392774;
   reg _392775_392775 ; 
   reg __392775_392775;
   reg _392776_392776 ; 
   reg __392776_392776;
   reg _392777_392777 ; 
   reg __392777_392777;
   reg _392778_392778 ; 
   reg __392778_392778;
   reg _392779_392779 ; 
   reg __392779_392779;
   reg _392780_392780 ; 
   reg __392780_392780;
   reg _392781_392781 ; 
   reg __392781_392781;
   reg _392782_392782 ; 
   reg __392782_392782;
   reg _392783_392783 ; 
   reg __392783_392783;
   reg _392784_392784 ; 
   reg __392784_392784;
   reg _392785_392785 ; 
   reg __392785_392785;
   reg _392786_392786 ; 
   reg __392786_392786;
   reg _392787_392787 ; 
   reg __392787_392787;
   reg _392788_392788 ; 
   reg __392788_392788;
   reg _392789_392789 ; 
   reg __392789_392789;
   reg _392790_392790 ; 
   reg __392790_392790;
   reg _392791_392791 ; 
   reg __392791_392791;
   reg _392792_392792 ; 
   reg __392792_392792;
   reg _392793_392793 ; 
   reg __392793_392793;
   reg _392794_392794 ; 
   reg __392794_392794;
   reg _392795_392795 ; 
   reg __392795_392795;
   reg _392796_392796 ; 
   reg __392796_392796;
   reg _392797_392797 ; 
   reg __392797_392797;
   reg _392798_392798 ; 
   reg __392798_392798;
   reg _392799_392799 ; 
   reg __392799_392799;
   reg _392800_392800 ; 
   reg __392800_392800;
   reg _392801_392801 ; 
   reg __392801_392801;
   reg _392802_392802 ; 
   reg __392802_392802;
   reg _392803_392803 ; 
   reg __392803_392803;
   reg _392804_392804 ; 
   reg __392804_392804;
   reg _392805_392805 ; 
   reg __392805_392805;
   reg _392806_392806 ; 
   reg __392806_392806;
   reg _392807_392807 ; 
   reg __392807_392807;
   reg _392808_392808 ; 
   reg __392808_392808;
   reg _392809_392809 ; 
   reg __392809_392809;
   reg _392810_392810 ; 
   reg __392810_392810;
   reg _392811_392811 ; 
   reg __392811_392811;
   reg _392812_392812 ; 
   reg __392812_392812;
   reg _392813_392813 ; 
   reg __392813_392813;
   reg _392814_392814 ; 
   reg __392814_392814;
   reg _392815_392815 ; 
   reg __392815_392815;
   reg _392816_392816 ; 
   reg __392816_392816;
   reg _392817_392817 ; 
   reg __392817_392817;
   reg _392818_392818 ; 
   reg __392818_392818;
   reg _392819_392819 ; 
   reg __392819_392819;
   reg _392820_392820 ; 
   reg __392820_392820;
   reg _392821_392821 ; 
   reg __392821_392821;
   reg _392822_392822 ; 
   reg __392822_392822;
   reg _392823_392823 ; 
   reg __392823_392823;
   reg _392824_392824 ; 
   reg __392824_392824;
   reg _392825_392825 ; 
   reg __392825_392825;
   reg _392826_392826 ; 
   reg __392826_392826;
   reg _392827_392827 ; 
   reg __392827_392827;
   reg _392828_392828 ; 
   reg __392828_392828;
   reg _392829_392829 ; 
   reg __392829_392829;
   reg _392830_392830 ; 
   reg __392830_392830;
   reg _392831_392831 ; 
   reg __392831_392831;
   reg _392832_392832 ; 
   reg __392832_392832;
   reg _392833_392833 ; 
   reg __392833_392833;
   reg _392834_392834 ; 
   reg __392834_392834;
   reg _392835_392835 ; 
   reg __392835_392835;
   reg _392836_392836 ; 
   reg __392836_392836;
   reg _392837_392837 ; 
   reg __392837_392837;
   reg _392838_392838 ; 
   reg __392838_392838;
   reg _392839_392839 ; 
   reg __392839_392839;
   reg _392840_392840 ; 
   reg __392840_392840;
   reg _392841_392841 ; 
   reg __392841_392841;
   reg _392842_392842 ; 
   reg __392842_392842;
   reg _392843_392843 ; 
   reg __392843_392843;
   reg _392844_392844 ; 
   reg __392844_392844;
   reg _392845_392845 ; 
   reg __392845_392845;
   reg _392846_392846 ; 
   reg __392846_392846;
   reg _392847_392847 ; 
   reg __392847_392847;
   reg _392848_392848 ; 
   reg __392848_392848;
   reg _392849_392849 ; 
   reg __392849_392849;
   reg _392850_392850 ; 
   reg __392850_392850;
   reg _392851_392851 ; 
   reg __392851_392851;
   reg _392852_392852 ; 
   reg __392852_392852;
   reg _392853_392853 ; 
   reg __392853_392853;
   reg _392854_392854 ; 
   reg __392854_392854;
   reg _392855_392855 ; 
   reg __392855_392855;
   reg _392856_392856 ; 
   reg __392856_392856;
   reg _392857_392857 ; 
   reg __392857_392857;
   reg _392858_392858 ; 
   reg __392858_392858;
   reg _392859_392859 ; 
   reg __392859_392859;
   reg _392860_392860 ; 
   reg __392860_392860;
   reg _392861_392861 ; 
   reg __392861_392861;
   reg _392862_392862 ; 
   reg __392862_392862;
   reg _392863_392863 ; 
   reg __392863_392863;
   reg _392864_392864 ; 
   reg __392864_392864;
   reg _392865_392865 ; 
   reg __392865_392865;
   reg _392866_392866 ; 
   reg __392866_392866;
   reg _392867_392867 ; 
   reg __392867_392867;
   reg _392868_392868 ; 
   reg __392868_392868;
   reg _392869_392869 ; 
   reg __392869_392869;
   reg _392870_392870 ; 
   reg __392870_392870;
   reg _392871_392871 ; 
   reg __392871_392871;
   reg _392872_392872 ; 
   reg __392872_392872;
   reg _392873_392873 ; 
   reg __392873_392873;
   reg _392874_392874 ; 
   reg __392874_392874;
   reg _392875_392875 ; 
   reg __392875_392875;
   reg _392876_392876 ; 
   reg __392876_392876;
   reg _392877_392877 ; 
   reg __392877_392877;
   reg _392878_392878 ; 
   reg __392878_392878;
   reg _392879_392879 ; 
   reg __392879_392879;
   reg _392880_392880 ; 
   reg __392880_392880;
   reg _392881_392881 ; 
   reg __392881_392881;
   reg _392882_392882 ; 
   reg __392882_392882;
   reg _392883_392883 ; 
   reg __392883_392883;
   reg _392884_392884 ; 
   reg __392884_392884;
   reg _392885_392885 ; 
   reg __392885_392885;
   reg _392886_392886 ; 
   reg __392886_392886;
   reg _392887_392887 ; 
   reg __392887_392887;
   reg _392888_392888 ; 
   reg __392888_392888;
   reg _392889_392889 ; 
   reg __392889_392889;
   reg _392890_392890 ; 
   reg __392890_392890;
   reg _392891_392891 ; 
   reg __392891_392891;
   reg _392892_392892 ; 
   reg __392892_392892;
   reg _392893_392893 ; 
   reg __392893_392893;
   reg _392894_392894 ; 
   reg __392894_392894;
   reg _392895_392895 ; 
   reg __392895_392895;
   reg _392896_392896 ; 
   reg __392896_392896;
   reg _392897_392897 ; 
   reg __392897_392897;
   reg _392898_392898 ; 
   reg __392898_392898;
   reg _392899_392899 ; 
   reg __392899_392899;
   reg _392900_392900 ; 
   reg __392900_392900;
   reg _392901_392901 ; 
   reg __392901_392901;
   reg _392902_392902 ; 
   reg __392902_392902;
   reg _392903_392903 ; 
   reg __392903_392903;
   reg _392904_392904 ; 
   reg __392904_392904;
   reg _392905_392905 ; 
   reg __392905_392905;
   reg _392906_392906 ; 
   reg __392906_392906;
   reg _392907_392907 ; 
   reg __392907_392907;
   reg _392908_392908 ; 
   reg __392908_392908;
   reg _392909_392909 ; 
   reg __392909_392909;
   reg _392910_392910 ; 
   reg __392910_392910;
   reg _392911_392911 ; 
   reg __392911_392911;
   reg _392912_392912 ; 
   reg __392912_392912;
   reg _392913_392913 ; 
   reg __392913_392913;
   reg _392914_392914 ; 
   reg __392914_392914;
   reg _392915_392915 ; 
   reg __392915_392915;
   reg _392916_392916 ; 
   reg __392916_392916;
   reg _392917_392917 ; 
   reg __392917_392917;
   reg _392918_392918 ; 
   reg __392918_392918;
   reg _392919_392919 ; 
   reg __392919_392919;
   reg _392920_392920 ; 
   reg __392920_392920;
   reg _392921_392921 ; 
   reg __392921_392921;
   reg _392922_392922 ; 
   reg __392922_392922;
   reg _392923_392923 ; 
   reg __392923_392923;
   reg _392924_392924 ; 
   reg __392924_392924;
   reg _392925_392925 ; 
   reg __392925_392925;
   reg _392926_392926 ; 
   reg __392926_392926;
   reg _392927_392927 ; 
   reg __392927_392927;
   reg _392928_392928 ; 
   reg __392928_392928;
   reg _392929_392929 ; 
   reg __392929_392929;
   reg _392930_392930 ; 
   reg __392930_392930;
   reg _392931_392931 ; 
   reg __392931_392931;
   reg _392932_392932 ; 
   reg __392932_392932;
   reg _392933_392933 ; 
   reg __392933_392933;
   reg _392934_392934 ; 
   reg __392934_392934;
   reg _392935_392935 ; 
   reg __392935_392935;
   reg _392936_392936 ; 
   reg __392936_392936;
   reg _392937_392937 ; 
   reg __392937_392937;
   reg _392938_392938 ; 
   reg __392938_392938;
   reg _392939_392939 ; 
   reg __392939_392939;
   reg _392940_392940 ; 
   reg __392940_392940;
   reg _392941_392941 ; 
   reg __392941_392941;
   reg _392942_392942 ; 
   reg __392942_392942;
   reg _392943_392943 ; 
   reg __392943_392943;
   reg _392944_392944 ; 
   reg __392944_392944;
   reg _392945_392945 ; 
   reg __392945_392945;
   reg _392946_392946 ; 
   reg __392946_392946;
   reg _392947_392947 ; 
   reg __392947_392947;
   reg _392948_392948 ; 
   reg __392948_392948;
   reg _392949_392949 ; 
   reg __392949_392949;
   reg _392950_392950 ; 
   reg __392950_392950;
   reg _392951_392951 ; 
   reg __392951_392951;
   reg _392952_392952 ; 
   reg __392952_392952;
   reg _392953_392953 ; 
   reg __392953_392953;
   reg _392954_392954 ; 
   reg __392954_392954;
   reg _392955_392955 ; 
   reg __392955_392955;
   reg _392956_392956 ; 
   reg __392956_392956;
   reg _392957_392957 ; 
   reg __392957_392957;
   reg _392958_392958 ; 
   reg __392958_392958;
   reg _392959_392959 ; 
   reg __392959_392959;
   reg _392960_392960 ; 
   reg __392960_392960;
   reg _392961_392961 ; 
   reg __392961_392961;
   reg _392962_392962 ; 
   reg __392962_392962;
   reg _392963_392963 ; 
   reg __392963_392963;
   reg _392964_392964 ; 
   reg __392964_392964;
   reg _392965_392965 ; 
   reg __392965_392965;
   reg _392966_392966 ; 
   reg __392966_392966;
   reg _392967_392967 ; 
   reg __392967_392967;
   reg _392968_392968 ; 
   reg __392968_392968;
   reg _392969_392969 ; 
   reg __392969_392969;
   reg _392970_392970 ; 
   reg __392970_392970;
   reg _392971_392971 ; 
   reg __392971_392971;
   reg _392972_392972 ; 
   reg __392972_392972;
   reg _392973_392973 ; 
   reg __392973_392973;
   reg _392974_392974 ; 
   reg __392974_392974;
   reg _392975_392975 ; 
   reg __392975_392975;
   reg _392976_392976 ; 
   reg __392976_392976;
   reg _392977_392977 ; 
   reg __392977_392977;
   reg _392978_392978 ; 
   reg __392978_392978;
   reg _392979_392979 ; 
   reg __392979_392979;
   reg _392980_392980 ; 
   reg __392980_392980;
   reg _392981_392981 ; 
   reg __392981_392981;
   reg _392982_392982 ; 
   reg __392982_392982;
   reg _392983_392983 ; 
   reg __392983_392983;
   reg _392984_392984 ; 
   reg __392984_392984;
   reg _392985_392985 ; 
   reg __392985_392985;
   reg _392986_392986 ; 
   reg __392986_392986;
   reg _392987_392987 ; 
   reg __392987_392987;
   reg _392988_392988 ; 
   reg __392988_392988;
   reg _392989_392989 ; 
   reg __392989_392989;
   reg _392990_392990 ; 
   reg __392990_392990;
   reg _392991_392991 ; 
   reg __392991_392991;
   reg _392992_392992 ; 
   reg __392992_392992;
   reg _392993_392993 ; 
   reg __392993_392993;
   reg _392994_392994 ; 
   reg __392994_392994;
   reg _392995_392995 ; 
   reg __392995_392995;
   reg _392996_392996 ; 
   reg __392996_392996;
   reg _392997_392997 ; 
   reg __392997_392997;
   reg _392998_392998 ; 
   reg __392998_392998;
   reg _392999_392999 ; 
   reg __392999_392999;
   reg _393000_393000 ; 
   reg __393000_393000;
   reg _393001_393001 ; 
   reg __393001_393001;
   reg _393002_393002 ; 
   reg __393002_393002;
   reg _393003_393003 ; 
   reg __393003_393003;
   reg _393004_393004 ; 
   reg __393004_393004;
   reg _393005_393005 ; 
   reg __393005_393005;
   reg _393006_393006 ; 
   reg __393006_393006;
   reg _393007_393007 ; 
   reg __393007_393007;
   reg _393008_393008 ; 
   reg __393008_393008;
   reg _393009_393009 ; 
   reg __393009_393009;
   reg _393010_393010 ; 
   reg __393010_393010;
   reg _393011_393011 ; 
   reg __393011_393011;
   reg _393012_393012 ; 
   reg __393012_393012;
   reg _393013_393013 ; 
   reg __393013_393013;
   reg _393014_393014 ; 
   reg __393014_393014;
   reg _393015_393015 ; 
   reg __393015_393015;
   reg _393016_393016 ; 
   reg __393016_393016;
   reg _393017_393017 ; 
   reg __393017_393017;
   reg _393018_393018 ; 
   reg __393018_393018;
   reg _393019_393019 ; 
   reg __393019_393019;
   reg _393020_393020 ; 
   reg __393020_393020;
   reg _393021_393021 ; 
   reg __393021_393021;
   reg _393022_393022 ; 
   reg __393022_393022;
   reg _393023_393023 ; 
   reg __393023_393023;
   reg _393024_393024 ; 
   reg __393024_393024;
   reg _393025_393025 ; 
   reg __393025_393025;
   reg _393026_393026 ; 
   reg __393026_393026;
   reg _393027_393027 ; 
   reg __393027_393027;
   reg _393028_393028 ; 
   reg __393028_393028;
   reg _393029_393029 ; 
   reg __393029_393029;
   reg _393030_393030 ; 
   reg __393030_393030;
   reg _393031_393031 ; 
   reg __393031_393031;
   reg _393032_393032 ; 
   reg __393032_393032;
   reg _393033_393033 ; 
   reg __393033_393033;
   reg _393034_393034 ; 
   reg __393034_393034;
   reg _393035_393035 ; 
   reg __393035_393035;
   reg _393036_393036 ; 
   reg __393036_393036;
   reg _393037_393037 ; 
   reg __393037_393037;
   reg _393038_393038 ; 
   reg __393038_393038;
   reg _393039_393039 ; 
   reg __393039_393039;
   reg _393040_393040 ; 
   reg __393040_393040;
   reg _393041_393041 ; 
   reg __393041_393041;
   reg _393042_393042 ; 
   reg __393042_393042;
   reg _393043_393043 ; 
   reg __393043_393043;
   reg _393044_393044 ; 
   reg __393044_393044;
   reg _393045_393045 ; 
   reg __393045_393045;
   reg _393046_393046 ; 
   reg __393046_393046;
   reg _393047_393047 ; 
   reg __393047_393047;
   reg _393048_393048 ; 
   reg __393048_393048;
   reg _393049_393049 ; 
   reg __393049_393049;
   reg _393050_393050 ; 
   reg __393050_393050;
   reg _393051_393051 ; 
   reg __393051_393051;
   reg _393052_393052 ; 
   reg __393052_393052;
   reg _393053_393053 ; 
   reg __393053_393053;
   reg _393054_393054 ; 
   reg __393054_393054;
   reg _393055_393055 ; 
   reg __393055_393055;
   reg _393056_393056 ; 
   reg __393056_393056;
   reg _393057_393057 ; 
   reg __393057_393057;
   reg _393058_393058 ; 
   reg __393058_393058;
   reg _393059_393059 ; 
   reg __393059_393059;
   reg _393060_393060 ; 
   reg __393060_393060;
   reg _393061_393061 ; 
   reg __393061_393061;
   reg _393062_393062 ; 
   reg __393062_393062;
   reg _393063_393063 ; 
   reg __393063_393063;
   reg _393064_393064 ; 
   reg __393064_393064;
   reg _393065_393065 ; 
   reg __393065_393065;
   reg _393066_393066 ; 
   reg __393066_393066;
   reg _393067_393067 ; 
   reg __393067_393067;
   reg _393068_393068 ; 
   reg __393068_393068;
   reg _393069_393069 ; 
   reg __393069_393069;
   reg _393070_393070 ; 
   reg __393070_393070;
   reg _393071_393071 ; 
   reg __393071_393071;
   reg _393072_393072 ; 
   reg __393072_393072;
   reg _393073_393073 ; 
   reg __393073_393073;
   reg _393074_393074 ; 
   reg __393074_393074;
   reg _393075_393075 ; 
   reg __393075_393075;
   reg _393076_393076 ; 
   reg __393076_393076;
   reg _393077_393077 ; 
   reg __393077_393077;
   reg _393078_393078 ; 
   reg __393078_393078;
   reg _393079_393079 ; 
   reg __393079_393079;
   reg _393080_393080 ; 
   reg __393080_393080;
   reg _393081_393081 ; 
   reg __393081_393081;
   reg _393082_393082 ; 
   reg __393082_393082;
   reg _393083_393083 ; 
   reg __393083_393083;
   reg _393084_393084 ; 
   reg __393084_393084;
   reg _393085_393085 ; 
   reg __393085_393085;
   reg _393086_393086 ; 
   reg __393086_393086;
   reg _393087_393087 ; 
   reg __393087_393087;
   reg _393088_393088 ; 
   reg __393088_393088;
   reg _393089_393089 ; 
   reg __393089_393089;
   reg _393090_393090 ; 
   reg __393090_393090;
   reg _393091_393091 ; 
   reg __393091_393091;
   reg _393092_393092 ; 
   reg __393092_393092;
   reg _393093_393093 ; 
   reg __393093_393093;
   reg _393094_393094 ; 
   reg __393094_393094;
   reg _393095_393095 ; 
   reg __393095_393095;
   reg _393096_393096 ; 
   reg __393096_393096;
   reg _393097_393097 ; 
   reg __393097_393097;
   reg _393098_393098 ; 
   reg __393098_393098;
   reg _393099_393099 ; 
   reg __393099_393099;
   reg _393100_393100 ; 
   reg __393100_393100;
   reg _393101_393101 ; 
   reg __393101_393101;
   reg _393102_393102 ; 
   reg __393102_393102;
   reg _393103_393103 ; 
   reg __393103_393103;
   reg _393104_393104 ; 
   reg __393104_393104;
   reg _393105_393105 ; 
   reg __393105_393105;
   reg _393106_393106 ; 
   reg __393106_393106;
   reg _393107_393107 ; 
   reg __393107_393107;
   reg _393108_393108 ; 
   reg __393108_393108;
   reg _393109_393109 ; 
   reg __393109_393109;
   reg _393110_393110 ; 
   reg __393110_393110;
   reg _393111_393111 ; 
   reg __393111_393111;
   reg _393112_393112 ; 
   reg __393112_393112;
   reg _393113_393113 ; 
   reg __393113_393113;
   reg _393114_393114 ; 
   reg __393114_393114;
   reg _393115_393115 ; 
   reg __393115_393115;
   reg _393116_393116 ; 
   reg __393116_393116;
   reg _393117_393117 ; 
   reg __393117_393117;
   reg _393118_393118 ; 
   reg __393118_393118;
   reg _393119_393119 ; 
   reg __393119_393119;
   reg _393120_393120 ; 
   reg __393120_393120;
   reg _393121_393121 ; 
   reg __393121_393121;
   reg _393122_393122 ; 
   reg __393122_393122;
   reg _393123_393123 ; 
   reg __393123_393123;
   reg _393124_393124 ; 
   reg __393124_393124;
   reg _393125_393125 ; 
   reg __393125_393125;
   reg _393126_393126 ; 
   reg __393126_393126;
   reg _393127_393127 ; 
   reg __393127_393127;
   reg _393128_393128 ; 
   reg __393128_393128;
   reg _393129_393129 ; 
   reg __393129_393129;
   reg _393130_393130 ; 
   reg __393130_393130;
   reg _393131_393131 ; 
   reg __393131_393131;
   reg _393132_393132 ; 
   reg __393132_393132;
   reg _393133_393133 ; 
   reg __393133_393133;
   reg _393134_393134 ; 
   reg __393134_393134;
   reg _393135_393135 ; 
   reg __393135_393135;
   reg _393136_393136 ; 
   reg __393136_393136;
   reg _393137_393137 ; 
   reg __393137_393137;
   reg _393138_393138 ; 
   reg __393138_393138;
   reg _393139_393139 ; 
   reg __393139_393139;
   reg _393140_393140 ; 
   reg __393140_393140;
   reg _393141_393141 ; 
   reg __393141_393141;
   reg _393142_393142 ; 
   reg __393142_393142;
   reg _393143_393143 ; 
   reg __393143_393143;
   reg _393144_393144 ; 
   reg __393144_393144;
   reg _393145_393145 ; 
   reg __393145_393145;
   reg _393146_393146 ; 
   reg __393146_393146;
   reg _393147_393147 ; 
   reg __393147_393147;
   reg _393148_393148 ; 
   reg __393148_393148;
   reg _393149_393149 ; 
   reg __393149_393149;
   reg _393150_393150 ; 
   reg __393150_393150;
   reg _393151_393151 ; 
   reg __393151_393151;
   reg _393152_393152 ; 
   reg __393152_393152;
   reg _393153_393153 ; 
   reg __393153_393153;
   reg _393154_393154 ; 
   reg __393154_393154;
   reg _393155_393155 ; 
   reg __393155_393155;
   reg _393156_393156 ; 
   reg __393156_393156;
   reg _393157_393157 ; 
   reg __393157_393157;
   reg _393158_393158 ; 
   reg __393158_393158;
   reg _393159_393159 ; 
   reg __393159_393159;
   reg _393160_393160 ; 
   reg __393160_393160;
   reg _393161_393161 ; 
   reg __393161_393161;
   reg _393162_393162 ; 
   reg __393162_393162;
   reg _393163_393163 ; 
   reg __393163_393163;
   reg _393164_393164 ; 
   reg __393164_393164;
   reg _393165_393165 ; 
   reg __393165_393165;
   reg _393166_393166 ; 
   reg __393166_393166;
   reg _393167_393167 ; 
   reg __393167_393167;
   reg _393168_393168 ; 
   reg __393168_393168;
   reg _393169_393169 ; 
   reg __393169_393169;
   reg _393170_393170 ; 
   reg __393170_393170;
   reg _393171_393171 ; 
   reg __393171_393171;
   reg _393172_393172 ; 
   reg __393172_393172;
   reg _393173_393173 ; 
   reg __393173_393173;
   reg _393174_393174 ; 
   reg __393174_393174;
   reg _393175_393175 ; 
   reg __393175_393175;
   reg _393176_393176 ; 
   reg __393176_393176;
   reg _393177_393177 ; 
   reg __393177_393177;
   reg _393178_393178 ; 
   reg __393178_393178;
   reg _393179_393179 ; 
   reg __393179_393179;
   reg _393180_393180 ; 
   reg __393180_393180;
   reg _393181_393181 ; 
   reg __393181_393181;
   reg _393182_393182 ; 
   reg __393182_393182;
   reg _393183_393183 ; 
   reg __393183_393183;
   reg _393184_393184 ; 
   reg __393184_393184;
   reg _393185_393185 ; 
   reg __393185_393185;
   reg _393186_393186 ; 
   reg __393186_393186;
   reg _393187_393187 ; 
   reg __393187_393187;
   reg _393188_393188 ; 
   reg __393188_393188;
   reg _393189_393189 ; 
   reg __393189_393189;
   reg _393190_393190 ; 
   reg __393190_393190;
   reg _393191_393191 ; 
   reg __393191_393191;
   reg _393192_393192 ; 
   reg __393192_393192;
   reg _393193_393193 ; 
   reg __393193_393193;
   reg _393194_393194 ; 
   reg __393194_393194;
   reg _393195_393195 ; 
   reg __393195_393195;
   reg _393196_393196 ; 
   reg __393196_393196;
   reg _393197_393197 ; 
   reg __393197_393197;
   reg _393198_393198 ; 
   reg __393198_393198;
   reg _393199_393199 ; 
   reg __393199_393199;
   reg _393200_393200 ; 
   reg __393200_393200;
   reg _393201_393201 ; 
   reg __393201_393201;
   reg _393202_393202 ; 
   reg __393202_393202;
   reg _393203_393203 ; 
   reg __393203_393203;
   reg _393204_393204 ; 
   reg __393204_393204;
   reg _393205_393205 ; 
   reg __393205_393205;
   reg _393206_393206 ; 
   reg __393206_393206;
   reg _393207_393207 ; 
   reg __393207_393207;
   reg _393208_393208 ; 
   reg __393208_393208;
   reg _393209_393209 ; 
   reg __393209_393209;
   reg _393210_393210 ; 
   reg __393210_393210;
   reg _393211_393211 ; 
   reg __393211_393211;
   reg _393212_393212 ; 
   reg __393212_393212;
   reg _393213_393213 ; 
   reg __393213_393213;
   reg _393214_393214 ; 
   reg __393214_393214;
   reg _393215_393215 ; 
   reg __393215_393215;
   reg _393216_393216 ; 
   reg __393216_393216;
   reg _393217_393217 ; 
   reg __393217_393217;
   reg _393218_393218 ; 
   reg __393218_393218;
   reg _393219_393219 ; 
   reg __393219_393219;
   reg _393220_393220 ; 
   reg __393220_393220;
   reg _393221_393221 ; 
   reg __393221_393221;
   reg _393222_393222 ; 
   reg __393222_393222;
   reg _393223_393223 ; 
   reg __393223_393223;
   reg _393224_393224 ; 
   reg __393224_393224;
   reg _393225_393225 ; 
   reg __393225_393225;
   reg _393226_393226 ; 
   reg __393226_393226;
   reg _393227_393227 ; 
   reg __393227_393227;
   reg _393228_393228 ; 
   reg __393228_393228;
   reg _393229_393229 ; 
   reg __393229_393229;
   reg _393230_393230 ; 
   reg __393230_393230;
   reg _393231_393231 ; 
   reg __393231_393231;
   reg _393232_393232 ; 
   reg __393232_393232;
   reg _393233_393233 ; 
   reg __393233_393233;
   reg _393234_393234 ; 
   reg __393234_393234;
   reg _393235_393235 ; 
   reg __393235_393235;
   reg _393236_393236 ; 
   reg __393236_393236;
   reg _393237_393237 ; 
   reg __393237_393237;
   reg _393238_393238 ; 
   reg __393238_393238;
   reg _393239_393239 ; 
   reg __393239_393239;
   reg _393240_393240 ; 
   reg __393240_393240;
   reg _393241_393241 ; 
   reg __393241_393241;
   reg _393242_393242 ; 
   reg __393242_393242;
   reg _393243_393243 ; 
   reg __393243_393243;
   reg _393244_393244 ; 
   reg __393244_393244;
   reg _393245_393245 ; 
   reg __393245_393245;
   reg _393246_393246 ; 
   reg __393246_393246;
   reg _393247_393247 ; 
   reg __393247_393247;
   reg _393248_393248 ; 
   reg __393248_393248;
   reg _393249_393249 ; 
   reg __393249_393249;
   reg _393250_393250 ; 
   reg __393250_393250;
   reg _393251_393251 ; 
   reg __393251_393251;
   reg _393252_393252 ; 
   reg __393252_393252;
   reg _393253_393253 ; 
   reg __393253_393253;
   reg _393254_393254 ; 
   reg __393254_393254;
   reg _393255_393255 ; 
   reg __393255_393255;
   reg _393256_393256 ; 
   reg __393256_393256;
   reg _393257_393257 ; 
   reg __393257_393257;
   reg _393258_393258 ; 
   reg __393258_393258;
   reg _393259_393259 ; 
   reg __393259_393259;
   reg _393260_393260 ; 
   reg __393260_393260;
   reg _393261_393261 ; 
   reg __393261_393261;
   reg _393262_393262 ; 
   reg __393262_393262;
   reg _393263_393263 ; 
   reg __393263_393263;
   reg _393264_393264 ; 
   reg __393264_393264;
   reg _393265_393265 ; 
   reg __393265_393265;
   reg _393266_393266 ; 
   reg __393266_393266;
   reg _393267_393267 ; 
   reg __393267_393267;
   reg _393268_393268 ; 
   reg __393268_393268;
   reg _393269_393269 ; 
   reg __393269_393269;
   reg _393270_393270 ; 
   reg __393270_393270;
   reg _393271_393271 ; 
   reg __393271_393271;
   reg _393272_393272 ; 
   reg __393272_393272;
   reg _393273_393273 ; 
   reg __393273_393273;
   reg _393274_393274 ; 
   reg __393274_393274;
   reg _393275_393275 ; 
   reg __393275_393275;
   reg _393276_393276 ; 
   reg __393276_393276;
   reg _393277_393277 ; 
   reg __393277_393277;
   reg _393278_393278 ; 
   reg __393278_393278;
   reg _393279_393279 ; 
   reg __393279_393279;
   reg _393280_393280 ; 
   reg __393280_393280;
   reg _393281_393281 ; 
   reg __393281_393281;
   reg _393282_393282 ; 
   reg __393282_393282;
   reg _393283_393283 ; 
   reg __393283_393283;
   reg _393284_393284 ; 
   reg __393284_393284;
   reg _393285_393285 ; 
   reg __393285_393285;
   reg _393286_393286 ; 
   reg __393286_393286;
   reg _393287_393287 ; 
   reg __393287_393287;
   reg _393288_393288 ; 
   reg __393288_393288;
   reg _393289_393289 ; 
   reg __393289_393289;
   reg _393290_393290 ; 
   reg __393290_393290;
   reg _393291_393291 ; 
   reg __393291_393291;
   reg _393292_393292 ; 
   reg __393292_393292;
   reg _393293_393293 ; 
   reg __393293_393293;
   reg _393294_393294 ; 
   reg __393294_393294;
   reg _393295_393295 ; 
   reg __393295_393295;
   reg _393296_393296 ; 
   reg __393296_393296;
   reg _393297_393297 ; 
   reg __393297_393297;
   reg _393298_393298 ; 
   reg __393298_393298;
   reg _393299_393299 ; 
   reg __393299_393299;
   reg _393300_393300 ; 
   reg __393300_393300;
   reg _393301_393301 ; 
   reg __393301_393301;
   reg _393302_393302 ; 
   reg __393302_393302;
   reg _393303_393303 ; 
   reg __393303_393303;
   reg _393304_393304 ; 
   reg __393304_393304;
   reg _393305_393305 ; 
   reg __393305_393305;
   reg _393306_393306 ; 
   reg __393306_393306;
   reg _393307_393307 ; 
   reg __393307_393307;
   reg _393308_393308 ; 
   reg __393308_393308;
   reg _393309_393309 ; 
   reg __393309_393309;
   reg _393310_393310 ; 
   reg __393310_393310;
   reg _393311_393311 ; 
   reg __393311_393311;
   reg _393312_393312 ; 
   reg __393312_393312;
   reg _393313_393313 ; 
   reg __393313_393313;
   reg _393314_393314 ; 
   reg __393314_393314;
   reg _393315_393315 ; 
   reg __393315_393315;
   reg _393316_393316 ; 
   reg __393316_393316;
   reg _393317_393317 ; 
   reg __393317_393317;
   reg _393318_393318 ; 
   reg __393318_393318;
   reg _393319_393319 ; 
   reg __393319_393319;
   reg _393320_393320 ; 
   reg __393320_393320;
   reg _393321_393321 ; 
   reg __393321_393321;
   reg _393322_393322 ; 
   reg __393322_393322;
   reg _393323_393323 ; 
   reg __393323_393323;
   reg _393324_393324 ; 
   reg __393324_393324;
   reg _393325_393325 ; 
   reg __393325_393325;
   reg _393326_393326 ; 
   reg __393326_393326;
   reg _393327_393327 ; 
   reg __393327_393327;
   reg _393328_393328 ; 
   reg __393328_393328;
   reg _393329_393329 ; 
   reg __393329_393329;
   reg _393330_393330 ; 
   reg __393330_393330;
   reg _393331_393331 ; 
   reg __393331_393331;
   reg _393332_393332 ; 
   reg __393332_393332;
   reg _393333_393333 ; 
   reg __393333_393333;
   reg _393334_393334 ; 
   reg __393334_393334;
   reg _393335_393335 ; 
   reg __393335_393335;
   reg _393336_393336 ; 
   reg __393336_393336;
   reg _393337_393337 ; 
   reg __393337_393337;
   reg _393338_393338 ; 
   reg __393338_393338;
   reg _393339_393339 ; 
   reg __393339_393339;
   reg _393340_393340 ; 
   reg __393340_393340;
   reg _393341_393341 ; 
   reg __393341_393341;
   reg _393342_393342 ; 
   reg __393342_393342;
   reg _393343_393343 ; 
   reg __393343_393343;
   reg _393344_393344 ; 
   reg __393344_393344;
   reg _393345_393345 ; 
   reg __393345_393345;
   reg _393346_393346 ; 
   reg __393346_393346;
   reg _393347_393347 ; 
   reg __393347_393347;
   reg _393348_393348 ; 
   reg __393348_393348;
   reg _393349_393349 ; 
   reg __393349_393349;
   reg _393350_393350 ; 
   reg __393350_393350;
   reg _393351_393351 ; 
   reg __393351_393351;
   reg _393352_393352 ; 
   reg __393352_393352;
   reg _393353_393353 ; 
   reg __393353_393353;
   reg _393354_393354 ; 
   reg __393354_393354;
   reg _393355_393355 ; 
   reg __393355_393355;
   reg _393356_393356 ; 
   reg __393356_393356;
   reg _393357_393357 ; 
   reg __393357_393357;
   reg _393358_393358 ; 
   reg __393358_393358;
   reg _393359_393359 ; 
   reg __393359_393359;
   reg _393360_393360 ; 
   reg __393360_393360;
   reg _393361_393361 ; 
   reg __393361_393361;
   reg _393362_393362 ; 
   reg __393362_393362;
   reg _393363_393363 ; 
   reg __393363_393363;
   reg _393364_393364 ; 
   reg __393364_393364;
   reg _393365_393365 ; 
   reg __393365_393365;
   reg _393366_393366 ; 
   reg __393366_393366;
   reg _393367_393367 ; 
   reg __393367_393367;
   reg _393368_393368 ; 
   reg __393368_393368;
   reg _393369_393369 ; 
   reg __393369_393369;
   reg _393370_393370 ; 
   reg __393370_393370;
   reg _393371_393371 ; 
   reg __393371_393371;
   reg _393372_393372 ; 
   reg __393372_393372;
   reg _393373_393373 ; 
   reg __393373_393373;
   reg _393374_393374 ; 
   reg __393374_393374;
   reg _393375_393375 ; 
   reg __393375_393375;
   reg _393376_393376 ; 
   reg __393376_393376;
   reg _393377_393377 ; 
   reg __393377_393377;
   reg _393378_393378 ; 
   reg __393378_393378;
   reg _393379_393379 ; 
   reg __393379_393379;
   reg _393380_393380 ; 
   reg __393380_393380;
   reg _393381_393381 ; 
   reg __393381_393381;
   reg _393382_393382 ; 
   reg __393382_393382;
   reg _393383_393383 ; 
   reg __393383_393383;
   reg _393384_393384 ; 
   reg __393384_393384;
   reg _393385_393385 ; 
   reg __393385_393385;
   reg _393386_393386 ; 
   reg __393386_393386;
   reg _393387_393387 ; 
   reg __393387_393387;
   reg _393388_393388 ; 
   reg __393388_393388;
   reg _393389_393389 ; 
   reg __393389_393389;
   reg _393390_393390 ; 
   reg __393390_393390;
   reg _393391_393391 ; 
   reg __393391_393391;
   reg _393392_393392 ; 
   reg __393392_393392;
   reg _393393_393393 ; 
   reg __393393_393393;
   reg _393394_393394 ; 
   reg __393394_393394;
   reg _393395_393395 ; 
   reg __393395_393395;
   reg _393396_393396 ; 
   reg __393396_393396;
   reg _393397_393397 ; 
   reg __393397_393397;
   reg _393398_393398 ; 
   reg __393398_393398;
   reg _393399_393399 ; 
   reg __393399_393399;
   reg _393400_393400 ; 
   reg __393400_393400;
   reg _393401_393401 ; 
   reg __393401_393401;
   reg _393402_393402 ; 
   reg __393402_393402;
   reg _393403_393403 ; 
   reg __393403_393403;
   reg _393404_393404 ; 
   reg __393404_393404;
   reg _393405_393405 ; 
   reg __393405_393405;
   reg _393406_393406 ; 
   reg __393406_393406;
   reg _393407_393407 ; 
   reg __393407_393407;
   reg _393408_393408 ; 
   reg __393408_393408;
   reg _393409_393409 ; 
   reg __393409_393409;
   reg _393410_393410 ; 
   reg __393410_393410;
   reg _393411_393411 ; 
   reg __393411_393411;
   reg _393412_393412 ; 
   reg __393412_393412;
   reg _393413_393413 ; 
   reg __393413_393413;
   reg _393414_393414 ; 
   reg __393414_393414;
   reg _393415_393415 ; 
   reg __393415_393415;
   reg _393416_393416 ; 
   reg __393416_393416;
   reg _393417_393417 ; 
   reg __393417_393417;
   reg _393418_393418 ; 
   reg __393418_393418;
   reg _393419_393419 ; 
   reg __393419_393419;
   reg _393420_393420 ; 
   reg __393420_393420;
   reg _393421_393421 ; 
   reg __393421_393421;
   reg _393422_393422 ; 
   reg __393422_393422;
   reg _393423_393423 ; 
   reg __393423_393423;
   reg _393424_393424 ; 
   reg __393424_393424;
   reg _393425_393425 ; 
   reg __393425_393425;
   reg _393426_393426 ; 
   reg __393426_393426;
   reg _393427_393427 ; 
   reg __393427_393427;
   reg _393428_393428 ; 
   reg __393428_393428;
   reg _393429_393429 ; 
   reg __393429_393429;
   reg _393430_393430 ; 
   reg __393430_393430;
   reg _393431_393431 ; 
   reg __393431_393431;
   reg _393432_393432 ; 
   reg __393432_393432;
   reg _393433_393433 ; 
   reg __393433_393433;
   reg _393434_393434 ; 
   reg __393434_393434;
   reg _393435_393435 ; 
   reg __393435_393435;
   reg _393436_393436 ; 
   reg __393436_393436;
   reg _393437_393437 ; 
   reg __393437_393437;
   reg _393438_393438 ; 
   reg __393438_393438;
   reg _393439_393439 ; 
   reg __393439_393439;
   reg _393440_393440 ; 
   reg __393440_393440;
   reg _393441_393441 ; 
   reg __393441_393441;
   reg _393442_393442 ; 
   reg __393442_393442;
   reg _393443_393443 ; 
   reg __393443_393443;
   reg _393444_393444 ; 
   reg __393444_393444;
   reg _393445_393445 ; 
   reg __393445_393445;
   reg _393446_393446 ; 
   reg __393446_393446;
   reg _393447_393447 ; 
   reg __393447_393447;
   reg _393448_393448 ; 
   reg __393448_393448;
   reg _393449_393449 ; 
   reg __393449_393449;
   reg _393450_393450 ; 
   reg __393450_393450;
   reg _393451_393451 ; 
   reg __393451_393451;
   reg _393452_393452 ; 
   reg __393452_393452;
   reg _393453_393453 ; 
   reg __393453_393453;
   reg _393454_393454 ; 
   reg __393454_393454;
   reg _393455_393455 ; 
   reg __393455_393455;
   reg _393456_393456 ; 
   reg __393456_393456;
   reg _393457_393457 ; 
   reg __393457_393457;
   reg _393458_393458 ; 
   reg __393458_393458;
   reg _393459_393459 ; 
   reg __393459_393459;
   reg _393460_393460 ; 
   reg __393460_393460;
   reg _393461_393461 ; 
   reg __393461_393461;
   reg _393462_393462 ; 
   reg __393462_393462;
   reg _393463_393463 ; 
   reg __393463_393463;
   reg _393464_393464 ; 
   reg __393464_393464;
   reg _393465_393465 ; 
   reg __393465_393465;
   reg _393466_393466 ; 
   reg __393466_393466;
   reg _393467_393467 ; 
   reg __393467_393467;
   reg _393468_393468 ; 
   reg __393468_393468;
   reg _393469_393469 ; 
   reg __393469_393469;
   reg _393470_393470 ; 
   reg __393470_393470;
   reg _393471_393471 ; 
   reg __393471_393471;
   reg _393472_393472 ; 
   reg __393472_393472;
   reg _393473_393473 ; 
   reg __393473_393473;
   reg _393474_393474 ; 
   reg __393474_393474;
   reg _393475_393475 ; 
   reg __393475_393475;
   reg _393476_393476 ; 
   reg __393476_393476;
   reg _393477_393477 ; 
   reg __393477_393477;
   reg _393478_393478 ; 
   reg __393478_393478;
   reg _393479_393479 ; 
   reg __393479_393479;
   reg _393480_393480 ; 
   reg __393480_393480;
   reg _393481_393481 ; 
   reg __393481_393481;
   reg _393482_393482 ; 
   reg __393482_393482;
   reg _393483_393483 ; 
   reg __393483_393483;
   reg _393484_393484 ; 
   reg __393484_393484;
   reg _393485_393485 ; 
   reg __393485_393485;
   reg _393486_393486 ; 
   reg __393486_393486;
   reg _393487_393487 ; 
   reg __393487_393487;
   reg _393488_393488 ; 
   reg __393488_393488;
   reg _393489_393489 ; 
   reg __393489_393489;
   reg _393490_393490 ; 
   reg __393490_393490;
   reg _393491_393491 ; 
   reg __393491_393491;
   reg _393492_393492 ; 
   reg __393492_393492;
   reg _393493_393493 ; 
   reg __393493_393493;
   reg _393494_393494 ; 
   reg __393494_393494;
   reg _393495_393495 ; 
   reg __393495_393495;
   reg _393496_393496 ; 
   reg __393496_393496;
   reg _393497_393497 ; 
   reg __393497_393497;
   reg _393498_393498 ; 
   reg __393498_393498;
   reg _393499_393499 ; 
   reg __393499_393499;
   reg _393500_393500 ; 
   reg __393500_393500;
   reg _393501_393501 ; 
   reg __393501_393501;
   reg _393502_393502 ; 
   reg __393502_393502;
   reg _393503_393503 ; 
   reg __393503_393503;
   reg _393504_393504 ; 
   reg __393504_393504;
   reg _393505_393505 ; 
   reg __393505_393505;
   reg _393506_393506 ; 
   reg __393506_393506;
   reg _393507_393507 ; 
   reg __393507_393507;
   reg _393508_393508 ; 
   reg __393508_393508;
   reg _393509_393509 ; 
   reg __393509_393509;
   reg _393510_393510 ; 
   reg __393510_393510;
   reg _393511_393511 ; 
   reg __393511_393511;
   reg _393512_393512 ; 
   reg __393512_393512;
   reg _393513_393513 ; 
   reg __393513_393513;
   reg _393514_393514 ; 
   reg __393514_393514;
   reg _393515_393515 ; 
   reg __393515_393515;
   reg _393516_393516 ; 
   reg __393516_393516;
   reg _393517_393517 ; 
   reg __393517_393517;
   reg _393518_393518 ; 
   reg __393518_393518;
   reg _393519_393519 ; 
   reg __393519_393519;
   reg _393520_393520 ; 
   reg __393520_393520;
   reg _393521_393521 ; 
   reg __393521_393521;
   reg _393522_393522 ; 
   reg __393522_393522;
   reg _393523_393523 ; 
   reg __393523_393523;
   reg _393524_393524 ; 
   reg __393524_393524;
   reg _393525_393525 ; 
   reg __393525_393525;
   reg _393526_393526 ; 
   reg __393526_393526;
   reg _393527_393527 ; 
   reg __393527_393527;
   reg _393528_393528 ; 
   reg __393528_393528;
   reg _393529_393529 ; 
   reg __393529_393529;
   reg _393530_393530 ; 
   reg __393530_393530;
   reg _393531_393531 ; 
   reg __393531_393531;
   reg _393532_393532 ; 
   reg __393532_393532;
   reg _393533_393533 ; 
   reg __393533_393533;
   reg _393534_393534 ; 
   reg __393534_393534;
   reg _393535_393535 ; 
   reg __393535_393535;
   reg _393536_393536 ; 
   reg __393536_393536;
   reg _393537_393537 ; 
   reg __393537_393537;
   reg _393538_393538 ; 
   reg __393538_393538;
   reg _393539_393539 ; 
   reg __393539_393539;
   reg _393540_393540 ; 
   reg __393540_393540;
   reg _393541_393541 ; 
   reg __393541_393541;
   reg _393542_393542 ; 
   reg __393542_393542;
   reg _393543_393543 ; 
   reg __393543_393543;
   reg _393544_393544 ; 
   reg __393544_393544;
   reg _393545_393545 ; 
   reg __393545_393545;
   reg _393546_393546 ; 
   reg __393546_393546;
   reg _393547_393547 ; 
   reg __393547_393547;
   reg _393548_393548 ; 
   reg __393548_393548;
   reg _393549_393549 ; 
   reg __393549_393549;
   reg _393550_393550 ; 
   reg __393550_393550;
   reg _393551_393551 ; 
   reg __393551_393551;
   reg _393552_393552 ; 
   reg __393552_393552;
   reg _393553_393553 ; 
   reg __393553_393553;
   reg _393554_393554 ; 
   reg __393554_393554;
   reg _393555_393555 ; 
   reg __393555_393555;
   reg _393556_393556 ; 
   reg __393556_393556;
   reg _393557_393557 ; 
   reg __393557_393557;
   reg _393558_393558 ; 
   reg __393558_393558;
   reg _393559_393559 ; 
   reg __393559_393559;
   reg _393560_393560 ; 
   reg __393560_393560;
   reg _393561_393561 ; 
   reg __393561_393561;
   reg _393562_393562 ; 
   reg __393562_393562;
   reg _393563_393563 ; 
   reg __393563_393563;
   reg _393564_393564 ; 
   reg __393564_393564;
   reg _393565_393565 ; 
   reg __393565_393565;
   reg _393566_393566 ; 
   reg __393566_393566;
   reg _393567_393567 ; 
   reg __393567_393567;
   reg _393568_393568 ; 
   reg __393568_393568;
   reg _393569_393569 ; 
   reg __393569_393569;
   reg _393570_393570 ; 
   reg __393570_393570;
   reg _393571_393571 ; 
   reg __393571_393571;
   reg _393572_393572 ; 
   reg __393572_393572;
   reg _393573_393573 ; 
   reg __393573_393573;
   reg _393574_393574 ; 
   reg __393574_393574;
   reg _393575_393575 ; 
   reg __393575_393575;
   reg _393576_393576 ; 
   reg __393576_393576;
   reg _393577_393577 ; 
   reg __393577_393577;
   reg _393578_393578 ; 
   reg __393578_393578;
   reg _393579_393579 ; 
   reg __393579_393579;
   reg _393580_393580 ; 
   reg __393580_393580;
   reg _393581_393581 ; 
   reg __393581_393581;
   reg _393582_393582 ; 
   reg __393582_393582;
   reg _393583_393583 ; 
   reg __393583_393583;
   reg _393584_393584 ; 
   reg __393584_393584;
   reg _393585_393585 ; 
   reg __393585_393585;
   reg _393586_393586 ; 
   reg __393586_393586;
   reg _393587_393587 ; 
   reg __393587_393587;
   reg _393588_393588 ; 
   reg __393588_393588;
   reg _393589_393589 ; 
   reg __393589_393589;
   reg _393590_393590 ; 
   reg __393590_393590;
   reg _393591_393591 ; 
   reg __393591_393591;
   reg _393592_393592 ; 
   reg __393592_393592;
   reg _393593_393593 ; 
   reg __393593_393593;
   reg _393594_393594 ; 
   reg __393594_393594;
   reg _393595_393595 ; 
   reg __393595_393595;
   reg _393596_393596 ; 
   reg __393596_393596;
   reg _393597_393597 ; 
   reg __393597_393597;
   reg _393598_393598 ; 
   reg __393598_393598;
   reg _393599_393599 ; 
   reg __393599_393599;
   reg _393600_393600 ; 
   reg __393600_393600;
   reg _393601_393601 ; 
   reg __393601_393601;
   reg _393602_393602 ; 
   reg __393602_393602;
   reg _393603_393603 ; 
   reg __393603_393603;
   reg _393604_393604 ; 
   reg __393604_393604;
   reg _393605_393605 ; 
   reg __393605_393605;
   reg _393606_393606 ; 
   reg __393606_393606;
   reg _393607_393607 ; 
   reg __393607_393607;
   reg _393608_393608 ; 
   reg __393608_393608;
   reg _393609_393609 ; 
   reg __393609_393609;
   reg _393610_393610 ; 
   reg __393610_393610;
   reg _393611_393611 ; 
   reg __393611_393611;
   reg _393612_393612 ; 
   reg __393612_393612;
   reg _393613_393613 ; 
   reg __393613_393613;
   reg _393614_393614 ; 
   reg __393614_393614;
   reg _393615_393615 ; 
   reg __393615_393615;
   reg _393616_393616 ; 
   reg __393616_393616;
   reg _393617_393617 ; 
   reg __393617_393617;
   reg _393618_393618 ; 
   reg __393618_393618;
   reg _393619_393619 ; 
   reg __393619_393619;
   reg _393620_393620 ; 
   reg __393620_393620;
   reg _393621_393621 ; 
   reg __393621_393621;
   reg _393622_393622 ; 
   reg __393622_393622;
   reg _393623_393623 ; 
   reg __393623_393623;
   reg _393624_393624 ; 
   reg __393624_393624;
   reg _393625_393625 ; 
   reg __393625_393625;
   reg _393626_393626 ; 
   reg __393626_393626;
   reg _393627_393627 ; 
   reg __393627_393627;
   reg _393628_393628 ; 
   reg __393628_393628;
   reg _393629_393629 ; 
   reg __393629_393629;
   reg _393630_393630 ; 
   reg __393630_393630;
   reg _393631_393631 ; 
   reg __393631_393631;
   reg _393632_393632 ; 
   reg __393632_393632;
   reg _393633_393633 ; 
   reg __393633_393633;
   reg _393634_393634 ; 
   reg __393634_393634;
   reg _393635_393635 ; 
   reg __393635_393635;
   reg _393636_393636 ; 
   reg __393636_393636;
   reg _393637_393637 ; 
   reg __393637_393637;
   reg _393638_393638 ; 
   reg __393638_393638;
   reg _393639_393639 ; 
   reg __393639_393639;
   reg _393640_393640 ; 
   reg __393640_393640;
   reg _393641_393641 ; 
   reg __393641_393641;
   reg _393642_393642 ; 
   reg __393642_393642;
   reg _393643_393643 ; 
   reg __393643_393643;
   reg _393644_393644 ; 
   reg __393644_393644;
   reg _393645_393645 ; 
   reg __393645_393645;
   reg _393646_393646 ; 
   reg __393646_393646;
   reg _393647_393647 ; 
   reg __393647_393647;
   reg _393648_393648 ; 
   reg __393648_393648;
   reg _393649_393649 ; 
   reg __393649_393649;
   reg _393650_393650 ; 
   reg __393650_393650;
   reg _393651_393651 ; 
   reg __393651_393651;
   reg _393652_393652 ; 
   reg __393652_393652;
   reg _393653_393653 ; 
   reg __393653_393653;
   reg _393654_393654 ; 
   reg __393654_393654;
   reg _393655_393655 ; 
   reg __393655_393655;
   reg _393656_393656 ; 
   reg __393656_393656;
   reg _393657_393657 ; 
   reg __393657_393657;
   reg _393658_393658 ; 
   reg __393658_393658;
   reg _393659_393659 ; 
   reg __393659_393659;
   reg _393660_393660 ; 
   reg __393660_393660;
   reg _393661_393661 ; 
   reg __393661_393661;
   reg _393662_393662 ; 
   reg __393662_393662;
   reg _393663_393663 ; 
   reg __393663_393663;
   reg _393664_393664 ; 
   reg __393664_393664;
   reg _393665_393665 ; 
   reg __393665_393665;
   reg _393666_393666 ; 
   reg __393666_393666;
   reg _393667_393667 ; 
   reg __393667_393667;
   reg _393668_393668 ; 
   reg __393668_393668;
   reg _393669_393669 ; 
   reg __393669_393669;
   reg _393670_393670 ; 
   reg __393670_393670;
   reg _393671_393671 ; 
   reg __393671_393671;
   reg _393672_393672 ; 
   reg __393672_393672;
   reg _393673_393673 ; 
   reg __393673_393673;
   reg _393674_393674 ; 
   reg __393674_393674;
   reg _393675_393675 ; 
   reg __393675_393675;
   reg _393676_393676 ; 
   reg __393676_393676;
   reg _393677_393677 ; 
   reg __393677_393677;
   reg _393678_393678 ; 
   reg __393678_393678;
   reg _393679_393679 ; 
   reg __393679_393679;
   reg _393680_393680 ; 
   reg __393680_393680;
   reg _393681_393681 ; 
   reg __393681_393681;
   reg _393682_393682 ; 
   reg __393682_393682;
   reg _393683_393683 ; 
   reg __393683_393683;
   reg _393684_393684 ; 
   reg __393684_393684;
   reg _393685_393685 ; 
   reg __393685_393685;
   reg _393686_393686 ; 
   reg __393686_393686;
   reg _393687_393687 ; 
   reg __393687_393687;
   reg _393688_393688 ; 
   reg __393688_393688;
   reg _393689_393689 ; 
   reg __393689_393689;
   reg _393690_393690 ; 
   reg __393690_393690;
   reg _393691_393691 ; 
   reg __393691_393691;
   reg _393692_393692 ; 
   reg __393692_393692;
   reg _393693_393693 ; 
   reg __393693_393693;
   reg _393694_393694 ; 
   reg __393694_393694;
   reg _393695_393695 ; 
   reg __393695_393695;
   reg _393696_393696 ; 
   reg __393696_393696;
   reg _393697_393697 ; 
   reg __393697_393697;
   reg _393698_393698 ; 
   reg __393698_393698;
   reg _393699_393699 ; 
   reg __393699_393699;
   reg _393700_393700 ; 
   reg __393700_393700;
   reg _393701_393701 ; 
   reg __393701_393701;
   reg _393702_393702 ; 
   reg __393702_393702;
   reg _393703_393703 ; 
   reg __393703_393703;
   reg _393704_393704 ; 
   reg __393704_393704;
   reg _393705_393705 ; 
   reg __393705_393705;
   reg _393706_393706 ; 
   reg __393706_393706;
   reg _393707_393707 ; 
   reg __393707_393707;
   reg _393708_393708 ; 
   reg __393708_393708;
   reg _393709_393709 ; 
   reg __393709_393709;
   reg _393710_393710 ; 
   reg __393710_393710;
   reg _393711_393711 ; 
   reg __393711_393711;
   reg _393712_393712 ; 
   reg __393712_393712;
   reg _393713_393713 ; 
   reg __393713_393713;
   reg _393714_393714 ; 
   reg __393714_393714;
   reg _393715_393715 ; 
   reg __393715_393715;
   reg _393716_393716 ; 
   reg __393716_393716;
   reg _393717_393717 ; 
   reg __393717_393717;
   reg _393718_393718 ; 
   reg __393718_393718;
   reg _393719_393719 ; 
   reg __393719_393719;
   reg _393720_393720 ; 
   reg __393720_393720;
   reg _393721_393721 ; 
   reg __393721_393721;
   reg _393722_393722 ; 
   reg __393722_393722;
   reg _393723_393723 ; 
   reg __393723_393723;
   reg _393724_393724 ; 
   reg __393724_393724;
   reg _393725_393725 ; 
   reg __393725_393725;
   reg _393726_393726 ; 
   reg __393726_393726;
   reg _393727_393727 ; 
   reg __393727_393727;
   reg _393728_393728 ; 
   reg __393728_393728;
   reg _393729_393729 ; 
   reg __393729_393729;
   reg _393730_393730 ; 
   reg __393730_393730;
   reg _393731_393731 ; 
   reg __393731_393731;
   reg _393732_393732 ; 
   reg __393732_393732;
   reg _393733_393733 ; 
   reg __393733_393733;
   reg _393734_393734 ; 
   reg __393734_393734;
   reg _393735_393735 ; 
   reg __393735_393735;
   reg _393736_393736 ; 
   reg __393736_393736;
   reg _393737_393737 ; 
   reg __393737_393737;
   reg _393738_393738 ; 
   reg __393738_393738;
   reg _393739_393739 ; 
   reg __393739_393739;
   reg _393740_393740 ; 
   reg __393740_393740;
   reg _393741_393741 ; 
   reg __393741_393741;
   reg _393742_393742 ; 
   reg __393742_393742;
   reg _393743_393743 ; 
   reg __393743_393743;
   reg _393744_393744 ; 
   reg __393744_393744;
   reg _393745_393745 ; 
   reg __393745_393745;
   reg _393746_393746 ; 
   reg __393746_393746;
   reg _393747_393747 ; 
   reg __393747_393747;
   reg _393748_393748 ; 
   reg __393748_393748;
   reg _393749_393749 ; 
   reg __393749_393749;
   reg _393750_393750 ; 
   reg __393750_393750;
   reg _393751_393751 ; 
   reg __393751_393751;
   reg _393752_393752 ; 
   reg __393752_393752;
   reg _393753_393753 ; 
   reg __393753_393753;
   reg _393754_393754 ; 
   reg __393754_393754;
   reg _393755_393755 ; 
   reg __393755_393755;
   reg _393756_393756 ; 
   reg __393756_393756;
   reg _393757_393757 ; 
   reg __393757_393757;
   reg _393758_393758 ; 
   reg __393758_393758;
   reg _393759_393759 ; 
   reg __393759_393759;
   reg _393760_393760 ; 
   reg __393760_393760;
   reg _393761_393761 ; 
   reg __393761_393761;
   reg _393762_393762 ; 
   reg __393762_393762;
   reg _393763_393763 ; 
   reg __393763_393763;
   reg _393764_393764 ; 
   reg __393764_393764;
   reg _393765_393765 ; 
   reg __393765_393765;
   reg _393766_393766 ; 
   reg __393766_393766;
   reg _393767_393767 ; 
   reg __393767_393767;
   reg _393768_393768 ; 
   reg __393768_393768;
   reg _393769_393769 ; 
   reg __393769_393769;
   reg _393770_393770 ; 
   reg __393770_393770;
   reg _393771_393771 ; 
   reg __393771_393771;
   reg _393772_393772 ; 
   reg __393772_393772;
   reg _393773_393773 ; 
   reg __393773_393773;
   reg _393774_393774 ; 
   reg __393774_393774;
   reg _393775_393775 ; 
   reg __393775_393775;
   reg _393776_393776 ; 
   reg __393776_393776;
   reg _393777_393777 ; 
   reg __393777_393777;
   reg _393778_393778 ; 
   reg __393778_393778;
   reg _393779_393779 ; 
   reg __393779_393779;
   reg _393780_393780 ; 
   reg __393780_393780;
   reg _393781_393781 ; 
   reg __393781_393781;
   reg _393782_393782 ; 
   reg __393782_393782;
   reg _393783_393783 ; 
   reg __393783_393783;
   reg _393784_393784 ; 
   reg __393784_393784;
   reg _393785_393785 ; 
   reg __393785_393785;
   reg _393786_393786 ; 
   reg __393786_393786;
   reg _393787_393787 ; 
   reg __393787_393787;
   reg _393788_393788 ; 
   reg __393788_393788;
   reg _393789_393789 ; 
   reg __393789_393789;
   reg _393790_393790 ; 
   reg __393790_393790;
   reg _393791_393791 ; 
   reg __393791_393791;
   reg _393792_393792 ; 
   reg __393792_393792;
   reg _393793_393793 ; 
   reg __393793_393793;
   reg _393794_393794 ; 
   reg __393794_393794;
   reg _393795_393795 ; 
   reg __393795_393795;
   reg _393796_393796 ; 
   reg __393796_393796;
   reg _393797_393797 ; 
   reg __393797_393797;
   reg _393798_393798 ; 
   reg __393798_393798;
   reg _393799_393799 ; 
   reg __393799_393799;
   reg _393800_393800 ; 
   reg __393800_393800;
   reg _393801_393801 ; 
   reg __393801_393801;
   reg _393802_393802 ; 
   reg __393802_393802;
   reg _393803_393803 ; 
   reg __393803_393803;
   reg _393804_393804 ; 
   reg __393804_393804;
   reg _393805_393805 ; 
   reg __393805_393805;
   reg _393806_393806 ; 
   reg __393806_393806;
   reg _393807_393807 ; 
   reg __393807_393807;
   reg _393808_393808 ; 
   reg __393808_393808;
   reg _393809_393809 ; 
   reg __393809_393809;
   reg _393810_393810 ; 
   reg __393810_393810;
   reg _393811_393811 ; 
   reg __393811_393811;
   reg _393812_393812 ; 
   reg __393812_393812;
   reg _393813_393813 ; 
   reg __393813_393813;
   reg _393814_393814 ; 
   reg __393814_393814;
   reg _393815_393815 ; 
   reg __393815_393815;
   reg _393816_393816 ; 
   reg __393816_393816;
   reg _393817_393817 ; 
   reg __393817_393817;
   reg _393818_393818 ; 
   reg __393818_393818;
   reg _393819_393819 ; 
   reg __393819_393819;
   reg _393820_393820 ; 
   reg __393820_393820;
   reg _393821_393821 ; 
   reg __393821_393821;
   reg _393822_393822 ; 
   reg __393822_393822;
   reg _393823_393823 ; 
   reg __393823_393823;
   reg _393824_393824 ; 
   reg __393824_393824;
   reg _393825_393825 ; 
   reg __393825_393825;
   reg _393826_393826 ; 
   reg __393826_393826;
   reg _393827_393827 ; 
   reg __393827_393827;
   reg _393828_393828 ; 
   reg __393828_393828;
   reg _393829_393829 ; 
   reg __393829_393829;
   reg _393830_393830 ; 
   reg __393830_393830;
   reg _393831_393831 ; 
   reg __393831_393831;
   reg _393832_393832 ; 
   reg __393832_393832;
   reg _393833_393833 ; 
   reg __393833_393833;
   reg _393834_393834 ; 
   reg __393834_393834;
   reg _393835_393835 ; 
   reg __393835_393835;
   reg _393836_393836 ; 
   reg __393836_393836;
   reg _393837_393837 ; 
   reg __393837_393837;
   reg _393838_393838 ; 
   reg __393838_393838;
   reg _393839_393839 ; 
   reg __393839_393839;
   reg _393840_393840 ; 
   reg __393840_393840;
   reg _393841_393841 ; 
   reg __393841_393841;
   reg _393842_393842 ; 
   reg __393842_393842;
   reg _393843_393843 ; 
   reg __393843_393843;
   reg _393844_393844 ; 
   reg __393844_393844;
   reg _393845_393845 ; 
   reg __393845_393845;
   reg _393846_393846 ; 
   reg __393846_393846;
   reg _393847_393847 ; 
   reg __393847_393847;
   reg _393848_393848 ; 
   reg __393848_393848;
   reg _393849_393849 ; 
   reg __393849_393849;
   reg _393850_393850 ; 
   reg __393850_393850;
   reg _393851_393851 ; 
   reg __393851_393851;
   reg _393852_393852 ; 
   reg __393852_393852;
   reg _393853_393853 ; 
   reg __393853_393853;
   reg _393854_393854 ; 
   reg __393854_393854;
   reg _393855_393855 ; 
   reg __393855_393855;
   reg _393856_393856 ; 
   reg __393856_393856;
   reg _393857_393857 ; 
   reg __393857_393857;
   reg _393858_393858 ; 
   reg __393858_393858;
   reg _393859_393859 ; 
   reg __393859_393859;
   reg _393860_393860 ; 
   reg __393860_393860;
   reg _393861_393861 ; 
   reg __393861_393861;
   reg _393862_393862 ; 
   reg __393862_393862;
   reg _393863_393863 ; 
   reg __393863_393863;
   reg _393864_393864 ; 
   reg __393864_393864;
   reg _393865_393865 ; 
   reg __393865_393865;
   reg _393866_393866 ; 
   reg __393866_393866;
   reg _393867_393867 ; 
   reg __393867_393867;
   reg _393868_393868 ; 
   reg __393868_393868;
   reg _393869_393869 ; 
   reg __393869_393869;
   reg _393870_393870 ; 
   reg __393870_393870;
   reg _393871_393871 ; 
   reg __393871_393871;
   reg _393872_393872 ; 
   reg __393872_393872;
   reg _393873_393873 ; 
   reg __393873_393873;
   reg _393874_393874 ; 
   reg __393874_393874;
   reg _393875_393875 ; 
   reg __393875_393875;
   reg _393876_393876 ; 
   reg __393876_393876;
   reg _393877_393877 ; 
   reg __393877_393877;
   reg _393878_393878 ; 
   reg __393878_393878;
   reg _393879_393879 ; 
   reg __393879_393879;
   reg _393880_393880 ; 
   reg __393880_393880;
   reg _393881_393881 ; 
   reg __393881_393881;
   reg _393882_393882 ; 
   reg __393882_393882;
   reg _393883_393883 ; 
   reg __393883_393883;
   reg _393884_393884 ; 
   reg __393884_393884;
   reg _393885_393885 ; 
   reg __393885_393885;
   reg _393886_393886 ; 
   reg __393886_393886;
   reg _393887_393887 ; 
   reg __393887_393887;
   reg _393888_393888 ; 
   reg __393888_393888;
   reg _393889_393889 ; 
   reg __393889_393889;
   reg _393890_393890 ; 
   reg __393890_393890;
   reg _393891_393891 ; 
   reg __393891_393891;
   reg _393892_393892 ; 
   reg __393892_393892;
   reg _393893_393893 ; 
   reg __393893_393893;
   reg _393894_393894 ; 
   reg __393894_393894;
   reg _393895_393895 ; 
   reg __393895_393895;
   reg _393896_393896 ; 
   reg __393896_393896;
   reg _393897_393897 ; 
   reg __393897_393897;
   reg _393898_393898 ; 
   reg __393898_393898;
   reg _393899_393899 ; 
   reg __393899_393899;
   reg _393900_393900 ; 
   reg __393900_393900;
   reg _393901_393901 ; 
   reg __393901_393901;
   reg _393902_393902 ; 
   reg __393902_393902;
   reg _393903_393903 ; 
   reg __393903_393903;
   reg _393904_393904 ; 
   reg __393904_393904;
   reg _393905_393905 ; 
   reg __393905_393905;
   reg _393906_393906 ; 
   reg __393906_393906;
   reg _393907_393907 ; 
   reg __393907_393907;
   reg _393908_393908 ; 
   reg __393908_393908;
   reg _393909_393909 ; 
   reg __393909_393909;
   reg _393910_393910 ; 
   reg __393910_393910;
   reg _393911_393911 ; 
   reg __393911_393911;
   reg _393912_393912 ; 
   reg __393912_393912;
   reg _393913_393913 ; 
   reg __393913_393913;
   reg _393914_393914 ; 
   reg __393914_393914;
   reg _393915_393915 ; 
   reg __393915_393915;
   reg _393916_393916 ; 
   reg __393916_393916;
   reg _393917_393917 ; 
   reg __393917_393917;
   reg _393918_393918 ; 
   reg __393918_393918;
   reg _393919_393919 ; 
   reg __393919_393919;
   reg _393920_393920 ; 
   reg __393920_393920;
   reg _393921_393921 ; 
   reg __393921_393921;
   reg _393922_393922 ; 
   reg __393922_393922;
   reg _393923_393923 ; 
   reg __393923_393923;
   reg _393924_393924 ; 
   reg __393924_393924;
   reg _393925_393925 ; 
   reg __393925_393925;
   reg _393926_393926 ; 
   reg __393926_393926;
   reg _393927_393927 ; 
   reg __393927_393927;
   reg _393928_393928 ; 
   reg __393928_393928;
   reg _393929_393929 ; 
   reg __393929_393929;
   reg _393930_393930 ; 
   reg __393930_393930;
   reg _393931_393931 ; 
   reg __393931_393931;
   reg _393932_393932 ; 
   reg __393932_393932;
   reg _393933_393933 ; 
   reg __393933_393933;
   reg _393934_393934 ; 
   reg __393934_393934;
   reg _393935_393935 ; 
   reg __393935_393935;
   reg _393936_393936 ; 
   reg __393936_393936;
   reg _393937_393937 ; 
   reg __393937_393937;
   reg _393938_393938 ; 
   reg __393938_393938;
   reg _393939_393939 ; 
   reg __393939_393939;
   reg _393940_393940 ; 
   reg __393940_393940;
   reg _393941_393941 ; 
   reg __393941_393941;
   reg _393942_393942 ; 
   reg __393942_393942;
   reg _393943_393943 ; 
   reg __393943_393943;
   reg _393944_393944 ; 
   reg __393944_393944;
   reg _393945_393945 ; 
   reg __393945_393945;
   reg _393946_393946 ; 
   reg __393946_393946;
   reg _393947_393947 ; 
   reg __393947_393947;
   reg _393948_393948 ; 
   reg __393948_393948;
   reg _393949_393949 ; 
   reg __393949_393949;
   reg _393950_393950 ; 
   reg __393950_393950;
   reg _393951_393951 ; 
   reg __393951_393951;
   reg _393952_393952 ; 
   reg __393952_393952;
   reg _393953_393953 ; 
   reg __393953_393953;
   reg _393954_393954 ; 
   reg __393954_393954;
   reg _393955_393955 ; 
   reg __393955_393955;
   reg _393956_393956 ; 
   reg __393956_393956;
   reg _393957_393957 ; 
   reg __393957_393957;
   reg _393958_393958 ; 
   reg __393958_393958;
   reg _393959_393959 ; 
   reg __393959_393959;
   reg _393960_393960 ; 
   reg __393960_393960;
   reg _393961_393961 ; 
   reg __393961_393961;
   reg _393962_393962 ; 
   reg __393962_393962;
   reg _393963_393963 ; 
   reg __393963_393963;
   reg _393964_393964 ; 
   reg __393964_393964;
   reg _393965_393965 ; 
   reg __393965_393965;
   reg _393966_393966 ; 
   reg __393966_393966;
   reg _393967_393967 ; 
   reg __393967_393967;
   reg _393968_393968 ; 
   reg __393968_393968;
   reg _393969_393969 ; 
   reg __393969_393969;
   reg _393970_393970 ; 
   reg __393970_393970;
   reg _393971_393971 ; 
   reg __393971_393971;
   reg _393972_393972 ; 
   reg __393972_393972;
   reg _393973_393973 ; 
   reg __393973_393973;
   reg _393974_393974 ; 
   reg __393974_393974;
   reg _393975_393975 ; 
   reg __393975_393975;
   reg _393976_393976 ; 
   reg __393976_393976;
   reg _393977_393977 ; 
   reg __393977_393977;
   reg _393978_393978 ; 
   reg __393978_393978;
   reg _393979_393979 ; 
   reg __393979_393979;
   reg _393980_393980 ; 
   reg __393980_393980;
   reg _393981_393981 ; 
   reg __393981_393981;
   reg _393982_393982 ; 
   reg __393982_393982;
   reg _393983_393983 ; 
   reg __393983_393983;
   reg _393984_393984 ; 
   reg __393984_393984;
   reg _393985_393985 ; 
   reg __393985_393985;
   reg _393986_393986 ; 
   reg __393986_393986;
   reg _393987_393987 ; 
   reg __393987_393987;
   reg _393988_393988 ; 
   reg __393988_393988;
   reg _393989_393989 ; 
   reg __393989_393989;
   reg _393990_393990 ; 
   reg __393990_393990;
   reg _393991_393991 ; 
   reg __393991_393991;
   reg _393992_393992 ; 
   reg __393992_393992;
   reg _393993_393993 ; 
   reg __393993_393993;
   reg _393994_393994 ; 
   reg __393994_393994;
   reg _393995_393995 ; 
   reg __393995_393995;
   reg _393996_393996 ; 
   reg __393996_393996;
   reg _393997_393997 ; 
   reg __393997_393997;
   reg _393998_393998 ; 
   reg __393998_393998;
   reg _393999_393999 ; 
   reg __393999_393999;
   reg _394000_394000 ; 
   reg __394000_394000;
   reg _394001_394001 ; 
   reg __394001_394001;
   reg _394002_394002 ; 
   reg __394002_394002;
   reg _394003_394003 ; 
   reg __394003_394003;
   reg _394004_394004 ; 
   reg __394004_394004;
   reg _394005_394005 ; 
   reg __394005_394005;
   reg _394006_394006 ; 
   reg __394006_394006;
   reg _394007_394007 ; 
   reg __394007_394007;
   reg _394008_394008 ; 
   reg __394008_394008;
   reg _394009_394009 ; 
   reg __394009_394009;
   reg _394010_394010 ; 
   reg __394010_394010;
   reg _394011_394011 ; 
   reg __394011_394011;
   reg _394012_394012 ; 
   reg __394012_394012;
   reg _394013_394013 ; 
   reg __394013_394013;
   reg _394014_394014 ; 
   reg __394014_394014;
   reg _394015_394015 ; 
   reg __394015_394015;
   reg _394016_394016 ; 
   reg __394016_394016;
   reg _394017_394017 ; 
   reg __394017_394017;
   reg _394018_394018 ; 
   reg __394018_394018;
   reg _394019_394019 ; 
   reg __394019_394019;
   reg _394020_394020 ; 
   reg __394020_394020;
   reg _394021_394021 ; 
   reg __394021_394021;
   reg _394022_394022 ; 
   reg __394022_394022;
   reg _394023_394023 ; 
   reg __394023_394023;
   reg _394024_394024 ; 
   reg __394024_394024;
   reg _394025_394025 ; 
   reg __394025_394025;
   reg _394026_394026 ; 
   reg __394026_394026;
   reg _394027_394027 ; 
   reg __394027_394027;
   reg _394028_394028 ; 
   reg __394028_394028;
   reg _394029_394029 ; 
   reg __394029_394029;
   reg _394030_394030 ; 
   reg __394030_394030;
   reg _394031_394031 ; 
   reg __394031_394031;
   reg _394032_394032 ; 
   reg __394032_394032;
   reg _394033_394033 ; 
   reg __394033_394033;
   reg _394034_394034 ; 
   reg __394034_394034;
   reg _394035_394035 ; 
   reg __394035_394035;
   reg _394036_394036 ; 
   reg __394036_394036;
   reg _394037_394037 ; 
   reg __394037_394037;
   reg _394038_394038 ; 
   reg __394038_394038;
   reg _394039_394039 ; 
   reg __394039_394039;
   reg _394040_394040 ; 
   reg __394040_394040;
   reg _394041_394041 ; 
   reg __394041_394041;
   reg _394042_394042 ; 
   reg __394042_394042;
   reg _394043_394043 ; 
   reg __394043_394043;
   reg _394044_394044 ; 
   reg __394044_394044;
   reg _394045_394045 ; 
   reg __394045_394045;
   reg _394046_394046 ; 
   reg __394046_394046;
   reg _394047_394047 ; 
   reg __394047_394047;
   reg _394048_394048 ; 
   reg __394048_394048;
   reg _394049_394049 ; 
   reg __394049_394049;
   reg _394050_394050 ; 
   reg __394050_394050;
   reg _394051_394051 ; 
   reg __394051_394051;
   reg _394052_394052 ; 
   reg __394052_394052;
   reg _394053_394053 ; 
   reg __394053_394053;
   reg _394054_394054 ; 
   reg __394054_394054;
   reg _394055_394055 ; 
   reg __394055_394055;
   reg _394056_394056 ; 
   reg __394056_394056;
   reg _394057_394057 ; 
   reg __394057_394057;
   reg _394058_394058 ; 
   reg __394058_394058;
   reg _394059_394059 ; 
   reg __394059_394059;
   reg _394060_394060 ; 
   reg __394060_394060;
   reg _394061_394061 ; 
   reg __394061_394061;
   reg _394062_394062 ; 
   reg __394062_394062;
   reg _394063_394063 ; 
   reg __394063_394063;
   reg _394064_394064 ; 
   reg __394064_394064;
   reg _394065_394065 ; 
   reg __394065_394065;
   reg _394066_394066 ; 
   reg __394066_394066;
   reg _394067_394067 ; 
   reg __394067_394067;
   reg _394068_394068 ; 
   reg __394068_394068;
   reg _394069_394069 ; 
   reg __394069_394069;
   reg _394070_394070 ; 
   reg __394070_394070;
   reg _394071_394071 ; 
   reg __394071_394071;
   reg _394072_394072 ; 
   reg __394072_394072;
   reg _394073_394073 ; 
   reg __394073_394073;
   reg _394074_394074 ; 
   reg __394074_394074;
   reg _394075_394075 ; 
   reg __394075_394075;
   reg _394076_394076 ; 
   reg __394076_394076;
   reg _394077_394077 ; 
   reg __394077_394077;
   reg _394078_394078 ; 
   reg __394078_394078;
   reg _394079_394079 ; 
   reg __394079_394079;
   reg _394080_394080 ; 
   reg __394080_394080;
   reg _394081_394081 ; 
   reg __394081_394081;
   reg _394082_394082 ; 
   reg __394082_394082;
   reg _394083_394083 ; 
   reg __394083_394083;
   reg _394084_394084 ; 
   reg __394084_394084;
   reg _394085_394085 ; 
   reg __394085_394085;
   reg _394086_394086 ; 
   reg __394086_394086;
   reg _394087_394087 ; 
   reg __394087_394087;
   reg _394088_394088 ; 
   reg __394088_394088;
   reg _394089_394089 ; 
   reg __394089_394089;
   reg _394090_394090 ; 
   reg __394090_394090;
   reg _394091_394091 ; 
   reg __394091_394091;
   reg _394092_394092 ; 
   reg __394092_394092;
   reg _394093_394093 ; 
   reg __394093_394093;
   reg _394094_394094 ; 
   reg __394094_394094;
   reg _394095_394095 ; 
   reg __394095_394095;
   reg _394096_394096 ; 
   reg __394096_394096;
   reg _394097_394097 ; 
   reg __394097_394097;
   reg _394098_394098 ; 
   reg __394098_394098;
   reg _394099_394099 ; 
   reg __394099_394099;
   reg _394100_394100 ; 
   reg __394100_394100;
   reg _394101_394101 ; 
   reg __394101_394101;
   reg _394102_394102 ; 
   reg __394102_394102;
   reg _394103_394103 ; 
   reg __394103_394103;
   reg _394104_394104 ; 
   reg __394104_394104;
   reg _394105_394105 ; 
   reg __394105_394105;
   reg _394106_394106 ; 
   reg __394106_394106;
   reg _394107_394107 ; 
   reg __394107_394107;
   reg _394108_394108 ; 
   reg __394108_394108;
   reg _394109_394109 ; 
   reg __394109_394109;
   reg _394110_394110 ; 
   reg __394110_394110;
   reg _394111_394111 ; 
   reg __394111_394111;
   reg _394112_394112 ; 
   reg __394112_394112;
   reg _394113_394113 ; 
   reg __394113_394113;
   reg _394114_394114 ; 
   reg __394114_394114;
   reg _394115_394115 ; 
   reg __394115_394115;
   reg _394116_394116 ; 
   reg __394116_394116;
   reg _394117_394117 ; 
   reg __394117_394117;
   reg _394118_394118 ; 
   reg __394118_394118;
   reg _394119_394119 ; 
   reg __394119_394119;
   reg _394120_394120 ; 
   reg __394120_394120;
   reg _394121_394121 ; 
   reg __394121_394121;
   reg _394122_394122 ; 
   reg __394122_394122;
   reg _394123_394123 ; 
   reg __394123_394123;
   reg _394124_394124 ; 
   reg __394124_394124;
   reg _394125_394125 ; 
   reg __394125_394125;
   reg _394126_394126 ; 
   reg __394126_394126;
   reg _394127_394127 ; 
   reg __394127_394127;
   reg _394128_394128 ; 
   reg __394128_394128;
   reg _394129_394129 ; 
   reg __394129_394129;
   reg _394130_394130 ; 
   reg __394130_394130;
   reg _394131_394131 ; 
   reg __394131_394131;
   reg _394132_394132 ; 
   reg __394132_394132;
   reg _394133_394133 ; 
   reg __394133_394133;
   reg _394134_394134 ; 
   reg __394134_394134;
   reg _394135_394135 ; 
   reg __394135_394135;
   reg _394136_394136 ; 
   reg __394136_394136;
   reg _394137_394137 ; 
   reg __394137_394137;
   reg _394138_394138 ; 
   reg __394138_394138;
   reg _394139_394139 ; 
   reg __394139_394139;
   reg _394140_394140 ; 
   reg __394140_394140;
   reg _394141_394141 ; 
   reg __394141_394141;
   reg _394142_394142 ; 
   reg __394142_394142;
   reg _394143_394143 ; 
   reg __394143_394143;
   reg _394144_394144 ; 
   reg __394144_394144;
   reg _394145_394145 ; 
   reg __394145_394145;
   reg _394146_394146 ; 
   reg __394146_394146;
   reg _394147_394147 ; 
   reg __394147_394147;
   reg _394148_394148 ; 
   reg __394148_394148;
   reg _394149_394149 ; 
   reg __394149_394149;
   reg _394150_394150 ; 
   reg __394150_394150;
   reg _394151_394151 ; 
   reg __394151_394151;
   reg _394152_394152 ; 
   reg __394152_394152;
   reg _394153_394153 ; 
   reg __394153_394153;
   reg _394154_394154 ; 
   reg __394154_394154;
   reg _394155_394155 ; 
   reg __394155_394155;
   reg _394156_394156 ; 
   reg __394156_394156;
   reg _394157_394157 ; 
   reg __394157_394157;
   reg _394158_394158 ; 
   reg __394158_394158;
   reg _394159_394159 ; 
   reg __394159_394159;
   reg _394160_394160 ; 
   reg __394160_394160;
   reg _394161_394161 ; 
   reg __394161_394161;
   reg _394162_394162 ; 
   reg __394162_394162;
   reg _394163_394163 ; 
   reg __394163_394163;
   reg _394164_394164 ; 
   reg __394164_394164;
   reg _394165_394165 ; 
   reg __394165_394165;
   reg _394166_394166 ; 
   reg __394166_394166;
   reg _394167_394167 ; 
   reg __394167_394167;
   reg _394168_394168 ; 
   reg __394168_394168;
   reg _394169_394169 ; 
   reg __394169_394169;
   reg _394170_394170 ; 
   reg __394170_394170;
   reg _394171_394171 ; 
   reg __394171_394171;
   reg _394172_394172 ; 
   reg __394172_394172;
   reg _394173_394173 ; 
   reg __394173_394173;
   reg _394174_394174 ; 
   reg __394174_394174;
   reg _394175_394175 ; 
   reg __394175_394175;
   reg _394176_394176 ; 
   reg __394176_394176;
   reg _394177_394177 ; 
   reg __394177_394177;
   reg _394178_394178 ; 
   reg __394178_394178;
   reg _394179_394179 ; 
   reg __394179_394179;
   reg _394180_394180 ; 
   reg __394180_394180;
   reg _394181_394181 ; 
   reg __394181_394181;
   reg _394182_394182 ; 
   reg __394182_394182;
   reg _394183_394183 ; 
   reg __394183_394183;
   reg _394184_394184 ; 
   reg __394184_394184;
   reg _394185_394185 ; 
   reg __394185_394185;
   reg _394186_394186 ; 
   reg __394186_394186;
   reg _394187_394187 ; 
   reg __394187_394187;
   reg _394188_394188 ; 
   reg __394188_394188;
   reg _394189_394189 ; 
   reg __394189_394189;
   reg _394190_394190 ; 
   reg __394190_394190;
   reg _394191_394191 ; 
   reg __394191_394191;
   reg _394192_394192 ; 
   reg __394192_394192;
   reg _394193_394193 ; 
   reg __394193_394193;
   reg _394194_394194 ; 
   reg __394194_394194;
   reg _394195_394195 ; 
   reg __394195_394195;
   reg _394196_394196 ; 
   reg __394196_394196;
   reg _394197_394197 ; 
   reg __394197_394197;
   reg _394198_394198 ; 
   reg __394198_394198;
   reg _394199_394199 ; 
   reg __394199_394199;
   reg _394200_394200 ; 
   reg __394200_394200;
   reg _394201_394201 ; 
   reg __394201_394201;
   reg _394202_394202 ; 
   reg __394202_394202;
   reg _394203_394203 ; 
   reg __394203_394203;
   reg _394204_394204 ; 
   reg __394204_394204;
   reg _394205_394205 ; 
   reg __394205_394205;
   reg _394206_394206 ; 
   reg __394206_394206;
   reg _394207_394207 ; 
   reg __394207_394207;
   reg _394208_394208 ; 
   reg __394208_394208;
   reg _394209_394209 ; 
   reg __394209_394209;
   reg _394210_394210 ; 
   reg __394210_394210;
   reg _394211_394211 ; 
   reg __394211_394211;
   reg _394212_394212 ; 
   reg __394212_394212;
   reg _394213_394213 ; 
   reg __394213_394213;
   reg _394214_394214 ; 
   reg __394214_394214;
   reg _394215_394215 ; 
   reg __394215_394215;
   reg _394216_394216 ; 
   reg __394216_394216;
   reg _394217_394217 ; 
   reg __394217_394217;
   reg _394218_394218 ; 
   reg __394218_394218;
   reg _394219_394219 ; 
   reg __394219_394219;
   reg _394220_394220 ; 
   reg __394220_394220;
   reg _394221_394221 ; 
   reg __394221_394221;
   reg _394222_394222 ; 
   reg __394222_394222;
   reg _394223_394223 ; 
   reg __394223_394223;
   reg _394224_394224 ; 
   reg __394224_394224;
   reg _394225_394225 ; 
   reg __394225_394225;
   reg _394226_394226 ; 
   reg __394226_394226;
   reg _394227_394227 ; 
   reg __394227_394227;
   reg _394228_394228 ; 
   reg __394228_394228;
   reg _394229_394229 ; 
   reg __394229_394229;
   reg _394230_394230 ; 
   reg __394230_394230;
   reg _394231_394231 ; 
   reg __394231_394231;
   reg _394232_394232 ; 
   reg __394232_394232;
   reg _394233_394233 ; 
   reg __394233_394233;
   reg _394234_394234 ; 
   reg __394234_394234;
   reg _394235_394235 ; 
   reg __394235_394235;
   reg _394236_394236 ; 
   reg __394236_394236;
   reg _394237_394237 ; 
   reg __394237_394237;
   reg _394238_394238 ; 
   reg __394238_394238;
   reg _394239_394239 ; 
   reg __394239_394239;
   reg _394240_394240 ; 
   reg __394240_394240;
   reg _394241_394241 ; 
   reg __394241_394241;
   reg _394242_394242 ; 
   reg __394242_394242;
   reg _394243_394243 ; 
   reg __394243_394243;
   reg _394244_394244 ; 
   reg __394244_394244;
   reg _394245_394245 ; 
   reg __394245_394245;
   reg _394246_394246 ; 
   reg __394246_394246;
   reg _394247_394247 ; 
   reg __394247_394247;
   reg _394248_394248 ; 
   reg __394248_394248;
   reg _394249_394249 ; 
   reg __394249_394249;
   reg _394250_394250 ; 
   reg __394250_394250;
   reg _394251_394251 ; 
   reg __394251_394251;
   reg _394252_394252 ; 
   reg __394252_394252;
   reg _394253_394253 ; 
   reg __394253_394253;
   reg _394254_394254 ; 
   reg __394254_394254;
   reg _394255_394255 ; 
   reg __394255_394255;
   reg _394256_394256 ; 
   reg __394256_394256;
   reg _394257_394257 ; 
   reg __394257_394257;
   reg _394258_394258 ; 
   reg __394258_394258;
   reg _394259_394259 ; 
   reg __394259_394259;
   reg _394260_394260 ; 
   reg __394260_394260;
   reg _394261_394261 ; 
   reg __394261_394261;
   reg _394262_394262 ; 
   reg __394262_394262;
   reg _394263_394263 ; 
   reg __394263_394263;
   reg _394264_394264 ; 
   reg __394264_394264;
   reg _394265_394265 ; 
   reg __394265_394265;
   reg _394266_394266 ; 
   reg __394266_394266;
   reg _394267_394267 ; 
   reg __394267_394267;
   reg _394268_394268 ; 
   reg __394268_394268;
   reg _394269_394269 ; 
   reg __394269_394269;
   reg _394270_394270 ; 
   reg __394270_394270;
   reg _394271_394271 ; 
   reg __394271_394271;
   reg _394272_394272 ; 
   reg __394272_394272;
   reg _394273_394273 ; 
   reg __394273_394273;
   reg _394274_394274 ; 
   reg __394274_394274;
   reg _394275_394275 ; 
   reg __394275_394275;
   reg _394276_394276 ; 
   reg __394276_394276;
   reg _394277_394277 ; 
   reg __394277_394277;
   reg _394278_394278 ; 
   reg __394278_394278;
   reg _394279_394279 ; 
   reg __394279_394279;
   reg _394280_394280 ; 
   reg __394280_394280;
   reg _394281_394281 ; 
   reg __394281_394281;
   reg _394282_394282 ; 
   reg __394282_394282;
   reg _394283_394283 ; 
   reg __394283_394283;
   reg _394284_394284 ; 
   reg __394284_394284;
   reg _394285_394285 ; 
   reg __394285_394285;
   reg _394286_394286 ; 
   reg __394286_394286;
   reg _394287_394287 ; 
   reg __394287_394287;
   reg _394288_394288 ; 
   reg __394288_394288;
   reg _394289_394289 ; 
   reg __394289_394289;
   reg _394290_394290 ; 
   reg __394290_394290;
   reg _394291_394291 ; 
   reg __394291_394291;
   reg _394292_394292 ; 
   reg __394292_394292;
   reg _394293_394293 ; 
   reg __394293_394293;
   reg _394294_394294 ; 
   reg __394294_394294;
   reg _394295_394295 ; 
   reg __394295_394295;
   reg _394296_394296 ; 
   reg __394296_394296;
   reg _394297_394297 ; 
   reg __394297_394297;
   reg _394298_394298 ; 
   reg __394298_394298;
   reg _394299_394299 ; 
   reg __394299_394299;
   reg _394300_394300 ; 
   reg __394300_394300;
   reg _394301_394301 ; 
   reg __394301_394301;
   reg _394302_394302 ; 
   reg __394302_394302;
   reg _394303_394303 ; 
   reg __394303_394303;
   reg _394304_394304 ; 
   reg __394304_394304;
   reg _394305_394305 ; 
   reg __394305_394305;
   reg _394306_394306 ; 
   reg __394306_394306;
   reg _394307_394307 ; 
   reg __394307_394307;
   reg _394308_394308 ; 
   reg __394308_394308;
   reg _394309_394309 ; 
   reg __394309_394309;
   reg _394310_394310 ; 
   reg __394310_394310;
   reg _394311_394311 ; 
   reg __394311_394311;
   reg _394312_394312 ; 
   reg __394312_394312;
   reg _394313_394313 ; 
   reg __394313_394313;
   reg _394314_394314 ; 
   reg __394314_394314;
   reg _394315_394315 ; 
   reg __394315_394315;
   reg _394316_394316 ; 
   reg __394316_394316;
   reg _394317_394317 ; 
   reg __394317_394317;
   reg _394318_394318 ; 
   reg __394318_394318;
   reg _394319_394319 ; 
   reg __394319_394319;
   reg _394320_394320 ; 
   reg __394320_394320;
   reg _394321_394321 ; 
   reg __394321_394321;
   reg _394322_394322 ; 
   reg __394322_394322;
   reg _394323_394323 ; 
   reg __394323_394323;
   reg _394324_394324 ; 
   reg __394324_394324;
   reg _394325_394325 ; 
   reg __394325_394325;
   reg _394326_394326 ; 
   reg __394326_394326;
   reg _394327_394327 ; 
   reg __394327_394327;
   reg _394328_394328 ; 
   reg __394328_394328;
   reg _394329_394329 ; 
   reg __394329_394329;
   reg _394330_394330 ; 
   reg __394330_394330;
   reg _394331_394331 ; 
   reg __394331_394331;
   reg _394332_394332 ; 
   reg __394332_394332;
   reg _394333_394333 ; 
   reg __394333_394333;
   reg _394334_394334 ; 
   reg __394334_394334;
   reg _394335_394335 ; 
   reg __394335_394335;
   reg _394336_394336 ; 
   reg __394336_394336;
   reg _394337_394337 ; 
   reg __394337_394337;
   reg _394338_394338 ; 
   reg __394338_394338;
   reg _394339_394339 ; 
   reg __394339_394339;
   reg _394340_394340 ; 
   reg __394340_394340;
   reg _394341_394341 ; 
   reg __394341_394341;
   reg _394342_394342 ; 
   reg __394342_394342;
   reg _394343_394343 ; 
   reg __394343_394343;
   reg _394344_394344 ; 
   reg __394344_394344;
   reg _394345_394345 ; 
   reg __394345_394345;
   reg _394346_394346 ; 
   reg __394346_394346;
   reg _394347_394347 ; 
   reg __394347_394347;
   reg _394348_394348 ; 
   reg __394348_394348;
   reg _394349_394349 ; 
   reg __394349_394349;
   reg _394350_394350 ; 
   reg __394350_394350;
   reg _394351_394351 ; 
   reg __394351_394351;
   reg _394352_394352 ; 
   reg __394352_394352;
   reg _394353_394353 ; 
   reg __394353_394353;
   reg _394354_394354 ; 
   reg __394354_394354;
   reg _394355_394355 ; 
   reg __394355_394355;
   reg _394356_394356 ; 
   reg __394356_394356;
   reg _394357_394357 ; 
   reg __394357_394357;
   reg _394358_394358 ; 
   reg __394358_394358;
   reg _394359_394359 ; 
   reg __394359_394359;
   reg _394360_394360 ; 
   reg __394360_394360;
   reg _394361_394361 ; 
   reg __394361_394361;
   reg _394362_394362 ; 
   reg __394362_394362;
   reg _394363_394363 ; 
   reg __394363_394363;
   reg _394364_394364 ; 
   reg __394364_394364;
   reg _394365_394365 ; 
   reg __394365_394365;
   reg _394366_394366 ; 
   reg __394366_394366;
   reg _394367_394367 ; 
   reg __394367_394367;
   reg _394368_394368 ; 
   reg __394368_394368;
   reg _394369_394369 ; 
   reg __394369_394369;
   reg _394370_394370 ; 
   reg __394370_394370;
   reg _394371_394371 ; 
   reg __394371_394371;
   reg _394372_394372 ; 
   reg __394372_394372;
   reg _394373_394373 ; 
   reg __394373_394373;
   reg _394374_394374 ; 
   reg __394374_394374;
   reg _394375_394375 ; 
   reg __394375_394375;
   reg _394376_394376 ; 
   reg __394376_394376;
   reg _394377_394377 ; 
   reg __394377_394377;
   reg _394378_394378 ; 
   reg __394378_394378;
   reg _394379_394379 ; 
   reg __394379_394379;
   reg _394380_394380 ; 
   reg __394380_394380;
   reg _394381_394381 ; 
   reg __394381_394381;
   reg _394382_394382 ; 
   reg __394382_394382;
   reg _394383_394383 ; 
   reg __394383_394383;
   reg _394384_394384 ; 
   reg __394384_394384;
   reg _394385_394385 ; 
   reg __394385_394385;
   reg _394386_394386 ; 
   reg __394386_394386;
   reg _394387_394387 ; 
   reg __394387_394387;
   reg _394388_394388 ; 
   reg __394388_394388;
   reg _394389_394389 ; 
   reg __394389_394389;
   reg _394390_394390 ; 
   reg __394390_394390;
   reg _394391_394391 ; 
   reg __394391_394391;
   reg _394392_394392 ; 
   reg __394392_394392;
   reg _394393_394393 ; 
   reg __394393_394393;
   reg _394394_394394 ; 
   reg __394394_394394;
   reg _394395_394395 ; 
   reg __394395_394395;
   reg _394396_394396 ; 
   reg __394396_394396;
   reg _394397_394397 ; 
   reg __394397_394397;
   reg _394398_394398 ; 
   reg __394398_394398;
   reg _394399_394399 ; 
   reg __394399_394399;
   reg _394400_394400 ; 
   reg __394400_394400;
   reg _394401_394401 ; 
   reg __394401_394401;
   reg _394402_394402 ; 
   reg __394402_394402;
   reg _394403_394403 ; 
   reg __394403_394403;
   reg _394404_394404 ; 
   reg __394404_394404;
   reg _394405_394405 ; 
   reg __394405_394405;
   reg _394406_394406 ; 
   reg __394406_394406;
   reg _394407_394407 ; 
   reg __394407_394407;
   reg _394408_394408 ; 
   reg __394408_394408;
   reg _394409_394409 ; 
   reg __394409_394409;
   reg _394410_394410 ; 
   reg __394410_394410;
   reg _394411_394411 ; 
   reg __394411_394411;
   reg _394412_394412 ; 
   reg __394412_394412;
   reg _394413_394413 ; 
   reg __394413_394413;
   reg _394414_394414 ; 
   reg __394414_394414;
   reg _394415_394415 ; 
   reg __394415_394415;
   reg _394416_394416 ; 
   reg __394416_394416;
   reg _394417_394417 ; 
   reg __394417_394417;
   reg _394418_394418 ; 
   reg __394418_394418;
   reg _394419_394419 ; 
   reg __394419_394419;
   reg _394420_394420 ; 
   reg __394420_394420;
   reg _394421_394421 ; 
   reg __394421_394421;
   reg _394422_394422 ; 
   reg __394422_394422;
   reg _394423_394423 ; 
   reg __394423_394423;
   reg _394424_394424 ; 
   reg __394424_394424;
   reg _394425_394425 ; 
   reg __394425_394425;
   reg _394426_394426 ; 
   reg __394426_394426;
   reg _394427_394427 ; 
   reg __394427_394427;
   reg _394428_394428 ; 
   reg __394428_394428;
   reg _394429_394429 ; 
   reg __394429_394429;
   reg _394430_394430 ; 
   reg __394430_394430;
   reg _394431_394431 ; 
   reg __394431_394431;
   reg _394432_394432 ; 
   reg __394432_394432;
   reg _394433_394433 ; 
   reg __394433_394433;
   reg _394434_394434 ; 
   reg __394434_394434;
   reg _394435_394435 ; 
   reg __394435_394435;
   reg _394436_394436 ; 
   reg __394436_394436;
   reg _394437_394437 ; 
   reg __394437_394437;
   reg _394438_394438 ; 
   reg __394438_394438;
   reg _394439_394439 ; 
   reg __394439_394439;
   reg _394440_394440 ; 
   reg __394440_394440;
   reg _394441_394441 ; 
   reg __394441_394441;
   reg _394442_394442 ; 
   reg __394442_394442;
   reg _394443_394443 ; 
   reg __394443_394443;
   reg _394444_394444 ; 
   reg __394444_394444;
   reg _394445_394445 ; 
   reg __394445_394445;
   reg _394446_394446 ; 
   reg __394446_394446;
   reg _394447_394447 ; 
   reg __394447_394447;
   reg _394448_394448 ; 
   reg __394448_394448;
   reg _394449_394449 ; 
   reg __394449_394449;
   reg _394450_394450 ; 
   reg __394450_394450;
   reg _394451_394451 ; 
   reg __394451_394451;
   reg _394452_394452 ; 
   reg __394452_394452;
   reg _394453_394453 ; 
   reg __394453_394453;
   reg _394454_394454 ; 
   reg __394454_394454;
   reg _394455_394455 ; 
   reg __394455_394455;
   reg _394456_394456 ; 
   reg __394456_394456;
   reg _394457_394457 ; 
   reg __394457_394457;
   reg _394458_394458 ; 
   reg __394458_394458;
   reg _394459_394459 ; 
   reg __394459_394459;
   reg _394460_394460 ; 
   reg __394460_394460;
   reg _394461_394461 ; 
   reg __394461_394461;
   reg _394462_394462 ; 
   reg __394462_394462;
   reg _394463_394463 ; 
   reg __394463_394463;
   reg _394464_394464 ; 
   reg __394464_394464;
   reg _394465_394465 ; 
   reg __394465_394465;
   reg _394466_394466 ; 
   reg __394466_394466;
   reg _394467_394467 ; 
   reg __394467_394467;
   reg _394468_394468 ; 
   reg __394468_394468;
   reg _394469_394469 ; 
   reg __394469_394469;
   reg _394470_394470 ; 
   reg __394470_394470;
   reg _394471_394471 ; 
   reg __394471_394471;
   reg _394472_394472 ; 
   reg __394472_394472;
   reg _394473_394473 ; 
   reg __394473_394473;
   reg _394474_394474 ; 
   reg __394474_394474;
   reg _394475_394475 ; 
   reg __394475_394475;
   reg _394476_394476 ; 
   reg __394476_394476;
   reg _394477_394477 ; 
   reg __394477_394477;
   reg _394478_394478 ; 
   reg __394478_394478;
   reg _394479_394479 ; 
   reg __394479_394479;
   reg _394480_394480 ; 
   reg __394480_394480;
   reg _394481_394481 ; 
   reg __394481_394481;
   reg _394482_394482 ; 
   reg __394482_394482;
   reg _394483_394483 ; 
   reg __394483_394483;
   reg _394484_394484 ; 
   reg __394484_394484;
   reg _394485_394485 ; 
   reg __394485_394485;
   reg _394486_394486 ; 
   reg __394486_394486;
   reg _394487_394487 ; 
   reg __394487_394487;
   reg _394488_394488 ; 
   reg __394488_394488;
   reg _394489_394489 ; 
   reg __394489_394489;
   reg _394490_394490 ; 
   reg __394490_394490;
   reg _394491_394491 ; 
   reg __394491_394491;
   reg _394492_394492 ; 
   reg __394492_394492;
   reg _394493_394493 ; 
   reg __394493_394493;
   reg _394494_394494 ; 
   reg __394494_394494;
   reg _394495_394495 ; 
   reg __394495_394495;
   reg _394496_394496 ; 
   reg __394496_394496;
   reg _394497_394497 ; 
   reg __394497_394497;
   reg _394498_394498 ; 
   reg __394498_394498;
   reg _394499_394499 ; 
   reg __394499_394499;
   reg _394500_394500 ; 
   reg __394500_394500;
   reg _394501_394501 ; 
   reg __394501_394501;
   reg _394502_394502 ; 
   reg __394502_394502;
   reg _394503_394503 ; 
   reg __394503_394503;
   reg _394504_394504 ; 
   reg __394504_394504;
   reg _394505_394505 ; 
   reg __394505_394505;
   reg _394506_394506 ; 
   reg __394506_394506;
   reg _394507_394507 ; 
   reg __394507_394507;
   reg _394508_394508 ; 
   reg __394508_394508;
   reg _394509_394509 ; 
   reg __394509_394509;
   reg _394510_394510 ; 
   reg __394510_394510;
   reg _394511_394511 ; 
   reg __394511_394511;
   reg _394512_394512 ; 
   reg __394512_394512;
   reg _394513_394513 ; 
   reg __394513_394513;
   reg _394514_394514 ; 
   reg __394514_394514;
   reg _394515_394515 ; 
   reg __394515_394515;
   reg _394516_394516 ; 
   reg __394516_394516;
   reg _394517_394517 ; 
   reg __394517_394517;
   reg _394518_394518 ; 
   reg __394518_394518;
   reg _394519_394519 ; 
   reg __394519_394519;
   reg _394520_394520 ; 
   reg __394520_394520;
   reg _394521_394521 ; 
   reg __394521_394521;
   reg _394522_394522 ; 
   reg __394522_394522;
   reg _394523_394523 ; 
   reg __394523_394523;
   reg _394524_394524 ; 
   reg __394524_394524;
   reg _394525_394525 ; 
   reg __394525_394525;
   reg _394526_394526 ; 
   reg __394526_394526;
   reg _394527_394527 ; 
   reg __394527_394527;
   reg _394528_394528 ; 
   reg __394528_394528;
   reg _394529_394529 ; 
   reg __394529_394529;
   reg _394530_394530 ; 
   reg __394530_394530;
   reg _394531_394531 ; 
   reg __394531_394531;
   reg _394532_394532 ; 
   reg __394532_394532;
   reg _394533_394533 ; 
   reg __394533_394533;
   reg _394534_394534 ; 
   reg __394534_394534;
   reg _394535_394535 ; 
   reg __394535_394535;
   reg _394536_394536 ; 
   reg __394536_394536;
   reg _394537_394537 ; 
   reg __394537_394537;
   reg _394538_394538 ; 
   reg __394538_394538;
   reg _394539_394539 ; 
   reg __394539_394539;
   reg _394540_394540 ; 
   reg __394540_394540;
   reg _394541_394541 ; 
   reg __394541_394541;
   reg _394542_394542 ; 
   reg __394542_394542;
   reg _394543_394543 ; 
   reg __394543_394543;
   reg _394544_394544 ; 
   reg __394544_394544;
   reg _394545_394545 ; 
   reg __394545_394545;
   reg _394546_394546 ; 
   reg __394546_394546;
   reg _394547_394547 ; 
   reg __394547_394547;
   reg _394548_394548 ; 
   reg __394548_394548;
   reg _394549_394549 ; 
   reg __394549_394549;
   reg _394550_394550 ; 
   reg __394550_394550;
   reg _394551_394551 ; 
   reg __394551_394551;
   reg _394552_394552 ; 
   reg __394552_394552;
   reg _394553_394553 ; 
   reg __394553_394553;
   reg _394554_394554 ; 
   reg __394554_394554;
   reg _394555_394555 ; 
   reg __394555_394555;
   reg _394556_394556 ; 
   reg __394556_394556;
   reg _394557_394557 ; 
   reg __394557_394557;
   reg _394558_394558 ; 
   reg __394558_394558;
   reg _394559_394559 ; 
   reg __394559_394559;
   reg _394560_394560 ; 
   reg __394560_394560;
   reg _394561_394561 ; 
   reg __394561_394561;
   reg _394562_394562 ; 
   reg __394562_394562;
   reg _394563_394563 ; 
   reg __394563_394563;
   reg _394564_394564 ; 
   reg __394564_394564;
   reg _394565_394565 ; 
   reg __394565_394565;
   reg _394566_394566 ; 
   reg __394566_394566;
   reg _394567_394567 ; 
   reg __394567_394567;
   reg _394568_394568 ; 
   reg __394568_394568;
   reg _394569_394569 ; 
   reg __394569_394569;
   reg _394570_394570 ; 
   reg __394570_394570;
   reg _394571_394571 ; 
   reg __394571_394571;
   reg _394572_394572 ; 
   reg __394572_394572;
   reg _394573_394573 ; 
   reg __394573_394573;
   reg _394574_394574 ; 
   reg __394574_394574;
   reg _394575_394575 ; 
   reg __394575_394575;
   reg _394576_394576 ; 
   reg __394576_394576;
   reg _394577_394577 ; 
   reg __394577_394577;
   reg _394578_394578 ; 
   reg __394578_394578;
   reg _394579_394579 ; 
   reg __394579_394579;
   reg _394580_394580 ; 
   reg __394580_394580;
   reg _394581_394581 ; 
   reg __394581_394581;
   reg _394582_394582 ; 
   reg __394582_394582;
   reg _394583_394583 ; 
   reg __394583_394583;
   reg _394584_394584 ; 
   reg __394584_394584;
   reg _394585_394585 ; 
   reg __394585_394585;
   reg _394586_394586 ; 
   reg __394586_394586;
   reg _394587_394587 ; 
   reg __394587_394587;
   reg _394588_394588 ; 
   reg __394588_394588;
   reg _394589_394589 ; 
   reg __394589_394589;
   reg _394590_394590 ; 
   reg __394590_394590;
   reg _394591_394591 ; 
   reg __394591_394591;
   reg _394592_394592 ; 
   reg __394592_394592;
   reg _394593_394593 ; 
   reg __394593_394593;
   reg _394594_394594 ; 
   reg __394594_394594;
   reg _394595_394595 ; 
   reg __394595_394595;
   reg _394596_394596 ; 
   reg __394596_394596;
   reg _394597_394597 ; 
   reg __394597_394597;
   reg _394598_394598 ; 
   reg __394598_394598;
   reg _394599_394599 ; 
   reg __394599_394599;
   reg _394600_394600 ; 
   reg __394600_394600;
   reg _394601_394601 ; 
   reg __394601_394601;
   reg _394602_394602 ; 
   reg __394602_394602;
   reg _394603_394603 ; 
   reg __394603_394603;
   reg _394604_394604 ; 
   reg __394604_394604;
   reg _394605_394605 ; 
   reg __394605_394605;
   reg _394606_394606 ; 
   reg __394606_394606;
   reg _394607_394607 ; 
   reg __394607_394607;
   reg _394608_394608 ; 
   reg __394608_394608;
   reg _394609_394609 ; 
   reg __394609_394609;
   reg _394610_394610 ; 
   reg __394610_394610;
   reg _394611_394611 ; 
   reg __394611_394611;
   reg _394612_394612 ; 
   reg __394612_394612;
   reg _394613_394613 ; 
   reg __394613_394613;
   reg _394614_394614 ; 
   reg __394614_394614;
   reg _394615_394615 ; 
   reg __394615_394615;
   reg _394616_394616 ; 
   reg __394616_394616;
   reg _394617_394617 ; 
   reg __394617_394617;
   reg _394618_394618 ; 
   reg __394618_394618;
   reg _394619_394619 ; 
   reg __394619_394619;
   reg _394620_394620 ; 
   reg __394620_394620;
   reg _394621_394621 ; 
   reg __394621_394621;
   reg _394622_394622 ; 
   reg __394622_394622;
   reg _394623_394623 ; 
   reg __394623_394623;
   reg _394624_394624 ; 
   reg __394624_394624;
   reg _394625_394625 ; 
   reg __394625_394625;
   reg _394626_394626 ; 
   reg __394626_394626;
   reg _394627_394627 ; 
   reg __394627_394627;
   reg _394628_394628 ; 
   reg __394628_394628;
   reg _394629_394629 ; 
   reg __394629_394629;
   reg _394630_394630 ; 
   reg __394630_394630;
   reg _394631_394631 ; 
   reg __394631_394631;
   reg _394632_394632 ; 
   reg __394632_394632;
   reg _394633_394633 ; 
   reg __394633_394633;
   reg _394634_394634 ; 
   reg __394634_394634;
   reg _394635_394635 ; 
   reg __394635_394635;
   reg _394636_394636 ; 
   reg __394636_394636;
   reg _394637_394637 ; 
   reg __394637_394637;
   reg _394638_394638 ; 
   reg __394638_394638;
   reg _394639_394639 ; 
   reg __394639_394639;
   reg _394640_394640 ; 
   reg __394640_394640;
   reg _394641_394641 ; 
   reg __394641_394641;
   reg _394642_394642 ; 
   reg __394642_394642;
   reg _394643_394643 ; 
   reg __394643_394643;
   reg _394644_394644 ; 
   reg __394644_394644;
   reg _394645_394645 ; 
   reg __394645_394645;
   reg _394646_394646 ; 
   reg __394646_394646;
   reg _394647_394647 ; 
   reg __394647_394647;
   reg _394648_394648 ; 
   reg __394648_394648;
   reg _394649_394649 ; 
   reg __394649_394649;
   reg _394650_394650 ; 
   reg __394650_394650;
   reg _394651_394651 ; 
   reg __394651_394651;
   reg _394652_394652 ; 
   reg __394652_394652;
   reg _394653_394653 ; 
   reg __394653_394653;
   reg _394654_394654 ; 
   reg __394654_394654;
   reg _394655_394655 ; 
   reg __394655_394655;
   reg _394656_394656 ; 
   reg __394656_394656;
   reg _394657_394657 ; 
   reg __394657_394657;
   reg _394658_394658 ; 
   reg __394658_394658;
   reg _394659_394659 ; 
   reg __394659_394659;
   reg _394660_394660 ; 
   reg __394660_394660;
   reg _394661_394661 ; 
   reg __394661_394661;
   reg _394662_394662 ; 
   reg __394662_394662;
   reg _394663_394663 ; 
   reg __394663_394663;
   reg _394664_394664 ; 
   reg __394664_394664;
   reg _394665_394665 ; 
   reg __394665_394665;
   reg _394666_394666 ; 
   reg __394666_394666;
   reg _394667_394667 ; 
   reg __394667_394667;
   reg _394668_394668 ; 
   reg __394668_394668;
   reg _394669_394669 ; 
   reg __394669_394669;
   reg _394670_394670 ; 
   reg __394670_394670;
   reg _394671_394671 ; 
   reg __394671_394671;
   reg _394672_394672 ; 
   reg __394672_394672;
   reg _394673_394673 ; 
   reg __394673_394673;
   reg _394674_394674 ; 
   reg __394674_394674;
   reg _394675_394675 ; 
   reg __394675_394675;
   reg _394676_394676 ; 
   reg __394676_394676;
   reg _394677_394677 ; 
   reg __394677_394677;
   reg _394678_394678 ; 
   reg __394678_394678;
   reg _394679_394679 ; 
   reg __394679_394679;
   reg _394680_394680 ; 
   reg __394680_394680;
   reg _394681_394681 ; 
   reg __394681_394681;
   reg _394682_394682 ; 
   reg __394682_394682;
   reg _394683_394683 ; 
   reg __394683_394683;
   reg _394684_394684 ; 
   reg __394684_394684;
   reg _394685_394685 ; 
   reg __394685_394685;
   reg _394686_394686 ; 
   reg __394686_394686;
   reg _394687_394687 ; 
   reg __394687_394687;
   reg _394688_394688 ; 
   reg __394688_394688;
   reg _394689_394689 ; 
   reg __394689_394689;
   reg _394690_394690 ; 
   reg __394690_394690;
   reg _394691_394691 ; 
   reg __394691_394691;
   reg _394692_394692 ; 
   reg __394692_394692;
   reg _394693_394693 ; 
   reg __394693_394693;
   reg _394694_394694 ; 
   reg __394694_394694;
   reg _394695_394695 ; 
   reg __394695_394695;
   reg _394696_394696 ; 
   reg __394696_394696;
   reg _394697_394697 ; 
   reg __394697_394697;
   reg _394698_394698 ; 
   reg __394698_394698;
   reg _394699_394699 ; 
   reg __394699_394699;
   reg _394700_394700 ; 
   reg __394700_394700;
   reg _394701_394701 ; 
   reg __394701_394701;
   reg _394702_394702 ; 
   reg __394702_394702;
   reg _394703_394703 ; 
   reg __394703_394703;
   reg _394704_394704 ; 
   reg __394704_394704;
   reg _394705_394705 ; 
   reg __394705_394705;
   reg _394706_394706 ; 
   reg __394706_394706;
   reg _394707_394707 ; 
   reg __394707_394707;
   reg _394708_394708 ; 
   reg __394708_394708;
   reg _394709_394709 ; 
   reg __394709_394709;
   reg _394710_394710 ; 
   reg __394710_394710;
   reg _394711_394711 ; 
   reg __394711_394711;
   reg _394712_394712 ; 
   reg __394712_394712;
   reg _394713_394713 ; 
   reg __394713_394713;
   reg _394714_394714 ; 
   reg __394714_394714;
   reg _394715_394715 ; 
   reg __394715_394715;
   reg _394716_394716 ; 
   reg __394716_394716;
   reg _394717_394717 ; 
   reg __394717_394717;
   reg _394718_394718 ; 
   reg __394718_394718;
   reg _394719_394719 ; 
   reg __394719_394719;
   reg _394720_394720 ; 
   reg __394720_394720;
   reg _394721_394721 ; 
   reg __394721_394721;
   reg _394722_394722 ; 
   reg __394722_394722;
   reg _394723_394723 ; 
   reg __394723_394723;
   reg _394724_394724 ; 
   reg __394724_394724;
   reg _394725_394725 ; 
   reg __394725_394725;
   reg _394726_394726 ; 
   reg __394726_394726;
   reg _394727_394727 ; 
   reg __394727_394727;
   reg _394728_394728 ; 
   reg __394728_394728;
   reg _394729_394729 ; 
   reg __394729_394729;
   reg _394730_394730 ; 
   reg __394730_394730;
   reg _394731_394731 ; 
   reg __394731_394731;
   reg _394732_394732 ; 
   reg __394732_394732;
   reg _394733_394733 ; 
   reg __394733_394733;
   reg _394734_394734 ; 
   reg __394734_394734;
   reg _394735_394735 ; 
   reg __394735_394735;
   reg _394736_394736 ; 
   reg __394736_394736;
   reg _394737_394737 ; 
   reg __394737_394737;
   reg _394738_394738 ; 
   reg __394738_394738;
   reg _394739_394739 ; 
   reg __394739_394739;
   reg _394740_394740 ; 
   reg __394740_394740;
   reg _394741_394741 ; 
   reg __394741_394741;
   reg _394742_394742 ; 
   reg __394742_394742;
   reg _394743_394743 ; 
   reg __394743_394743;
   reg _394744_394744 ; 
   reg __394744_394744;
   reg _394745_394745 ; 
   reg __394745_394745;
   reg _394746_394746 ; 
   reg __394746_394746;
   reg _394747_394747 ; 
   reg __394747_394747;
   reg _394748_394748 ; 
   reg __394748_394748;
   reg _394749_394749 ; 
   reg __394749_394749;
   reg _394750_394750 ; 
   reg __394750_394750;
   reg _394751_394751 ; 
   reg __394751_394751;
   reg _394752_394752 ; 
   reg __394752_394752;
   reg _394753_394753 ; 
   reg __394753_394753;
   reg _394754_394754 ; 
   reg __394754_394754;
   reg _394755_394755 ; 
   reg __394755_394755;
   reg _394756_394756 ; 
   reg __394756_394756;
   reg _394757_394757 ; 
   reg __394757_394757;
   reg _394758_394758 ; 
   reg __394758_394758;
   reg _394759_394759 ; 
   reg __394759_394759;
   reg _394760_394760 ; 
   reg __394760_394760;
   reg _394761_394761 ; 
   reg __394761_394761;
   reg _394762_394762 ; 
   reg __394762_394762;
   reg _394763_394763 ; 
   reg __394763_394763;
   reg _394764_394764 ; 
   reg __394764_394764;
   reg _394765_394765 ; 
   reg __394765_394765;
   reg _394766_394766 ; 
   reg __394766_394766;
   reg _394767_394767 ; 
   reg __394767_394767;
   reg _394768_394768 ; 
   reg __394768_394768;
   reg _394769_394769 ; 
   reg __394769_394769;
   reg _394770_394770 ; 
   reg __394770_394770;
   reg _394771_394771 ; 
   reg __394771_394771;
   reg _394772_394772 ; 
   reg __394772_394772;
   reg _394773_394773 ; 
   reg __394773_394773;
   reg _394774_394774 ; 
   reg __394774_394774;
   reg _394775_394775 ; 
   reg __394775_394775;
   reg _394776_394776 ; 
   reg __394776_394776;
   reg _394777_394777 ; 
   reg __394777_394777;
   reg _394778_394778 ; 
   reg __394778_394778;
   reg _394779_394779 ; 
   reg __394779_394779;
   reg _394780_394780 ; 
   reg __394780_394780;
   reg _394781_394781 ; 
   reg __394781_394781;
   reg _394782_394782 ; 
   reg __394782_394782;
   reg _394783_394783 ; 
   reg __394783_394783;
   reg _394784_394784 ; 
   reg __394784_394784;
   reg _394785_394785 ; 
   reg __394785_394785;
   reg _394786_394786 ; 
   reg __394786_394786;
   reg _394787_394787 ; 
   reg __394787_394787;
   reg _394788_394788 ; 
   reg __394788_394788;
   reg _394789_394789 ; 
   reg __394789_394789;
   reg _394790_394790 ; 
   reg __394790_394790;
   reg _394791_394791 ; 
   reg __394791_394791;
   reg _394792_394792 ; 
   reg __394792_394792;
   reg _394793_394793 ; 
   reg __394793_394793;
   reg _394794_394794 ; 
   reg __394794_394794;
   reg _394795_394795 ; 
   reg __394795_394795;
   reg _394796_394796 ; 
   reg __394796_394796;
   reg _394797_394797 ; 
   reg __394797_394797;
   reg _394798_394798 ; 
   reg __394798_394798;
   reg _394799_394799 ; 
   reg __394799_394799;
   reg _394800_394800 ; 
   reg __394800_394800;
   reg _394801_394801 ; 
   reg __394801_394801;
   reg _394802_394802 ; 
   reg __394802_394802;
   reg _394803_394803 ; 
   reg __394803_394803;
   reg _394804_394804 ; 
   reg __394804_394804;
   reg _394805_394805 ; 
   reg __394805_394805;
   reg _394806_394806 ; 
   reg __394806_394806;
   reg _394807_394807 ; 
   reg __394807_394807;
   reg _394808_394808 ; 
   reg __394808_394808;
   reg _394809_394809 ; 
   reg __394809_394809;
   reg _394810_394810 ; 
   reg __394810_394810;
   reg _394811_394811 ; 
   reg __394811_394811;
   reg _394812_394812 ; 
   reg __394812_394812;
   reg _394813_394813 ; 
   reg __394813_394813;
   reg _394814_394814 ; 
   reg __394814_394814;
   reg _394815_394815 ; 
   reg __394815_394815;
   reg _394816_394816 ; 
   reg __394816_394816;
   reg _394817_394817 ; 
   reg __394817_394817;
   reg _394818_394818 ; 
   reg __394818_394818;
   reg _394819_394819 ; 
   reg __394819_394819;
   reg _394820_394820 ; 
   reg __394820_394820;
   reg _394821_394821 ; 
   reg __394821_394821;
   reg _394822_394822 ; 
   reg __394822_394822;
   reg _394823_394823 ; 
   reg __394823_394823;
   reg _394824_394824 ; 
   reg __394824_394824;
   reg _394825_394825 ; 
   reg __394825_394825;
   reg _394826_394826 ; 
   reg __394826_394826;
   reg _394827_394827 ; 
   reg __394827_394827;
   reg _394828_394828 ; 
   reg __394828_394828;
   reg _394829_394829 ; 
   reg __394829_394829;
   reg _394830_394830 ; 
   reg __394830_394830;
   reg _394831_394831 ; 
   reg __394831_394831;
   reg _394832_394832 ; 
   reg __394832_394832;
   reg _394833_394833 ; 
   reg __394833_394833;
   reg _394834_394834 ; 
   reg __394834_394834;
   reg _394835_394835 ; 
   reg __394835_394835;
   reg _394836_394836 ; 
   reg __394836_394836;
   reg _394837_394837 ; 
   reg __394837_394837;
   reg _394838_394838 ; 
   reg __394838_394838;
   reg _394839_394839 ; 
   reg __394839_394839;
   reg _394840_394840 ; 
   reg __394840_394840;
   reg _394841_394841 ; 
   reg __394841_394841;
   reg _394842_394842 ; 
   reg __394842_394842;
   reg _394843_394843 ; 
   reg __394843_394843;
   reg _394844_394844 ; 
   reg __394844_394844;
   reg _394845_394845 ; 
   reg __394845_394845;
   reg _394846_394846 ; 
   reg __394846_394846;
   reg _394847_394847 ; 
   reg __394847_394847;
   reg _394848_394848 ; 
   reg __394848_394848;
   reg _394849_394849 ; 
   reg __394849_394849;
   reg _394850_394850 ; 
   reg __394850_394850;
   reg _394851_394851 ; 
   reg __394851_394851;
   reg _394852_394852 ; 
   reg __394852_394852;
   reg _394853_394853 ; 
   reg __394853_394853;
   reg _394854_394854 ; 
   reg __394854_394854;
   reg _394855_394855 ; 
   reg __394855_394855;
   reg _394856_394856 ; 
   reg __394856_394856;
   reg _394857_394857 ; 
   reg __394857_394857;
   reg _394858_394858 ; 
   reg __394858_394858;
   reg _394859_394859 ; 
   reg __394859_394859;
   reg _394860_394860 ; 
   reg __394860_394860;
   reg _394861_394861 ; 
   reg __394861_394861;
   reg _394862_394862 ; 
   reg __394862_394862;
   reg _394863_394863 ; 
   reg __394863_394863;
   reg _394864_394864 ; 
   reg __394864_394864;
   reg _394865_394865 ; 
   reg __394865_394865;
   reg _394866_394866 ; 
   reg __394866_394866;
   reg _394867_394867 ; 
   reg __394867_394867;
   reg _394868_394868 ; 
   reg __394868_394868;
   reg _394869_394869 ; 
   reg __394869_394869;
   reg _394870_394870 ; 
   reg __394870_394870;
   reg _394871_394871 ; 
   reg __394871_394871;
   reg _394872_394872 ; 
   reg __394872_394872;
   reg _394873_394873 ; 
   reg __394873_394873;
   reg _394874_394874 ; 
   reg __394874_394874;
   reg _394875_394875 ; 
   reg __394875_394875;
   reg _394876_394876 ; 
   reg __394876_394876;
   reg _394877_394877 ; 
   reg __394877_394877;
   reg _394878_394878 ; 
   reg __394878_394878;
   reg _394879_394879 ; 
   reg __394879_394879;
   reg _394880_394880 ; 
   reg __394880_394880;
   reg _394881_394881 ; 
   reg __394881_394881;
   reg _394882_394882 ; 
   reg __394882_394882;
   reg _394883_394883 ; 
   reg __394883_394883;
   reg _394884_394884 ; 
   reg __394884_394884;
   reg _394885_394885 ; 
   reg __394885_394885;
   reg _394886_394886 ; 
   reg __394886_394886;
   reg _394887_394887 ; 
   reg __394887_394887;
   reg _394888_394888 ; 
   reg __394888_394888;
   reg _394889_394889 ; 
   reg __394889_394889;
   reg _394890_394890 ; 
   reg __394890_394890;
   reg _394891_394891 ; 
   reg __394891_394891;
   reg _394892_394892 ; 
   reg __394892_394892;
   reg _394893_394893 ; 
   reg __394893_394893;
   reg _394894_394894 ; 
   reg __394894_394894;
   reg _394895_394895 ; 
   reg __394895_394895;
   reg _394896_394896 ; 
   reg __394896_394896;
   reg _394897_394897 ; 
   reg __394897_394897;
   reg _394898_394898 ; 
   reg __394898_394898;
   reg _394899_394899 ; 
   reg __394899_394899;
   reg _394900_394900 ; 
   reg __394900_394900;
   reg _394901_394901 ; 
   reg __394901_394901;
   reg _394902_394902 ; 
   reg __394902_394902;
   reg _394903_394903 ; 
   reg __394903_394903;
   reg _394904_394904 ; 
   reg __394904_394904;
   reg _394905_394905 ; 
   reg __394905_394905;
   reg _394906_394906 ; 
   reg __394906_394906;
   reg _394907_394907 ; 
   reg __394907_394907;
   reg _394908_394908 ; 
   reg __394908_394908;
   reg _394909_394909 ; 
   reg __394909_394909;
   reg _394910_394910 ; 
   reg __394910_394910;
   reg _394911_394911 ; 
   reg __394911_394911;
   reg _394912_394912 ; 
   reg __394912_394912;
   reg _394913_394913 ; 
   reg __394913_394913;
   reg _394914_394914 ; 
   reg __394914_394914;
   reg _394915_394915 ; 
   reg __394915_394915;
   reg _394916_394916 ; 
   reg __394916_394916;
   reg _394917_394917 ; 
   reg __394917_394917;
   reg _394918_394918 ; 
   reg __394918_394918;
   reg _394919_394919 ; 
   reg __394919_394919;
   reg _394920_394920 ; 
   reg __394920_394920;
   reg _394921_394921 ; 
   reg __394921_394921;
   reg _394922_394922 ; 
   reg __394922_394922;
   reg _394923_394923 ; 
   reg __394923_394923;
   reg _394924_394924 ; 
   reg __394924_394924;
   reg _394925_394925 ; 
   reg __394925_394925;
   reg _394926_394926 ; 
   reg __394926_394926;
   reg _394927_394927 ; 
   reg __394927_394927;
   reg _394928_394928 ; 
   reg __394928_394928;
   reg _394929_394929 ; 
   reg __394929_394929;
   reg _394930_394930 ; 
   reg __394930_394930;
   reg _394931_394931 ; 
   reg __394931_394931;
   reg _394932_394932 ; 
   reg __394932_394932;
   reg _394933_394933 ; 
   reg __394933_394933;
   reg _394934_394934 ; 
   reg __394934_394934;
   reg _394935_394935 ; 
   reg __394935_394935;
   reg _394936_394936 ; 
   reg __394936_394936;
   reg _394937_394937 ; 
   reg __394937_394937;
   reg _394938_394938 ; 
   reg __394938_394938;
   reg _394939_394939 ; 
   reg __394939_394939;
   reg _394940_394940 ; 
   reg __394940_394940;
   reg _394941_394941 ; 
   reg __394941_394941;
   reg _394942_394942 ; 
   reg __394942_394942;
   reg _394943_394943 ; 
   reg __394943_394943;
   reg _394944_394944 ; 
   reg __394944_394944;
   reg _394945_394945 ; 
   reg __394945_394945;
   reg _394946_394946 ; 
   reg __394946_394946;
   reg _394947_394947 ; 
   reg __394947_394947;
   reg _394948_394948 ; 
   reg __394948_394948;
   reg _394949_394949 ; 
   reg __394949_394949;
   reg _394950_394950 ; 
   reg __394950_394950;
   reg _394951_394951 ; 
   reg __394951_394951;
   reg _394952_394952 ; 
   reg __394952_394952;
   reg _394953_394953 ; 
   reg __394953_394953;
   reg _394954_394954 ; 
   reg __394954_394954;
   reg _394955_394955 ; 
   reg __394955_394955;
   reg _394956_394956 ; 
   reg __394956_394956;
   reg _394957_394957 ; 
   reg __394957_394957;
   reg _394958_394958 ; 
   reg __394958_394958;
   reg _394959_394959 ; 
   reg __394959_394959;
   reg _394960_394960 ; 
   reg __394960_394960;
   reg _394961_394961 ; 
   reg __394961_394961;
   reg _394962_394962 ; 
   reg __394962_394962;
   reg _394963_394963 ; 
   reg __394963_394963;
   reg _394964_394964 ; 
   reg __394964_394964;
   reg _394965_394965 ; 
   reg __394965_394965;
   reg _394966_394966 ; 
   reg __394966_394966;
   reg _394967_394967 ; 
   reg __394967_394967;
   reg _394968_394968 ; 
   reg __394968_394968;
   reg _394969_394969 ; 
   reg __394969_394969;
   reg _394970_394970 ; 
   reg __394970_394970;
   reg _394971_394971 ; 
   reg __394971_394971;
   reg _394972_394972 ; 
   reg __394972_394972;
   reg _394973_394973 ; 
   reg __394973_394973;
   reg _394974_394974 ; 
   reg __394974_394974;
   reg _394975_394975 ; 
   reg __394975_394975;
   reg _394976_394976 ; 
   reg __394976_394976;
   reg _394977_394977 ; 
   reg __394977_394977;
   reg _394978_394978 ; 
   reg __394978_394978;
   reg _394979_394979 ; 
   reg __394979_394979;
   reg _394980_394980 ; 
   reg __394980_394980;
   reg _394981_394981 ; 
   reg __394981_394981;
   reg _394982_394982 ; 
   reg __394982_394982;
   reg _394983_394983 ; 
   reg __394983_394983;
   reg _394984_394984 ; 
   reg __394984_394984;
   reg _394985_394985 ; 
   reg __394985_394985;
   reg _394986_394986 ; 
   reg __394986_394986;
   reg _394987_394987 ; 
   reg __394987_394987;
   reg _394988_394988 ; 
   reg __394988_394988;
   reg _394989_394989 ; 
   reg __394989_394989;
   reg _394990_394990 ; 
   reg __394990_394990;
   reg _394991_394991 ; 
   reg __394991_394991;
   reg _394992_394992 ; 
   reg __394992_394992;
   reg _394993_394993 ; 
   reg __394993_394993;
   reg _394994_394994 ; 
   reg __394994_394994;
   reg _394995_394995 ; 
   reg __394995_394995;
   reg _394996_394996 ; 
   reg __394996_394996;
   reg _394997_394997 ; 
   reg __394997_394997;
   reg _394998_394998 ; 
   reg __394998_394998;
   reg _394999_394999 ; 
   reg __394999_394999;
   reg _395000_395000 ; 
   reg __395000_395000;
   reg _395001_395001 ; 
   reg __395001_395001;
   reg _395002_395002 ; 
   reg __395002_395002;
   reg _395003_395003 ; 
   reg __395003_395003;
   reg _395004_395004 ; 
   reg __395004_395004;
   reg _395005_395005 ; 
   reg __395005_395005;
   reg _395006_395006 ; 
   reg __395006_395006;
   reg _395007_395007 ; 
   reg __395007_395007;
   reg _395008_395008 ; 
   reg __395008_395008;
   reg _395009_395009 ; 
   reg __395009_395009;
   reg _395010_395010 ; 
   reg __395010_395010;
   reg _395011_395011 ; 
   reg __395011_395011;
   reg _395012_395012 ; 
   reg __395012_395012;
   reg _395013_395013 ; 
   reg __395013_395013;
   reg _395014_395014 ; 
   reg __395014_395014;
   reg _395015_395015 ; 
   reg __395015_395015;
   reg _395016_395016 ; 
   reg __395016_395016;
   reg _395017_395017 ; 
   reg __395017_395017;
   reg _395018_395018 ; 
   reg __395018_395018;
   reg _395019_395019 ; 
   reg __395019_395019;
   reg _395020_395020 ; 
   reg __395020_395020;
   reg _395021_395021 ; 
   reg __395021_395021;
   reg _395022_395022 ; 
   reg __395022_395022;
   reg _395023_395023 ; 
   reg __395023_395023;
   reg _395024_395024 ; 
   reg __395024_395024;
   reg _395025_395025 ; 
   reg __395025_395025;
   reg _395026_395026 ; 
   reg __395026_395026;
   reg _395027_395027 ; 
   reg __395027_395027;
   reg _395028_395028 ; 
   reg __395028_395028;
   reg _395029_395029 ; 
   reg __395029_395029;
   reg _395030_395030 ; 
   reg __395030_395030;
   reg _395031_395031 ; 
   reg __395031_395031;
   reg _395032_395032 ; 
   reg __395032_395032;
   reg _395033_395033 ; 
   reg __395033_395033;
   reg _395034_395034 ; 
   reg __395034_395034;
   reg _395035_395035 ; 
   reg __395035_395035;
   reg _395036_395036 ; 
   reg __395036_395036;
   reg _395037_395037 ; 
   reg __395037_395037;
   reg _395038_395038 ; 
   reg __395038_395038;
   reg _395039_395039 ; 
   reg __395039_395039;
   reg _395040_395040 ; 
   reg __395040_395040;
   reg _395041_395041 ; 
   reg __395041_395041;
   reg _395042_395042 ; 
   reg __395042_395042;
   reg _395043_395043 ; 
   reg __395043_395043;
   reg _395044_395044 ; 
   reg __395044_395044;
   reg _395045_395045 ; 
   reg __395045_395045;
   reg _395046_395046 ; 
   reg __395046_395046;
   reg _395047_395047 ; 
   reg __395047_395047;
   reg _395048_395048 ; 
   reg __395048_395048;
   reg _395049_395049 ; 
   reg __395049_395049;
   reg _395050_395050 ; 
   reg __395050_395050;
   reg _395051_395051 ; 
   reg __395051_395051;
   reg _395052_395052 ; 
   reg __395052_395052;
   reg _395053_395053 ; 
   reg __395053_395053;
   reg _395054_395054 ; 
   reg __395054_395054;
   reg _395055_395055 ; 
   reg __395055_395055;
   reg _395056_395056 ; 
   reg __395056_395056;
   reg _395057_395057 ; 
   reg __395057_395057;
   reg _395058_395058 ; 
   reg __395058_395058;
   reg _395059_395059 ; 
   reg __395059_395059;
   reg _395060_395060 ; 
   reg __395060_395060;
   reg _395061_395061 ; 
   reg __395061_395061;
   reg _395062_395062 ; 
   reg __395062_395062;
   reg _395063_395063 ; 
   reg __395063_395063;
   reg _395064_395064 ; 
   reg __395064_395064;
   reg _395065_395065 ; 
   reg __395065_395065;
   reg _395066_395066 ; 
   reg __395066_395066;
   reg _395067_395067 ; 
   reg __395067_395067;
   reg _395068_395068 ; 
   reg __395068_395068;
   reg _395069_395069 ; 
   reg __395069_395069;
   reg _395070_395070 ; 
   reg __395070_395070;
   reg _395071_395071 ; 
   reg __395071_395071;
   reg _395072_395072 ; 
   reg __395072_395072;
   reg _395073_395073 ; 
   reg __395073_395073;
   reg _395074_395074 ; 
   reg __395074_395074;
   reg _395075_395075 ; 
   reg __395075_395075;
   reg _395076_395076 ; 
   reg __395076_395076;
   reg _395077_395077 ; 
   reg __395077_395077;
   reg _395078_395078 ; 
   reg __395078_395078;
   reg _395079_395079 ; 
   reg __395079_395079;
   reg _395080_395080 ; 
   reg __395080_395080;
   reg _395081_395081 ; 
   reg __395081_395081;
   reg _395082_395082 ; 
   reg __395082_395082;
   reg _395083_395083 ; 
   reg __395083_395083;
   reg _395084_395084 ; 
   reg __395084_395084;
   reg _395085_395085 ; 
   reg __395085_395085;
   reg _395086_395086 ; 
   reg __395086_395086;
   reg _395087_395087 ; 
   reg __395087_395087;
   reg _395088_395088 ; 
   reg __395088_395088;
   reg _395089_395089 ; 
   reg __395089_395089;
   reg _395090_395090 ; 
   reg __395090_395090;
   reg _395091_395091 ; 
   reg __395091_395091;
   reg _395092_395092 ; 
   reg __395092_395092;
   reg _395093_395093 ; 
   reg __395093_395093;
   reg _395094_395094 ; 
   reg __395094_395094;
   reg _395095_395095 ; 
   reg __395095_395095;
   reg _395096_395096 ; 
   reg __395096_395096;
   reg _395097_395097 ; 
   reg __395097_395097;
   reg _395098_395098 ; 
   reg __395098_395098;
   reg _395099_395099 ; 
   reg __395099_395099;
   reg _395100_395100 ; 
   reg __395100_395100;
   reg _395101_395101 ; 
   reg __395101_395101;
   reg _395102_395102 ; 
   reg __395102_395102;
   reg _395103_395103 ; 
   reg __395103_395103;
   reg _395104_395104 ; 
   reg __395104_395104;
   reg _395105_395105 ; 
   reg __395105_395105;
   reg _395106_395106 ; 
   reg __395106_395106;
   reg _395107_395107 ; 
   reg __395107_395107;
   reg _395108_395108 ; 
   reg __395108_395108;
   reg _395109_395109 ; 
   reg __395109_395109;
   reg _395110_395110 ; 
   reg __395110_395110;
   reg _395111_395111 ; 
   reg __395111_395111;
   reg _395112_395112 ; 
   reg __395112_395112;
   reg _395113_395113 ; 
   reg __395113_395113;
   reg _395114_395114 ; 
   reg __395114_395114;
   reg _395115_395115 ; 
   reg __395115_395115;
   reg _395116_395116 ; 
   reg __395116_395116;
   reg _395117_395117 ; 
   reg __395117_395117;
   reg _395118_395118 ; 
   reg __395118_395118;
   reg _395119_395119 ; 
   reg __395119_395119;
   reg _395120_395120 ; 
   reg __395120_395120;
   reg _395121_395121 ; 
   reg __395121_395121;
   reg _395122_395122 ; 
   reg __395122_395122;
   reg _395123_395123 ; 
   reg __395123_395123;
   reg _395124_395124 ; 
   reg __395124_395124;
   reg _395125_395125 ; 
   reg __395125_395125;
   reg _395126_395126 ; 
   reg __395126_395126;
   reg _395127_395127 ; 
   reg __395127_395127;
   reg _395128_395128 ; 
   reg __395128_395128;
   reg _395129_395129 ; 
   reg __395129_395129;
   reg _395130_395130 ; 
   reg __395130_395130;
   reg _395131_395131 ; 
   reg __395131_395131;
   reg _395132_395132 ; 
   reg __395132_395132;
   reg _395133_395133 ; 
   reg __395133_395133;
   reg _395134_395134 ; 
   reg __395134_395134;
   reg _395135_395135 ; 
   reg __395135_395135;
   reg _395136_395136 ; 
   reg __395136_395136;
   reg _395137_395137 ; 
   reg __395137_395137;
   reg _395138_395138 ; 
   reg __395138_395138;
   reg _395139_395139 ; 
   reg __395139_395139;
   reg _395140_395140 ; 
   reg __395140_395140;
   reg _395141_395141 ; 
   reg __395141_395141;
   reg _395142_395142 ; 
   reg __395142_395142;
   reg _395143_395143 ; 
   reg __395143_395143;
   reg _395144_395144 ; 
   reg __395144_395144;
   reg _395145_395145 ; 
   reg __395145_395145;
   reg _395146_395146 ; 
   reg __395146_395146;
   reg _395147_395147 ; 
   reg __395147_395147;
   reg _395148_395148 ; 
   reg __395148_395148;
   reg _395149_395149 ; 
   reg __395149_395149;
   reg _395150_395150 ; 
   reg __395150_395150;
   reg _395151_395151 ; 
   reg __395151_395151;
   reg _395152_395152 ; 
   reg __395152_395152;
   reg _395153_395153 ; 
   reg __395153_395153;
   reg _395154_395154 ; 
   reg __395154_395154;
   reg _395155_395155 ; 
   reg __395155_395155;
   reg _395156_395156 ; 
   reg __395156_395156;
   reg _395157_395157 ; 
   reg __395157_395157;
   reg _395158_395158 ; 
   reg __395158_395158;
   reg _395159_395159 ; 
   reg __395159_395159;
   reg _395160_395160 ; 
   reg __395160_395160;
   reg _395161_395161 ; 
   reg __395161_395161;
   reg _395162_395162 ; 
   reg __395162_395162;
   reg _395163_395163 ; 
   reg __395163_395163;
   reg _395164_395164 ; 
   reg __395164_395164;
   reg _395165_395165 ; 
   reg __395165_395165;
   reg _395166_395166 ; 
   reg __395166_395166;
   reg _395167_395167 ; 
   reg __395167_395167;
   reg _395168_395168 ; 
   reg __395168_395168;
   reg _395169_395169 ; 
   reg __395169_395169;
   reg _395170_395170 ; 
   reg __395170_395170;
   reg _395171_395171 ; 
   reg __395171_395171;
   reg _395172_395172 ; 
   reg __395172_395172;
   reg _395173_395173 ; 
   reg __395173_395173;
   reg _395174_395174 ; 
   reg __395174_395174;
   reg _395175_395175 ; 
   reg __395175_395175;
   reg _395176_395176 ; 
   reg __395176_395176;
   reg _395177_395177 ; 
   reg __395177_395177;
   reg _395178_395178 ; 
   reg __395178_395178;
   reg _395179_395179 ; 
   reg __395179_395179;
   reg _395180_395180 ; 
   reg __395180_395180;
   reg _395181_395181 ; 
   reg __395181_395181;
   reg _395182_395182 ; 
   reg __395182_395182;
   reg _395183_395183 ; 
   reg __395183_395183;
   reg _395184_395184 ; 
   reg __395184_395184;
   reg _395185_395185 ; 
   reg __395185_395185;
   reg _395186_395186 ; 
   reg __395186_395186;
   reg _395187_395187 ; 
   reg __395187_395187;
   reg _395188_395188 ; 
   reg __395188_395188;
   reg _395189_395189 ; 
   reg __395189_395189;
   reg _395190_395190 ; 
   reg __395190_395190;
   reg _395191_395191 ; 
   reg __395191_395191;
   reg _395192_395192 ; 
   reg __395192_395192;
   reg _395193_395193 ; 
   reg __395193_395193;
   reg _395194_395194 ; 
   reg __395194_395194;
   reg _395195_395195 ; 
   reg __395195_395195;
   reg _395196_395196 ; 
   reg __395196_395196;
   reg _395197_395197 ; 
   reg __395197_395197;
   reg _395198_395198 ; 
   reg __395198_395198;
   reg _395199_395199 ; 
   reg __395199_395199;
   reg _395200_395200 ; 
   reg __395200_395200;
   reg _395201_395201 ; 
   reg __395201_395201;
   reg _395202_395202 ; 
   reg __395202_395202;
   reg _395203_395203 ; 
   reg __395203_395203;
   reg _395204_395204 ; 
   reg __395204_395204;
   reg _395205_395205 ; 
   reg __395205_395205;
   reg _395206_395206 ; 
   reg __395206_395206;
   reg _395207_395207 ; 
   reg __395207_395207;
   reg _395208_395208 ; 
   reg __395208_395208;
   reg _395209_395209 ; 
   reg __395209_395209;
   reg _395210_395210 ; 
   reg __395210_395210;
   reg _395211_395211 ; 
   reg __395211_395211;
   reg _395212_395212 ; 
   reg __395212_395212;
   reg _395213_395213 ; 
   reg __395213_395213;
   reg _395214_395214 ; 
   reg __395214_395214;
   reg _395215_395215 ; 
   reg __395215_395215;
   reg _395216_395216 ; 
   reg __395216_395216;
   reg _395217_395217 ; 
   reg __395217_395217;
   reg _395218_395218 ; 
   reg __395218_395218;
   reg _395219_395219 ; 
   reg __395219_395219;
   reg _395220_395220 ; 
   reg __395220_395220;
   reg _395221_395221 ; 
   reg __395221_395221;
   reg _395222_395222 ; 
   reg __395222_395222;
   reg _395223_395223 ; 
   reg __395223_395223;
   reg _395224_395224 ; 
   reg __395224_395224;
   reg _395225_395225 ; 
   reg __395225_395225;
   reg _395226_395226 ; 
   reg __395226_395226;
   reg _395227_395227 ; 
   reg __395227_395227;
   reg _395228_395228 ; 
   reg __395228_395228;
   reg _395229_395229 ; 
   reg __395229_395229;
   reg _395230_395230 ; 
   reg __395230_395230;
   reg _395231_395231 ; 
   reg __395231_395231;
   reg _395232_395232 ; 
   reg __395232_395232;
   reg _395233_395233 ; 
   reg __395233_395233;
   reg _395234_395234 ; 
   reg __395234_395234;
   reg _395235_395235 ; 
   reg __395235_395235;
   reg _395236_395236 ; 
   reg __395236_395236;
   reg _395237_395237 ; 
   reg __395237_395237;
   reg _395238_395238 ; 
   reg __395238_395238;
   reg _395239_395239 ; 
   reg __395239_395239;
   reg _395240_395240 ; 
   reg __395240_395240;
   reg _395241_395241 ; 
   reg __395241_395241;
   reg _395242_395242 ; 
   reg __395242_395242;
   reg _395243_395243 ; 
   reg __395243_395243;
   reg _395244_395244 ; 
   reg __395244_395244;
   reg _395245_395245 ; 
   reg __395245_395245;
   reg _395246_395246 ; 
   reg __395246_395246;
   reg _395247_395247 ; 
   reg __395247_395247;
   reg _395248_395248 ; 
   reg __395248_395248;
   reg _395249_395249 ; 
   reg __395249_395249;
   reg _395250_395250 ; 
   reg __395250_395250;
   reg _395251_395251 ; 
   reg __395251_395251;
   reg _395252_395252 ; 
   reg __395252_395252;
   reg _395253_395253 ; 
   reg __395253_395253;
   reg _395254_395254 ; 
   reg __395254_395254;
   reg _395255_395255 ; 
   reg __395255_395255;
   reg _395256_395256 ; 
   reg __395256_395256;
   reg _395257_395257 ; 
   reg __395257_395257;
   reg _395258_395258 ; 
   reg __395258_395258;
   reg _395259_395259 ; 
   reg __395259_395259;
   reg _395260_395260 ; 
   reg __395260_395260;
   reg _395261_395261 ; 
   reg __395261_395261;
   reg _395262_395262 ; 
   reg __395262_395262;
   reg _395263_395263 ; 
   reg __395263_395263;
   reg _395264_395264 ; 
   reg __395264_395264;
   reg _395265_395265 ; 
   reg __395265_395265;
   reg _395266_395266 ; 
   reg __395266_395266;
   reg _395267_395267 ; 
   reg __395267_395267;
   reg _395268_395268 ; 
   reg __395268_395268;
   reg _395269_395269 ; 
   reg __395269_395269;
   reg _395270_395270 ; 
   reg __395270_395270;
   reg _395271_395271 ; 
   reg __395271_395271;
   reg _395272_395272 ; 
   reg __395272_395272;
   reg _395273_395273 ; 
   reg __395273_395273;
   reg _395274_395274 ; 
   reg __395274_395274;
   reg _395275_395275 ; 
   reg __395275_395275;
   reg _395276_395276 ; 
   reg __395276_395276;
   reg _395277_395277 ; 
   reg __395277_395277;
   reg _395278_395278 ; 
   reg __395278_395278;
   reg _395279_395279 ; 
   reg __395279_395279;
   reg _395280_395280 ; 
   reg __395280_395280;
   reg _395281_395281 ; 
   reg __395281_395281;
   reg _395282_395282 ; 
   reg __395282_395282;
   reg _395283_395283 ; 
   reg __395283_395283;
   reg _395284_395284 ; 
   reg __395284_395284;
   reg _395285_395285 ; 
   reg __395285_395285;
   reg _395286_395286 ; 
   reg __395286_395286;
   reg _395287_395287 ; 
   reg __395287_395287;
   reg _395288_395288 ; 
   reg __395288_395288;
   reg _395289_395289 ; 
   reg __395289_395289;
   reg _395290_395290 ; 
   reg __395290_395290;
   reg _395291_395291 ; 
   reg __395291_395291;
   reg _395292_395292 ; 
   reg __395292_395292;
   reg _395293_395293 ; 
   reg __395293_395293;
   reg _395294_395294 ; 
   reg __395294_395294;
   reg _395295_395295 ; 
   reg __395295_395295;
   reg _395296_395296 ; 
   reg __395296_395296;
   reg _395297_395297 ; 
   reg __395297_395297;
   reg _395298_395298 ; 
   reg __395298_395298;
   reg _395299_395299 ; 
   reg __395299_395299;
   reg _395300_395300 ; 
   reg __395300_395300;
   reg _395301_395301 ; 
   reg __395301_395301;
   reg _395302_395302 ; 
   reg __395302_395302;
   reg _395303_395303 ; 
   reg __395303_395303;
   reg _395304_395304 ; 
   reg __395304_395304;
   reg _395305_395305 ; 
   reg __395305_395305;
   reg _395306_395306 ; 
   reg __395306_395306;
   reg _395307_395307 ; 
   reg __395307_395307;
   reg _395308_395308 ; 
   reg __395308_395308;
   reg _395309_395309 ; 
   reg __395309_395309;
   reg _395310_395310 ; 
   reg __395310_395310;
   reg _395311_395311 ; 
   reg __395311_395311;
   reg _395312_395312 ; 
   reg __395312_395312;
   reg _395313_395313 ; 
   reg __395313_395313;
   reg _395314_395314 ; 
   reg __395314_395314;
   reg _395315_395315 ; 
   reg __395315_395315;
   reg _395316_395316 ; 
   reg __395316_395316;
   reg _395317_395317 ; 
   reg __395317_395317;
   reg _395318_395318 ; 
   reg __395318_395318;
   reg _395319_395319 ; 
   reg __395319_395319;
   reg _395320_395320 ; 
   reg __395320_395320;
   reg _395321_395321 ; 
   reg __395321_395321;
   reg _395322_395322 ; 
   reg __395322_395322;
   reg _395323_395323 ; 
   reg __395323_395323;
   reg _395324_395324 ; 
   reg __395324_395324;
   reg _395325_395325 ; 
   reg __395325_395325;
   reg _395326_395326 ; 
   reg __395326_395326;
   reg _395327_395327 ; 
   reg __395327_395327;
   reg _395328_395328 ; 
   reg __395328_395328;
   reg _395329_395329 ; 
   reg __395329_395329;
   reg _395330_395330 ; 
   reg __395330_395330;
   reg _395331_395331 ; 
   reg __395331_395331;
   reg _395332_395332 ; 
   reg __395332_395332;
   reg _395333_395333 ; 
   reg __395333_395333;
   reg _395334_395334 ; 
   reg __395334_395334;
   reg _395335_395335 ; 
   reg __395335_395335;
   reg _395336_395336 ; 
   reg __395336_395336;
   reg _395337_395337 ; 
   reg __395337_395337;
   reg _395338_395338 ; 
   reg __395338_395338;
   reg _395339_395339 ; 
   reg __395339_395339;
   reg _395340_395340 ; 
   reg __395340_395340;
   reg _395341_395341 ; 
   reg __395341_395341;
   reg _395342_395342 ; 
   reg __395342_395342;
   reg _395343_395343 ; 
   reg __395343_395343;
   reg _395344_395344 ; 
   reg __395344_395344;
   reg _395345_395345 ; 
   reg __395345_395345;
   reg _395346_395346 ; 
   reg __395346_395346;
   reg _395347_395347 ; 
   reg __395347_395347;
   reg _395348_395348 ; 
   reg __395348_395348;
   reg _395349_395349 ; 
   reg __395349_395349;
   reg _395350_395350 ; 
   reg __395350_395350;
   reg _395351_395351 ; 
   reg __395351_395351;
   reg _395352_395352 ; 
   reg __395352_395352;
   reg _395353_395353 ; 
   reg __395353_395353;
   reg _395354_395354 ; 
   reg __395354_395354;
   reg _395355_395355 ; 
   reg __395355_395355;
   reg _395356_395356 ; 
   reg __395356_395356;
   reg _395357_395357 ; 
   reg __395357_395357;
   reg _395358_395358 ; 
   reg __395358_395358;
   reg _395359_395359 ; 
   reg __395359_395359;
   reg _395360_395360 ; 
   reg __395360_395360;
   reg _395361_395361 ; 
   reg __395361_395361;
   reg _395362_395362 ; 
   reg __395362_395362;
   reg _395363_395363 ; 
   reg __395363_395363;
   reg _395364_395364 ; 
   reg __395364_395364;
   reg _395365_395365 ; 
   reg __395365_395365;
   reg _395366_395366 ; 
   reg __395366_395366;
   reg _395367_395367 ; 
   reg __395367_395367;
   reg _395368_395368 ; 
   reg __395368_395368;
   reg _395369_395369 ; 
   reg __395369_395369;
   reg _395370_395370 ; 
   reg __395370_395370;
   reg _395371_395371 ; 
   reg __395371_395371;
   reg _395372_395372 ; 
   reg __395372_395372;
   reg _395373_395373 ; 
   reg __395373_395373;
   reg _395374_395374 ; 
   reg __395374_395374;
   reg _395375_395375 ; 
   reg __395375_395375;
   reg _395376_395376 ; 
   reg __395376_395376;
   reg _395377_395377 ; 
   reg __395377_395377;
   reg _395378_395378 ; 
   reg __395378_395378;
   reg _395379_395379 ; 
   reg __395379_395379;
   reg _395380_395380 ; 
   reg __395380_395380;
   reg _395381_395381 ; 
   reg __395381_395381;
   reg _395382_395382 ; 
   reg __395382_395382;
   reg _395383_395383 ; 
   reg __395383_395383;
   reg _395384_395384 ; 
   reg __395384_395384;
   reg _395385_395385 ; 
   reg __395385_395385;
   reg _395386_395386 ; 
   reg __395386_395386;
   reg _395387_395387 ; 
   reg __395387_395387;
   reg _395388_395388 ; 
   reg __395388_395388;
   reg _395389_395389 ; 
   reg __395389_395389;
   reg _395390_395390 ; 
   reg __395390_395390;
   reg _395391_395391 ; 
   reg __395391_395391;
   reg _395392_395392 ; 
   reg __395392_395392;
   reg _395393_395393 ; 
   reg __395393_395393;
   reg _395394_395394 ; 
   reg __395394_395394;
   reg _395395_395395 ; 
   reg __395395_395395;
   reg _395396_395396 ; 
   reg __395396_395396;
   reg _395397_395397 ; 
   reg __395397_395397;
   reg _395398_395398 ; 
   reg __395398_395398;
   reg _395399_395399 ; 
   reg __395399_395399;
   reg _395400_395400 ; 
   reg __395400_395400;
   reg _395401_395401 ; 
   reg __395401_395401;
   reg _395402_395402 ; 
   reg __395402_395402;
   reg _395403_395403 ; 
   reg __395403_395403;
   reg _395404_395404 ; 
   reg __395404_395404;
   reg _395405_395405 ; 
   reg __395405_395405;
   reg _395406_395406 ; 
   reg __395406_395406;
   reg _395407_395407 ; 
   reg __395407_395407;
   reg _395408_395408 ; 
   reg __395408_395408;
   reg _395409_395409 ; 
   reg __395409_395409;
   reg _395410_395410 ; 
   reg __395410_395410;
   reg _395411_395411 ; 
   reg __395411_395411;
   reg _395412_395412 ; 
   reg __395412_395412;
   reg _395413_395413 ; 
   reg __395413_395413;
   reg _395414_395414 ; 
   reg __395414_395414;
   reg _395415_395415 ; 
   reg __395415_395415;
   reg _395416_395416 ; 
   reg __395416_395416;
   reg _395417_395417 ; 
   reg __395417_395417;
   reg _395418_395418 ; 
   reg __395418_395418;
   reg _395419_395419 ; 
   reg __395419_395419;
   reg _395420_395420 ; 
   reg __395420_395420;
   reg _395421_395421 ; 
   reg __395421_395421;
   reg _395422_395422 ; 
   reg __395422_395422;
   reg _395423_395423 ; 
   reg __395423_395423;
   reg _395424_395424 ; 
   reg __395424_395424;
   reg _395425_395425 ; 
   reg __395425_395425;
   reg _395426_395426 ; 
   reg __395426_395426;
   reg _395427_395427 ; 
   reg __395427_395427;
   reg _395428_395428 ; 
   reg __395428_395428;
   reg _395429_395429 ; 
   reg __395429_395429;
   reg _395430_395430 ; 
   reg __395430_395430;
   reg _395431_395431 ; 
   reg __395431_395431;
   reg _395432_395432 ; 
   reg __395432_395432;
   reg _395433_395433 ; 
   reg __395433_395433;
   reg _395434_395434 ; 
   reg __395434_395434;
   reg _395435_395435 ; 
   reg __395435_395435;
   reg _395436_395436 ; 
   reg __395436_395436;
   reg _395437_395437 ; 
   reg __395437_395437;
   reg _395438_395438 ; 
   reg __395438_395438;
   reg _395439_395439 ; 
   reg __395439_395439;
   reg _395440_395440 ; 
   reg __395440_395440;
   reg _395441_395441 ; 
   reg __395441_395441;
   reg _395442_395442 ; 
   reg __395442_395442;
   reg _395443_395443 ; 
   reg __395443_395443;
   reg _395444_395444 ; 
   reg __395444_395444;
   reg _395445_395445 ; 
   reg __395445_395445;
   reg _395446_395446 ; 
   reg __395446_395446;
   reg _395447_395447 ; 
   reg __395447_395447;
   reg _395448_395448 ; 
   reg __395448_395448;
   reg _395449_395449 ; 
   reg __395449_395449;
   reg _395450_395450 ; 
   reg __395450_395450;
   reg _395451_395451 ; 
   reg __395451_395451;
   reg _395452_395452 ; 
   reg __395452_395452;
   reg _395453_395453 ; 
   reg __395453_395453;
   reg _395454_395454 ; 
   reg __395454_395454;
   reg _395455_395455 ; 
   reg __395455_395455;
   reg _395456_395456 ; 
   reg __395456_395456;
   reg _395457_395457 ; 
   reg __395457_395457;
   reg _395458_395458 ; 
   reg __395458_395458;
   reg _395459_395459 ; 
   reg __395459_395459;
   reg _395460_395460 ; 
   reg __395460_395460;
   reg _395461_395461 ; 
   reg __395461_395461;
   reg _395462_395462 ; 
   reg __395462_395462;
   reg _395463_395463 ; 
   reg __395463_395463;
   reg _395464_395464 ; 
   reg __395464_395464;
   reg _395465_395465 ; 
   reg __395465_395465;
   reg _395466_395466 ; 
   reg __395466_395466;
   reg _395467_395467 ; 
   reg __395467_395467;
   reg _395468_395468 ; 
   reg __395468_395468;
   reg _395469_395469 ; 
   reg __395469_395469;
   reg _395470_395470 ; 
   reg __395470_395470;
   reg _395471_395471 ; 
   reg __395471_395471;
   reg _395472_395472 ; 
   reg __395472_395472;
   reg _395473_395473 ; 
   reg __395473_395473;
   reg _395474_395474 ; 
   reg __395474_395474;
   reg _395475_395475 ; 
   reg __395475_395475;
   reg _395476_395476 ; 
   reg __395476_395476;
   reg _395477_395477 ; 
   reg __395477_395477;
   reg _395478_395478 ; 
   reg __395478_395478;
   reg _395479_395479 ; 
   reg __395479_395479;
   reg _395480_395480 ; 
   reg __395480_395480;
   reg _395481_395481 ; 
   reg __395481_395481;
   reg _395482_395482 ; 
   reg __395482_395482;
   reg _395483_395483 ; 
   reg __395483_395483;
   reg _395484_395484 ; 
   reg __395484_395484;
   reg _395485_395485 ; 
   reg __395485_395485;
   reg _395486_395486 ; 
   reg __395486_395486;
   reg _395487_395487 ; 
   reg __395487_395487;
   reg _395488_395488 ; 
   reg __395488_395488;
   reg _395489_395489 ; 
   reg __395489_395489;
   reg _395490_395490 ; 
   reg __395490_395490;
   reg _395491_395491 ; 
   reg __395491_395491;
   reg _395492_395492 ; 
   reg __395492_395492;
   reg _395493_395493 ; 
   reg __395493_395493;
   reg _395494_395494 ; 
   reg __395494_395494;
   reg _395495_395495 ; 
   reg __395495_395495;
   reg _395496_395496 ; 
   reg __395496_395496;
   reg _395497_395497 ; 
   reg __395497_395497;
   reg _395498_395498 ; 
   reg __395498_395498;
   reg _395499_395499 ; 
   reg __395499_395499;
   reg _395500_395500 ; 
   reg __395500_395500;
   reg _395501_395501 ; 
   reg __395501_395501;
   reg _395502_395502 ; 
   reg __395502_395502;
   reg _395503_395503 ; 
   reg __395503_395503;
   reg _395504_395504 ; 
   reg __395504_395504;
   reg _395505_395505 ; 
   reg __395505_395505;
   reg _395506_395506 ; 
   reg __395506_395506;
   reg _395507_395507 ; 
   reg __395507_395507;
   reg _395508_395508 ; 
   reg __395508_395508;
   reg _395509_395509 ; 
   reg __395509_395509;
   reg _395510_395510 ; 
   reg __395510_395510;
   reg _395511_395511 ; 
   reg __395511_395511;
   reg _395512_395512 ; 
   reg __395512_395512;
   reg _395513_395513 ; 
   reg __395513_395513;
   reg _395514_395514 ; 
   reg __395514_395514;
   reg _395515_395515 ; 
   reg __395515_395515;
   reg _395516_395516 ; 
   reg __395516_395516;
   reg _395517_395517 ; 
   reg __395517_395517;
   reg _395518_395518 ; 
   reg __395518_395518;
   reg _395519_395519 ; 
   reg __395519_395519;
   reg _395520_395520 ; 
   reg __395520_395520;
   reg _395521_395521 ; 
   reg __395521_395521;
   reg _395522_395522 ; 
   reg __395522_395522;
   reg _395523_395523 ; 
   reg __395523_395523;
   reg _395524_395524 ; 
   reg __395524_395524;
   reg _395525_395525 ; 
   reg __395525_395525;
   reg _395526_395526 ; 
   reg __395526_395526;
   reg _395527_395527 ; 
   reg __395527_395527;
   reg _395528_395528 ; 
   reg __395528_395528;
   reg _395529_395529 ; 
   reg __395529_395529;
   reg _395530_395530 ; 
   reg __395530_395530;
   reg _395531_395531 ; 
   reg __395531_395531;
   reg _395532_395532 ; 
   reg __395532_395532;
   reg _395533_395533 ; 
   reg __395533_395533;
   reg _395534_395534 ; 
   reg __395534_395534;
   reg _395535_395535 ; 
   reg __395535_395535;
   reg _395536_395536 ; 
   reg __395536_395536;
   reg _395537_395537 ; 
   reg __395537_395537;
   reg _395538_395538 ; 
   reg __395538_395538;
   reg _395539_395539 ; 
   reg __395539_395539;
   reg _395540_395540 ; 
   reg __395540_395540;
   reg _395541_395541 ; 
   reg __395541_395541;
   reg _395542_395542 ; 
   reg __395542_395542;
   reg _395543_395543 ; 
   reg __395543_395543;
   reg _395544_395544 ; 
   reg __395544_395544;
   reg _395545_395545 ; 
   reg __395545_395545;
   reg _395546_395546 ; 
   reg __395546_395546;
   reg _395547_395547 ; 
   reg __395547_395547;
   reg _395548_395548 ; 
   reg __395548_395548;
   reg _395549_395549 ; 
   reg __395549_395549;
   reg _395550_395550 ; 
   reg __395550_395550;
   reg _395551_395551 ; 
   reg __395551_395551;
   reg _395552_395552 ; 
   reg __395552_395552;
   reg _395553_395553 ; 
   reg __395553_395553;
   reg _395554_395554 ; 
   reg __395554_395554;
   reg _395555_395555 ; 
   reg __395555_395555;
   reg _395556_395556 ; 
   reg __395556_395556;
   reg _395557_395557 ; 
   reg __395557_395557;
   reg _395558_395558 ; 
   reg __395558_395558;
   reg _395559_395559 ; 
   reg __395559_395559;
   reg _395560_395560 ; 
   reg __395560_395560;
   reg _395561_395561 ; 
   reg __395561_395561;
   reg _395562_395562 ; 
   reg __395562_395562;
   reg _395563_395563 ; 
   reg __395563_395563;
   reg _395564_395564 ; 
   reg __395564_395564;
   reg _395565_395565 ; 
   reg __395565_395565;
   reg _395566_395566 ; 
   reg __395566_395566;
   reg _395567_395567 ; 
   reg __395567_395567;
   reg _395568_395568 ; 
   reg __395568_395568;
   reg _395569_395569 ; 
   reg __395569_395569;
   reg _395570_395570 ; 
   reg __395570_395570;
   reg _395571_395571 ; 
   reg __395571_395571;
   reg _395572_395572 ; 
   reg __395572_395572;
   reg _395573_395573 ; 
   reg __395573_395573;
   reg _395574_395574 ; 
   reg __395574_395574;
   reg _395575_395575 ; 
   reg __395575_395575;
   reg _395576_395576 ; 
   reg __395576_395576;
   reg _395577_395577 ; 
   reg __395577_395577;
   reg _395578_395578 ; 
   reg __395578_395578;
   reg _395579_395579 ; 
   reg __395579_395579;
   reg _395580_395580 ; 
   reg __395580_395580;
   reg _395581_395581 ; 
   reg __395581_395581;
   reg _395582_395582 ; 
   reg __395582_395582;
   reg _395583_395583 ; 
   reg __395583_395583;
   reg _395584_395584 ; 
   reg __395584_395584;
   reg _395585_395585 ; 
   reg __395585_395585;
   reg _395586_395586 ; 
   reg __395586_395586;
   reg _395587_395587 ; 
   reg __395587_395587;
   reg _395588_395588 ; 
   reg __395588_395588;
   reg _395589_395589 ; 
   reg __395589_395589;
   reg _395590_395590 ; 
   reg __395590_395590;
   reg _395591_395591 ; 
   reg __395591_395591;
   reg _395592_395592 ; 
   reg __395592_395592;
   reg _395593_395593 ; 
   reg __395593_395593;
   reg _395594_395594 ; 
   reg __395594_395594;
   reg _395595_395595 ; 
   reg __395595_395595;
   reg _395596_395596 ; 
   reg __395596_395596;
   reg _395597_395597 ; 
   reg __395597_395597;
   reg _395598_395598 ; 
   reg __395598_395598;
   reg _395599_395599 ; 
   reg __395599_395599;
   reg _395600_395600 ; 
   reg __395600_395600;
   reg _395601_395601 ; 
   reg __395601_395601;
   reg _395602_395602 ; 
   reg __395602_395602;
   reg _395603_395603 ; 
   reg __395603_395603;
   reg _395604_395604 ; 
   reg __395604_395604;
   reg _395605_395605 ; 
   reg __395605_395605;
   reg _395606_395606 ; 
   reg __395606_395606;
   reg _395607_395607 ; 
   reg __395607_395607;
   reg _395608_395608 ; 
   reg __395608_395608;
   reg _395609_395609 ; 
   reg __395609_395609;
   reg _395610_395610 ; 
   reg __395610_395610;
   reg _395611_395611 ; 
   reg __395611_395611;
   reg _395612_395612 ; 
   reg __395612_395612;
   reg _395613_395613 ; 
   reg __395613_395613;
   reg _395614_395614 ; 
   reg __395614_395614;
   reg _395615_395615 ; 
   reg __395615_395615;
   reg _395616_395616 ; 
   reg __395616_395616;
   reg _395617_395617 ; 
   reg __395617_395617;
   reg _395618_395618 ; 
   reg __395618_395618;
   reg _395619_395619 ; 
   reg __395619_395619;
   reg _395620_395620 ; 
   reg __395620_395620;
   reg _395621_395621 ; 
   reg __395621_395621;
   reg _395622_395622 ; 
   reg __395622_395622;
   reg _395623_395623 ; 
   reg __395623_395623;
   reg _395624_395624 ; 
   reg __395624_395624;
   reg _395625_395625 ; 
   reg __395625_395625;
   reg _395626_395626 ; 
   reg __395626_395626;
   reg _395627_395627 ; 
   reg __395627_395627;
   reg _395628_395628 ; 
   reg __395628_395628;
   reg _395629_395629 ; 
   reg __395629_395629;
   reg _395630_395630 ; 
   reg __395630_395630;
   reg _395631_395631 ; 
   reg __395631_395631;
   reg _395632_395632 ; 
   reg __395632_395632;
   reg _395633_395633 ; 
   reg __395633_395633;
   reg _395634_395634 ; 
   reg __395634_395634;
   reg _395635_395635 ; 
   reg __395635_395635;
   reg _395636_395636 ; 
   reg __395636_395636;
   reg _395637_395637 ; 
   reg __395637_395637;
   reg _395638_395638 ; 
   reg __395638_395638;
   reg _395639_395639 ; 
   reg __395639_395639;
   reg _395640_395640 ; 
   reg __395640_395640;
   reg _395641_395641 ; 
   reg __395641_395641;
   reg _395642_395642 ; 
   reg __395642_395642;
   reg _395643_395643 ; 
   reg __395643_395643;
   reg _395644_395644 ; 
   reg __395644_395644;
   reg _395645_395645 ; 
   reg __395645_395645;
   reg _395646_395646 ; 
   reg __395646_395646;
   reg _395647_395647 ; 
   reg __395647_395647;
   reg _395648_395648 ; 
   reg __395648_395648;
   reg _395649_395649 ; 
   reg __395649_395649;
   reg _395650_395650 ; 
   reg __395650_395650;
   reg _395651_395651 ; 
   reg __395651_395651;
   reg _395652_395652 ; 
   reg __395652_395652;
   reg _395653_395653 ; 
   reg __395653_395653;
   reg _395654_395654 ; 
   reg __395654_395654;
   reg _395655_395655 ; 
   reg __395655_395655;
   reg _395656_395656 ; 
   reg __395656_395656;
   reg _395657_395657 ; 
   reg __395657_395657;
   reg _395658_395658 ; 
   reg __395658_395658;
   reg _395659_395659 ; 
   reg __395659_395659;
   reg _395660_395660 ; 
   reg __395660_395660;
   reg _395661_395661 ; 
   reg __395661_395661;
   reg _395662_395662 ; 
   reg __395662_395662;
   reg _395663_395663 ; 
   reg __395663_395663;
   reg _395664_395664 ; 
   reg __395664_395664;
   reg _395665_395665 ; 
   reg __395665_395665;
   reg _395666_395666 ; 
   reg __395666_395666;
   reg _395667_395667 ; 
   reg __395667_395667;
   reg _395668_395668 ; 
   reg __395668_395668;
   reg _395669_395669 ; 
   reg __395669_395669;
   reg _395670_395670 ; 
   reg __395670_395670;
   reg _395671_395671 ; 
   reg __395671_395671;
   reg _395672_395672 ; 
   reg __395672_395672;
   reg _395673_395673 ; 
   reg __395673_395673;
   reg _395674_395674 ; 
   reg __395674_395674;
   reg _395675_395675 ; 
   reg __395675_395675;
   reg _395676_395676 ; 
   reg __395676_395676;
   reg _395677_395677 ; 
   reg __395677_395677;
   reg _395678_395678 ; 
   reg __395678_395678;
   reg _395679_395679 ; 
   reg __395679_395679;
   reg _395680_395680 ; 
   reg __395680_395680;
   reg _395681_395681 ; 
   reg __395681_395681;
   reg _395682_395682 ; 
   reg __395682_395682;
   reg _395683_395683 ; 
   reg __395683_395683;
   reg _395684_395684 ; 
   reg __395684_395684;
   reg _395685_395685 ; 
   reg __395685_395685;
   reg _395686_395686 ; 
   reg __395686_395686;
   reg _395687_395687 ; 
   reg __395687_395687;
   reg _395688_395688 ; 
   reg __395688_395688;
   reg _395689_395689 ; 
   reg __395689_395689;
   reg _395690_395690 ; 
   reg __395690_395690;
   reg _395691_395691 ; 
   reg __395691_395691;
   reg _395692_395692 ; 
   reg __395692_395692;
   reg _395693_395693 ; 
   reg __395693_395693;
   reg _395694_395694 ; 
   reg __395694_395694;
   reg _395695_395695 ; 
   reg __395695_395695;
   reg _395696_395696 ; 
   reg __395696_395696;
   reg _395697_395697 ; 
   reg __395697_395697;
   reg _395698_395698 ; 
   reg __395698_395698;
   reg _395699_395699 ; 
   reg __395699_395699;
   reg _395700_395700 ; 
   reg __395700_395700;
   reg _395701_395701 ; 
   reg __395701_395701;
   reg _395702_395702 ; 
   reg __395702_395702;
   reg _395703_395703 ; 
   reg __395703_395703;
   reg _395704_395704 ; 
   reg __395704_395704;
   reg _395705_395705 ; 
   reg __395705_395705;
   reg _395706_395706 ; 
   reg __395706_395706;
   reg _395707_395707 ; 
   reg __395707_395707;
   reg _395708_395708 ; 
   reg __395708_395708;
   reg _395709_395709 ; 
   reg __395709_395709;
   reg _395710_395710 ; 
   reg __395710_395710;
   reg _395711_395711 ; 
   reg __395711_395711;
   reg _395712_395712 ; 
   reg __395712_395712;
   reg _395713_395713 ; 
   reg __395713_395713;
   reg _395714_395714 ; 
   reg __395714_395714;
   reg _395715_395715 ; 
   reg __395715_395715;
   reg _395716_395716 ; 
   reg __395716_395716;
   reg _395717_395717 ; 
   reg __395717_395717;
   reg _395718_395718 ; 
   reg __395718_395718;
   reg _395719_395719 ; 
   reg __395719_395719;
   reg _395720_395720 ; 
   reg __395720_395720;
   reg _395721_395721 ; 
   reg __395721_395721;
   reg _395722_395722 ; 
   reg __395722_395722;
   reg _395723_395723 ; 
   reg __395723_395723;
   reg _395724_395724 ; 
   reg __395724_395724;
   reg _395725_395725 ; 
   reg __395725_395725;
   reg _395726_395726 ; 
   reg __395726_395726;
   reg _395727_395727 ; 
   reg __395727_395727;
   reg _395728_395728 ; 
   reg __395728_395728;
   reg _395729_395729 ; 
   reg __395729_395729;
   reg _395730_395730 ; 
   reg __395730_395730;
   reg _395731_395731 ; 
   reg __395731_395731;
   reg _395732_395732 ; 
   reg __395732_395732;
   reg _395733_395733 ; 
   reg __395733_395733;
   reg _395734_395734 ; 
   reg __395734_395734;
   reg _395735_395735 ; 
   reg __395735_395735;
   reg _395736_395736 ; 
   reg __395736_395736;
   reg _395737_395737 ; 
   reg __395737_395737;
   reg _395738_395738 ; 
   reg __395738_395738;
   reg _395739_395739 ; 
   reg __395739_395739;
   reg _395740_395740 ; 
   reg __395740_395740;
   reg _395741_395741 ; 
   reg __395741_395741;
   reg _395742_395742 ; 
   reg __395742_395742;
   reg _395743_395743 ; 
   reg __395743_395743;
   reg _395744_395744 ; 
   reg __395744_395744;
   reg _395745_395745 ; 
   reg __395745_395745;
   reg _395746_395746 ; 
   reg __395746_395746;
   reg _395747_395747 ; 
   reg __395747_395747;
   reg _395748_395748 ; 
   reg __395748_395748;
   reg _395749_395749 ; 
   reg __395749_395749;
   reg _395750_395750 ; 
   reg __395750_395750;
   reg _395751_395751 ; 
   reg __395751_395751;
   reg _395752_395752 ; 
   reg __395752_395752;
   reg _395753_395753 ; 
   reg __395753_395753;
   reg _395754_395754 ; 
   reg __395754_395754;
   reg _395755_395755 ; 
   reg __395755_395755;
   reg _395756_395756 ; 
   reg __395756_395756;
   reg _395757_395757 ; 
   reg __395757_395757;
   reg _395758_395758 ; 
   reg __395758_395758;
   reg _395759_395759 ; 
   reg __395759_395759;
   reg _395760_395760 ; 
   reg __395760_395760;
   reg _395761_395761 ; 
   reg __395761_395761;
   reg _395762_395762 ; 
   reg __395762_395762;
   reg _395763_395763 ; 
   reg __395763_395763;
   reg _395764_395764 ; 
   reg __395764_395764;
   reg _395765_395765 ; 
   reg __395765_395765;
   reg _395766_395766 ; 
   reg __395766_395766;
   reg _395767_395767 ; 
   reg __395767_395767;
   reg _395768_395768 ; 
   reg __395768_395768;
   reg _395769_395769 ; 
   reg __395769_395769;
   reg _395770_395770 ; 
   reg __395770_395770;
   reg _395771_395771 ; 
   reg __395771_395771;
   reg _395772_395772 ; 
   reg __395772_395772;
   reg _395773_395773 ; 
   reg __395773_395773;
   reg _395774_395774 ; 
   reg __395774_395774;
   reg _395775_395775 ; 
   reg __395775_395775;
   reg _395776_395776 ; 
   reg __395776_395776;
   reg _395777_395777 ; 
   reg __395777_395777;
   reg _395778_395778 ; 
   reg __395778_395778;
   reg _395779_395779 ; 
   reg __395779_395779;
   reg _395780_395780 ; 
   reg __395780_395780;
   reg _395781_395781 ; 
   reg __395781_395781;
   reg _395782_395782 ; 
   reg __395782_395782;
   reg _395783_395783 ; 
   reg __395783_395783;
   reg _395784_395784 ; 
   reg __395784_395784;
   reg _395785_395785 ; 
   reg __395785_395785;
   reg _395786_395786 ; 
   reg __395786_395786;
   reg _395787_395787 ; 
   reg __395787_395787;
   reg _395788_395788 ; 
   reg __395788_395788;
   reg _395789_395789 ; 
   reg __395789_395789;
   reg _395790_395790 ; 
   reg __395790_395790;
   reg _395791_395791 ; 
   reg __395791_395791;
   reg _395792_395792 ; 
   reg __395792_395792;
   reg _395793_395793 ; 
   reg __395793_395793;
   reg _395794_395794 ; 
   reg __395794_395794;
   reg _395795_395795 ; 
   reg __395795_395795;
   reg _395796_395796 ; 
   reg __395796_395796;
   reg _395797_395797 ; 
   reg __395797_395797;
   reg _395798_395798 ; 
   reg __395798_395798;
   reg _395799_395799 ; 
   reg __395799_395799;
   reg _395800_395800 ; 
   reg __395800_395800;
   reg _395801_395801 ; 
   reg __395801_395801;
   reg _395802_395802 ; 
   reg __395802_395802;
   reg _395803_395803 ; 
   reg __395803_395803;
   reg _395804_395804 ; 
   reg __395804_395804;
   reg _395805_395805 ; 
   reg __395805_395805;
   reg _395806_395806 ; 
   reg __395806_395806;
   reg _395807_395807 ; 
   reg __395807_395807;
   reg _395808_395808 ; 
   reg __395808_395808;
   reg _395809_395809 ; 
   reg __395809_395809;
   reg _395810_395810 ; 
   reg __395810_395810;
   reg _395811_395811 ; 
   reg __395811_395811;
   reg _395812_395812 ; 
   reg __395812_395812;
   reg _395813_395813 ; 
   reg __395813_395813;
   reg _395814_395814 ; 
   reg __395814_395814;
   reg _395815_395815 ; 
   reg __395815_395815;
   reg _395816_395816 ; 
   reg __395816_395816;
   reg _395817_395817 ; 
   reg __395817_395817;
   reg _395818_395818 ; 
   reg __395818_395818;
   reg _395819_395819 ; 
   reg __395819_395819;
   reg _395820_395820 ; 
   reg __395820_395820;
   reg _395821_395821 ; 
   reg __395821_395821;
   reg _395822_395822 ; 
   reg __395822_395822;
   reg _395823_395823 ; 
   reg __395823_395823;
   reg _395824_395824 ; 
   reg __395824_395824;
   reg _395825_395825 ; 
   reg __395825_395825;
   reg _395826_395826 ; 
   reg __395826_395826;
   reg _395827_395827 ; 
   reg __395827_395827;
   reg _395828_395828 ; 
   reg __395828_395828;
   reg _395829_395829 ; 
   reg __395829_395829;
   reg _395830_395830 ; 
   reg __395830_395830;
   reg _395831_395831 ; 
   reg __395831_395831;
   reg _395832_395832 ; 
   reg __395832_395832;
   reg _395833_395833 ; 
   reg __395833_395833;
   reg _395834_395834 ; 
   reg __395834_395834;
   reg _395835_395835 ; 
   reg __395835_395835;
   reg _395836_395836 ; 
   reg __395836_395836;
   reg _395837_395837 ; 
   reg __395837_395837;
   reg _395838_395838 ; 
   reg __395838_395838;
   reg _395839_395839 ; 
   reg __395839_395839;
   reg _395840_395840 ; 
   reg __395840_395840;
   reg _395841_395841 ; 
   reg __395841_395841;
   reg _395842_395842 ; 
   reg __395842_395842;
   reg _395843_395843 ; 
   reg __395843_395843;
   reg _395844_395844 ; 
   reg __395844_395844;
   reg _395845_395845 ; 
   reg __395845_395845;
   reg _395846_395846 ; 
   reg __395846_395846;
   reg _395847_395847 ; 
   reg __395847_395847;
   reg _395848_395848 ; 
   reg __395848_395848;
   reg _395849_395849 ; 
   reg __395849_395849;
   reg _395850_395850 ; 
   reg __395850_395850;
   reg _395851_395851 ; 
   reg __395851_395851;
   reg _395852_395852 ; 
   reg __395852_395852;
   reg _395853_395853 ; 
   reg __395853_395853;
   reg _395854_395854 ; 
   reg __395854_395854;
   reg _395855_395855 ; 
   reg __395855_395855;
   reg _395856_395856 ; 
   reg __395856_395856;
   reg _395857_395857 ; 
   reg __395857_395857;
   reg _395858_395858 ; 
   reg __395858_395858;
   reg _395859_395859 ; 
   reg __395859_395859;
   reg _395860_395860 ; 
   reg __395860_395860;
   reg _395861_395861 ; 
   reg __395861_395861;
   reg _395862_395862 ; 
   reg __395862_395862;
   reg _395863_395863 ; 
   reg __395863_395863;
   reg _395864_395864 ; 
   reg __395864_395864;
   reg _395865_395865 ; 
   reg __395865_395865;
   reg _395866_395866 ; 
   reg __395866_395866;
   reg _395867_395867 ; 
   reg __395867_395867;
   reg _395868_395868 ; 
   reg __395868_395868;
   reg _395869_395869 ; 
   reg __395869_395869;
   reg _395870_395870 ; 
   reg __395870_395870;
   reg _395871_395871 ; 
   reg __395871_395871;
   reg _395872_395872 ; 
   reg __395872_395872;
   reg _395873_395873 ; 
   reg __395873_395873;
   reg _395874_395874 ; 
   reg __395874_395874;
   reg _395875_395875 ; 
   reg __395875_395875;
   reg _395876_395876 ; 
   reg __395876_395876;
   reg _395877_395877 ; 
   reg __395877_395877;
   reg _395878_395878 ; 
   reg __395878_395878;
   reg _395879_395879 ; 
   reg __395879_395879;
   reg _395880_395880 ; 
   reg __395880_395880;
   reg _395881_395881 ; 
   reg __395881_395881;
   reg _395882_395882 ; 
   reg __395882_395882;
   reg _395883_395883 ; 
   reg __395883_395883;
   reg _395884_395884 ; 
   reg __395884_395884;
   reg _395885_395885 ; 
   reg __395885_395885;
   reg _395886_395886 ; 
   reg __395886_395886;
   reg _395887_395887 ; 
   reg __395887_395887;
   reg _395888_395888 ; 
   reg __395888_395888;
   reg _395889_395889 ; 
   reg __395889_395889;
   reg _395890_395890 ; 
   reg __395890_395890;
   reg _395891_395891 ; 
   reg __395891_395891;
   reg _395892_395892 ; 
   reg __395892_395892;
   reg _395893_395893 ; 
   reg __395893_395893;
   reg _395894_395894 ; 
   reg __395894_395894;
   reg _395895_395895 ; 
   reg __395895_395895;
   reg _395896_395896 ; 
   reg __395896_395896;
   reg _395897_395897 ; 
   reg __395897_395897;
   reg _395898_395898 ; 
   reg __395898_395898;
   reg _395899_395899 ; 
   reg __395899_395899;
   reg _395900_395900 ; 
   reg __395900_395900;
   reg _395901_395901 ; 
   reg __395901_395901;
   reg _395902_395902 ; 
   reg __395902_395902;
   reg _395903_395903 ; 
   reg __395903_395903;
   reg _395904_395904 ; 
   reg __395904_395904;
   reg _395905_395905 ; 
   reg __395905_395905;
   reg _395906_395906 ; 
   reg __395906_395906;
   reg _395907_395907 ; 
   reg __395907_395907;
   reg _395908_395908 ; 
   reg __395908_395908;
   reg _395909_395909 ; 
   reg __395909_395909;
   reg _395910_395910 ; 
   reg __395910_395910;
   reg _395911_395911 ; 
   reg __395911_395911;
   reg _395912_395912 ; 
   reg __395912_395912;
   reg _395913_395913 ; 
   reg __395913_395913;
   reg _395914_395914 ; 
   reg __395914_395914;
   reg _395915_395915 ; 
   reg __395915_395915;
   reg _395916_395916 ; 
   reg __395916_395916;
   reg _395917_395917 ; 
   reg __395917_395917;
   reg _395918_395918 ; 
   reg __395918_395918;
   reg _395919_395919 ; 
   reg __395919_395919;
   reg _395920_395920 ; 
   reg __395920_395920;
   reg _395921_395921 ; 
   reg __395921_395921;
   reg _395922_395922 ; 
   reg __395922_395922;
   reg _395923_395923 ; 
   reg __395923_395923;
   reg _395924_395924 ; 
   reg __395924_395924;
   reg _395925_395925 ; 
   reg __395925_395925;
   reg _395926_395926 ; 
   reg __395926_395926;
   reg _395927_395927 ; 
   reg __395927_395927;
   reg _395928_395928 ; 
   reg __395928_395928;
   reg _395929_395929 ; 
   reg __395929_395929;
   reg _395930_395930 ; 
   reg __395930_395930;
   reg _395931_395931 ; 
   reg __395931_395931;
   reg _395932_395932 ; 
   reg __395932_395932;
   reg _395933_395933 ; 
   reg __395933_395933;
   reg _395934_395934 ; 
   reg __395934_395934;
   reg _395935_395935 ; 
   reg __395935_395935;
   reg _395936_395936 ; 
   reg __395936_395936;
   reg _395937_395937 ; 
   reg __395937_395937;
   reg _395938_395938 ; 
   reg __395938_395938;
   reg _395939_395939 ; 
   reg __395939_395939;
   reg _395940_395940 ; 
   reg __395940_395940;
   reg _395941_395941 ; 
   reg __395941_395941;
   reg _395942_395942 ; 
   reg __395942_395942;
   reg _395943_395943 ; 
   reg __395943_395943;
   reg _395944_395944 ; 
   reg __395944_395944;
   reg _395945_395945 ; 
   reg __395945_395945;
   reg _395946_395946 ; 
   reg __395946_395946;
   reg _395947_395947 ; 
   reg __395947_395947;
   reg _395948_395948 ; 
   reg __395948_395948;
   reg _395949_395949 ; 
   reg __395949_395949;
   reg _395950_395950 ; 
   reg __395950_395950;
   reg _395951_395951 ; 
   reg __395951_395951;
   reg _395952_395952 ; 
   reg __395952_395952;
   reg _395953_395953 ; 
   reg __395953_395953;
   reg _395954_395954 ; 
   reg __395954_395954;
   reg _395955_395955 ; 
   reg __395955_395955;
   reg _395956_395956 ; 
   reg __395956_395956;
   reg _395957_395957 ; 
   reg __395957_395957;
   reg _395958_395958 ; 
   reg __395958_395958;
   reg _395959_395959 ; 
   reg __395959_395959;
   reg _395960_395960 ; 
   reg __395960_395960;
   reg _395961_395961 ; 
   reg __395961_395961;
   reg _395962_395962 ; 
   reg __395962_395962;
   reg _395963_395963 ; 
   reg __395963_395963;
   reg _395964_395964 ; 
   reg __395964_395964;
   reg _395965_395965 ; 
   reg __395965_395965;
   reg _395966_395966 ; 
   reg __395966_395966;
   reg _395967_395967 ; 
   reg __395967_395967;
   reg _395968_395968 ; 
   reg __395968_395968;
   reg _395969_395969 ; 
   reg __395969_395969;
   reg _395970_395970 ; 
   reg __395970_395970;
   reg _395971_395971 ; 
   reg __395971_395971;
   reg _395972_395972 ; 
   reg __395972_395972;
   reg _395973_395973 ; 
   reg __395973_395973;
   reg _395974_395974 ; 
   reg __395974_395974;
   reg _395975_395975 ; 
   reg __395975_395975;
   reg _395976_395976 ; 
   reg __395976_395976;
   reg _395977_395977 ; 
   reg __395977_395977;
   reg _395978_395978 ; 
   reg __395978_395978;
   reg _395979_395979 ; 
   reg __395979_395979;
   reg _395980_395980 ; 
   reg __395980_395980;
   reg _395981_395981 ; 
   reg __395981_395981;
   reg _395982_395982 ; 
   reg __395982_395982;
   reg _395983_395983 ; 
   reg __395983_395983;
   reg _395984_395984 ; 
   reg __395984_395984;
   reg _395985_395985 ; 
   reg __395985_395985;
   reg _395986_395986 ; 
   reg __395986_395986;
   reg _395987_395987 ; 
   reg __395987_395987;
   reg _395988_395988 ; 
   reg __395988_395988;
   reg _395989_395989 ; 
   reg __395989_395989;
   reg _395990_395990 ; 
   reg __395990_395990;
   reg _395991_395991 ; 
   reg __395991_395991;
   reg _395992_395992 ; 
   reg __395992_395992;
   reg _395993_395993 ; 
   reg __395993_395993;
   reg _395994_395994 ; 
   reg __395994_395994;
   reg _395995_395995 ; 
   reg __395995_395995;
   reg _395996_395996 ; 
   reg __395996_395996;
   reg _395997_395997 ; 
   reg __395997_395997;
   reg _395998_395998 ; 
   reg __395998_395998;
   reg _395999_395999 ; 
   reg __395999_395999;
   reg _396000_396000 ; 
   reg __396000_396000;
   reg _396001_396001 ; 
   reg __396001_396001;
   reg _396002_396002 ; 
   reg __396002_396002;
   reg _396003_396003 ; 
   reg __396003_396003;
   reg _396004_396004 ; 
   reg __396004_396004;
   reg _396005_396005 ; 
   reg __396005_396005;
   reg _396006_396006 ; 
   reg __396006_396006;
   reg _396007_396007 ; 
   reg __396007_396007;
   reg _396008_396008 ; 
   reg __396008_396008;
   reg _396009_396009 ; 
   reg __396009_396009;
   reg _396010_396010 ; 
   reg __396010_396010;
   reg _396011_396011 ; 
   reg __396011_396011;
   reg _396012_396012 ; 
   reg __396012_396012;
   reg _396013_396013 ; 
   reg __396013_396013;
   reg _396014_396014 ; 
   reg __396014_396014;
   reg _396015_396015 ; 
   reg __396015_396015;
   reg _396016_396016 ; 
   reg __396016_396016;
   reg _396017_396017 ; 
   reg __396017_396017;
   reg _396018_396018 ; 
   reg __396018_396018;
   reg _396019_396019 ; 
   reg __396019_396019;
   reg _396020_396020 ; 
   reg __396020_396020;
   reg _396021_396021 ; 
   reg __396021_396021;
   reg _396022_396022 ; 
   reg __396022_396022;
   reg _396023_396023 ; 
   reg __396023_396023;
   reg _396024_396024 ; 
   reg __396024_396024;
   reg _396025_396025 ; 
   reg __396025_396025;
   reg _396026_396026 ; 
   reg __396026_396026;
   reg _396027_396027 ; 
   reg __396027_396027;
   reg _396028_396028 ; 
   reg __396028_396028;
   reg _396029_396029 ; 
   reg __396029_396029;
   reg _396030_396030 ; 
   reg __396030_396030;
   reg _396031_396031 ; 
   reg __396031_396031;
   reg _396032_396032 ; 
   reg __396032_396032;
   reg _396033_396033 ; 
   reg __396033_396033;
   reg _396034_396034 ; 
   reg __396034_396034;
   reg _396035_396035 ; 
   reg __396035_396035;
   reg _396036_396036 ; 
   reg __396036_396036;
   reg _396037_396037 ; 
   reg __396037_396037;
   reg _396038_396038 ; 
   reg __396038_396038;
   reg _396039_396039 ; 
   reg __396039_396039;
   reg _396040_396040 ; 
   reg __396040_396040;
   reg _396041_396041 ; 
   reg __396041_396041;
   reg _396042_396042 ; 
   reg __396042_396042;
   reg _396043_396043 ; 
   reg __396043_396043;
   reg _396044_396044 ; 
   reg __396044_396044;
   reg _396045_396045 ; 
   reg __396045_396045;
   reg _396046_396046 ; 
   reg __396046_396046;
   reg _396047_396047 ; 
   reg __396047_396047;
   reg _396048_396048 ; 
   reg __396048_396048;
   reg _396049_396049 ; 
   reg __396049_396049;
   reg _396050_396050 ; 
   reg __396050_396050;
   reg _396051_396051 ; 
   reg __396051_396051;
   reg _396052_396052 ; 
   reg __396052_396052;
   reg _396053_396053 ; 
   reg __396053_396053;
   reg _396054_396054 ; 
   reg __396054_396054;
   reg _396055_396055 ; 
   reg __396055_396055;
   reg _396056_396056 ; 
   reg __396056_396056;
   reg _396057_396057 ; 
   reg __396057_396057;
   reg _396058_396058 ; 
   reg __396058_396058;
   reg _396059_396059 ; 
   reg __396059_396059;
   reg _396060_396060 ; 
   reg __396060_396060;
   reg _396061_396061 ; 
   reg __396061_396061;
   reg _396062_396062 ; 
   reg __396062_396062;
   reg _396063_396063 ; 
   reg __396063_396063;
   reg _396064_396064 ; 
   reg __396064_396064;
   reg _396065_396065 ; 
   reg __396065_396065;
   reg _396066_396066 ; 
   reg __396066_396066;
   reg _396067_396067 ; 
   reg __396067_396067;
   reg _396068_396068 ; 
   reg __396068_396068;
   reg _396069_396069 ; 
   reg __396069_396069;
   reg _396070_396070 ; 
   reg __396070_396070;
   reg _396071_396071 ; 
   reg __396071_396071;
   reg _396072_396072 ; 
   reg __396072_396072;
   reg _396073_396073 ; 
   reg __396073_396073;
   reg _396074_396074 ; 
   reg __396074_396074;
   reg _396075_396075 ; 
   reg __396075_396075;
   reg _396076_396076 ; 
   reg __396076_396076;
   reg _396077_396077 ; 
   reg __396077_396077;
   reg _396078_396078 ; 
   reg __396078_396078;
   reg _396079_396079 ; 
   reg __396079_396079;
   reg _396080_396080 ; 
   reg __396080_396080;
   reg _396081_396081 ; 
   reg __396081_396081;
   reg _396082_396082 ; 
   reg __396082_396082;
   reg _396083_396083 ; 
   reg __396083_396083;
   reg _396084_396084 ; 
   reg __396084_396084;
   reg _396085_396085 ; 
   reg __396085_396085;
   reg _396086_396086 ; 
   reg __396086_396086;
   reg _396087_396087 ; 
   reg __396087_396087;
   reg _396088_396088 ; 
   reg __396088_396088;
   reg _396089_396089 ; 
   reg __396089_396089;
   reg _396090_396090 ; 
   reg __396090_396090;
   reg _396091_396091 ; 
   reg __396091_396091;
   reg _396092_396092 ; 
   reg __396092_396092;
   reg _396093_396093 ; 
   reg __396093_396093;
   reg _396094_396094 ; 
   reg __396094_396094;
   reg _396095_396095 ; 
   reg __396095_396095;
   reg _396096_396096 ; 
   reg __396096_396096;
   reg _396097_396097 ; 
   reg __396097_396097;
   reg _396098_396098 ; 
   reg __396098_396098;
   reg _396099_396099 ; 
   reg __396099_396099;
   reg _396100_396100 ; 
   reg __396100_396100;
   reg _396101_396101 ; 
   reg __396101_396101;
   reg _396102_396102 ; 
   reg __396102_396102;
   reg _396103_396103 ; 
   reg __396103_396103;
   reg _396104_396104 ; 
   reg __396104_396104;
   reg _396105_396105 ; 
   reg __396105_396105;
   reg _396106_396106 ; 
   reg __396106_396106;
   reg _396107_396107 ; 
   reg __396107_396107;
   reg _396108_396108 ; 
   reg __396108_396108;
   reg _396109_396109 ; 
   reg __396109_396109;
   reg _396110_396110 ; 
   reg __396110_396110;
   reg _396111_396111 ; 
   reg __396111_396111;
   reg _396112_396112 ; 
   reg __396112_396112;
   reg _396113_396113 ; 
   reg __396113_396113;
   reg _396114_396114 ; 
   reg __396114_396114;
   reg _396115_396115 ; 
   reg __396115_396115;
   reg _396116_396116 ; 
   reg __396116_396116;
   reg _396117_396117 ; 
   reg __396117_396117;
   reg _396118_396118 ; 
   reg __396118_396118;
   reg _396119_396119 ; 
   reg __396119_396119;
   reg _396120_396120 ; 
   reg __396120_396120;
   reg _396121_396121 ; 
   reg __396121_396121;
   reg _396122_396122 ; 
   reg __396122_396122;
   reg _396123_396123 ; 
   reg __396123_396123;
   reg _396124_396124 ; 
   reg __396124_396124;
   reg _396125_396125 ; 
   reg __396125_396125;
   reg _396126_396126 ; 
   reg __396126_396126;
   reg _396127_396127 ; 
   reg __396127_396127;
   reg _396128_396128 ; 
   reg __396128_396128;
   reg _396129_396129 ; 
   reg __396129_396129;
   reg _396130_396130 ; 
   reg __396130_396130;
   reg _396131_396131 ; 
   reg __396131_396131;
   reg _396132_396132 ; 
   reg __396132_396132;
   reg _396133_396133 ; 
   reg __396133_396133;
   reg _396134_396134 ; 
   reg __396134_396134;
   reg _396135_396135 ; 
   reg __396135_396135;
   reg _396136_396136 ; 
   reg __396136_396136;
   reg _396137_396137 ; 
   reg __396137_396137;
   reg _396138_396138 ; 
   reg __396138_396138;
   reg _396139_396139 ; 
   reg __396139_396139;
   reg _396140_396140 ; 
   reg __396140_396140;
   reg _396141_396141 ; 
   reg __396141_396141;
   reg _396142_396142 ; 
   reg __396142_396142;
   reg _396143_396143 ; 
   reg __396143_396143;
   reg _396144_396144 ; 
   reg __396144_396144;
   reg _396145_396145 ; 
   reg __396145_396145;
   reg _396146_396146 ; 
   reg __396146_396146;
   reg _396147_396147 ; 
   reg __396147_396147;
   reg _396148_396148 ; 
   reg __396148_396148;
   reg _396149_396149 ; 
   reg __396149_396149;
   reg _396150_396150 ; 
   reg __396150_396150;
   reg _396151_396151 ; 
   reg __396151_396151;
   reg _396152_396152 ; 
   reg __396152_396152;
   reg _396153_396153 ; 
   reg __396153_396153;
   reg _396154_396154 ; 
   reg __396154_396154;
   reg _396155_396155 ; 
   reg __396155_396155;
   reg _396156_396156 ; 
   reg __396156_396156;
   reg _396157_396157 ; 
   reg __396157_396157;
   reg _396158_396158 ; 
   reg __396158_396158;
   reg _396159_396159 ; 
   reg __396159_396159;
   reg _396160_396160 ; 
   reg __396160_396160;
   reg _396161_396161 ; 
   reg __396161_396161;
   reg _396162_396162 ; 
   reg __396162_396162;
   reg _396163_396163 ; 
   reg __396163_396163;
   reg _396164_396164 ; 
   reg __396164_396164;
   reg _396165_396165 ; 
   reg __396165_396165;
   reg _396166_396166 ; 
   reg __396166_396166;
   reg _396167_396167 ; 
   reg __396167_396167;
   reg _396168_396168 ; 
   reg __396168_396168;
   reg _396169_396169 ; 
   reg __396169_396169;
   reg _396170_396170 ; 
   reg __396170_396170;
   reg _396171_396171 ; 
   reg __396171_396171;
   reg _396172_396172 ; 
   reg __396172_396172;
   reg _396173_396173 ; 
   reg __396173_396173;
   reg _396174_396174 ; 
   reg __396174_396174;
   reg _396175_396175 ; 
   reg __396175_396175;
   reg _396176_396176 ; 
   reg __396176_396176;
   reg _396177_396177 ; 
   reg __396177_396177;
   reg _396178_396178 ; 
   reg __396178_396178;
   reg _396179_396179 ; 
   reg __396179_396179;
   reg _396180_396180 ; 
   reg __396180_396180;
   reg _396181_396181 ; 
   reg __396181_396181;
   reg _396182_396182 ; 
   reg __396182_396182;
   reg _396183_396183 ; 
   reg __396183_396183;
   reg _396184_396184 ; 
   reg __396184_396184;
   reg _396185_396185 ; 
   reg __396185_396185;
   reg _396186_396186 ; 
   reg __396186_396186;
   reg _396187_396187 ; 
   reg __396187_396187;
   reg _396188_396188 ; 
   reg __396188_396188;
   reg _396189_396189 ; 
   reg __396189_396189;
   reg _396190_396190 ; 
   reg __396190_396190;
   reg _396191_396191 ; 
   reg __396191_396191;
   reg _396192_396192 ; 
   reg __396192_396192;
   reg _396193_396193 ; 
   reg __396193_396193;
   reg _396194_396194 ; 
   reg __396194_396194;
   reg _396195_396195 ; 
   reg __396195_396195;
   reg _396196_396196 ; 
   reg __396196_396196;
   reg _396197_396197 ; 
   reg __396197_396197;
   reg _396198_396198 ; 
   reg __396198_396198;
   reg _396199_396199 ; 
   reg __396199_396199;
   reg _396200_396200 ; 
   reg __396200_396200;
   reg _396201_396201 ; 
   reg __396201_396201;
   reg _396202_396202 ; 
   reg __396202_396202;
   reg _396203_396203 ; 
   reg __396203_396203;
   reg _396204_396204 ; 
   reg __396204_396204;
   reg _396205_396205 ; 
   reg __396205_396205;
   reg _396206_396206 ; 
   reg __396206_396206;
   reg _396207_396207 ; 
   reg __396207_396207;
   reg _396208_396208 ; 
   reg __396208_396208;
   reg _396209_396209 ; 
   reg __396209_396209;
   reg _396210_396210 ; 
   reg __396210_396210;
   reg _396211_396211 ; 
   reg __396211_396211;
   reg _396212_396212 ; 
   reg __396212_396212;
   reg _396213_396213 ; 
   reg __396213_396213;
   reg _396214_396214 ; 
   reg __396214_396214;
   reg _396215_396215 ; 
   reg __396215_396215;
   reg _396216_396216 ; 
   reg __396216_396216;
   reg _396217_396217 ; 
   reg __396217_396217;
   reg _396218_396218 ; 
   reg __396218_396218;
   reg _396219_396219 ; 
   reg __396219_396219;
   reg _396220_396220 ; 
   reg __396220_396220;
   reg _396221_396221 ; 
   reg __396221_396221;
   reg _396222_396222 ; 
   reg __396222_396222;
   reg _396223_396223 ; 
   reg __396223_396223;
   reg _396224_396224 ; 
   reg __396224_396224;
   reg _396225_396225 ; 
   reg __396225_396225;
   reg _396226_396226 ; 
   reg __396226_396226;
   reg _396227_396227 ; 
   reg __396227_396227;
   reg _396228_396228 ; 
   reg __396228_396228;
   reg _396229_396229 ; 
   reg __396229_396229;
   reg _396230_396230 ; 
   reg __396230_396230;
   reg _396231_396231 ; 
   reg __396231_396231;
   reg _396232_396232 ; 
   reg __396232_396232;
   reg _396233_396233 ; 
   reg __396233_396233;
   reg _396234_396234 ; 
   reg __396234_396234;
   reg _396235_396235 ; 
   reg __396235_396235;
   reg _396236_396236 ; 
   reg __396236_396236;
   reg _396237_396237 ; 
   reg __396237_396237;
   reg _396238_396238 ; 
   reg __396238_396238;
   reg _396239_396239 ; 
   reg __396239_396239;
   reg _396240_396240 ; 
   reg __396240_396240;
   reg _396241_396241 ; 
   reg __396241_396241;
   reg _396242_396242 ; 
   reg __396242_396242;
   reg _396243_396243 ; 
   reg __396243_396243;
   reg _396244_396244 ; 
   reg __396244_396244;
   reg _396245_396245 ; 
   reg __396245_396245;
   reg _396246_396246 ; 
   reg __396246_396246;
   reg _396247_396247 ; 
   reg __396247_396247;
   reg _396248_396248 ; 
   reg __396248_396248;
   reg _396249_396249 ; 
   reg __396249_396249;
   reg _396250_396250 ; 
   reg __396250_396250;
   reg _396251_396251 ; 
   reg __396251_396251;
   reg _396252_396252 ; 
   reg __396252_396252;
   reg _396253_396253 ; 
   reg __396253_396253;
   reg _396254_396254 ; 
   reg __396254_396254;
   reg _396255_396255 ; 
   reg __396255_396255;
   reg _396256_396256 ; 
   reg __396256_396256;
   reg _396257_396257 ; 
   reg __396257_396257;
   reg _396258_396258 ; 
   reg __396258_396258;
   reg _396259_396259 ; 
   reg __396259_396259;
   reg _396260_396260 ; 
   reg __396260_396260;
   reg _396261_396261 ; 
   reg __396261_396261;
   reg _396262_396262 ; 
   reg __396262_396262;
   reg _396263_396263 ; 
   reg __396263_396263;
   reg _396264_396264 ; 
   reg __396264_396264;
   reg _396265_396265 ; 
   reg __396265_396265;
   reg _396266_396266 ; 
   reg __396266_396266;
   reg _396267_396267 ; 
   reg __396267_396267;
   reg _396268_396268 ; 
   reg __396268_396268;
   reg _396269_396269 ; 
   reg __396269_396269;
   reg _396270_396270 ; 
   reg __396270_396270;
   reg _396271_396271 ; 
   reg __396271_396271;
   reg _396272_396272 ; 
   reg __396272_396272;
   reg _396273_396273 ; 
   reg __396273_396273;
   reg _396274_396274 ; 
   reg __396274_396274;
   reg _396275_396275 ; 
   reg __396275_396275;
   reg _396276_396276 ; 
   reg __396276_396276;
   reg _396277_396277 ; 
   reg __396277_396277;
   reg _396278_396278 ; 
   reg __396278_396278;
   reg _396279_396279 ; 
   reg __396279_396279;
   reg _396280_396280 ; 
   reg __396280_396280;
   reg _396281_396281 ; 
   reg __396281_396281;
   reg _396282_396282 ; 
   reg __396282_396282;
   reg _396283_396283 ; 
   reg __396283_396283;
   reg _396284_396284 ; 
   reg __396284_396284;
   reg _396285_396285 ; 
   reg __396285_396285;
   reg _396286_396286 ; 
   reg __396286_396286;
   reg _396287_396287 ; 
   reg __396287_396287;
   reg _396288_396288 ; 
   reg __396288_396288;
   reg _396289_396289 ; 
   reg __396289_396289;
   reg _396290_396290 ; 
   reg __396290_396290;
   reg _396291_396291 ; 
   reg __396291_396291;
   reg _396292_396292 ; 
   reg __396292_396292;
   reg _396293_396293 ; 
   reg __396293_396293;
   reg _396294_396294 ; 
   reg __396294_396294;
   reg _396295_396295 ; 
   reg __396295_396295;
   reg _396296_396296 ; 
   reg __396296_396296;
   reg _396297_396297 ; 
   reg __396297_396297;
   reg _396298_396298 ; 
   reg __396298_396298;
   reg _396299_396299 ; 
   reg __396299_396299;
   reg _396300_396300 ; 
   reg __396300_396300;
   reg _396301_396301 ; 
   reg __396301_396301;
   reg _396302_396302 ; 
   reg __396302_396302;
   reg _396303_396303 ; 
   reg __396303_396303;
   reg _396304_396304 ; 
   reg __396304_396304;
   reg _396305_396305 ; 
   reg __396305_396305;
   reg _396306_396306 ; 
   reg __396306_396306;
   reg _396307_396307 ; 
   reg __396307_396307;
   reg _396308_396308 ; 
   reg __396308_396308;
   reg _396309_396309 ; 
   reg __396309_396309;
   reg _396310_396310 ; 
   reg __396310_396310;
   reg _396311_396311 ; 
   reg __396311_396311;
   reg _396312_396312 ; 
   reg __396312_396312;
   reg _396313_396313 ; 
   reg __396313_396313;
   reg _396314_396314 ; 
   reg __396314_396314;
   reg _396315_396315 ; 
   reg __396315_396315;
   reg _396316_396316 ; 
   reg __396316_396316;
   reg _396317_396317 ; 
   reg __396317_396317;
   reg _396318_396318 ; 
   reg __396318_396318;
   reg _396319_396319 ; 
   reg __396319_396319;
   reg _396320_396320 ; 
   reg __396320_396320;
   reg _396321_396321 ; 
   reg __396321_396321;
   reg _396322_396322 ; 
   reg __396322_396322;
   reg _396323_396323 ; 
   reg __396323_396323;
   reg _396324_396324 ; 
   reg __396324_396324;
   reg _396325_396325 ; 
   reg __396325_396325;
   reg _396326_396326 ; 
   reg __396326_396326;
   reg _396327_396327 ; 
   reg __396327_396327;
   reg _396328_396328 ; 
   reg __396328_396328;
   reg _396329_396329 ; 
   reg __396329_396329;
   reg _396330_396330 ; 
   reg __396330_396330;
   reg _396331_396331 ; 
   reg __396331_396331;
   reg _396332_396332 ; 
   reg __396332_396332;
   reg _396333_396333 ; 
   reg __396333_396333;
   reg _396334_396334 ; 
   reg __396334_396334;
   reg _396335_396335 ; 
   reg __396335_396335;
   reg _396336_396336 ; 
   reg __396336_396336;
   reg _396337_396337 ; 
   reg __396337_396337;
   reg _396338_396338 ; 
   reg __396338_396338;
   reg _396339_396339 ; 
   reg __396339_396339;
   reg _396340_396340 ; 
   reg __396340_396340;
   reg _396341_396341 ; 
   reg __396341_396341;
   reg _396342_396342 ; 
   reg __396342_396342;
   reg _396343_396343 ; 
   reg __396343_396343;
   reg _396344_396344 ; 
   reg __396344_396344;
   reg _396345_396345 ; 
   reg __396345_396345;
   reg _396346_396346 ; 
   reg __396346_396346;
   reg _396347_396347 ; 
   reg __396347_396347;
   reg _396348_396348 ; 
   reg __396348_396348;
   reg _396349_396349 ; 
   reg __396349_396349;
   reg _396350_396350 ; 
   reg __396350_396350;
   reg _396351_396351 ; 
   reg __396351_396351;
   reg _396352_396352 ; 
   reg __396352_396352;
   reg _396353_396353 ; 
   reg __396353_396353;
   reg _396354_396354 ; 
   reg __396354_396354;
   reg _396355_396355 ; 
   reg __396355_396355;
   reg _396356_396356 ; 
   reg __396356_396356;
   reg _396357_396357 ; 
   reg __396357_396357;
   reg _396358_396358 ; 
   reg __396358_396358;
   reg _396359_396359 ; 
   reg __396359_396359;
   reg _396360_396360 ; 
   reg __396360_396360;
   reg _396361_396361 ; 
   reg __396361_396361;
   reg _396362_396362 ; 
   reg __396362_396362;
   reg _396363_396363 ; 
   reg __396363_396363;
   reg _396364_396364 ; 
   reg __396364_396364;
   reg _396365_396365 ; 
   reg __396365_396365;
   reg _396366_396366 ; 
   reg __396366_396366;
   reg _396367_396367 ; 
   reg __396367_396367;
   reg _396368_396368 ; 
   reg __396368_396368;
   reg _396369_396369 ; 
   reg __396369_396369;
   reg _396370_396370 ; 
   reg __396370_396370;
   reg _396371_396371 ; 
   reg __396371_396371;
   reg _396372_396372 ; 
   reg __396372_396372;
   reg _396373_396373 ; 
   reg __396373_396373;
   reg _396374_396374 ; 
   reg __396374_396374;
   reg _396375_396375 ; 
   reg __396375_396375;
   reg _396376_396376 ; 
   reg __396376_396376;
   reg _396377_396377 ; 
   reg __396377_396377;
   reg _396378_396378 ; 
   reg __396378_396378;
   reg _396379_396379 ; 
   reg __396379_396379;
   reg _396380_396380 ; 
   reg __396380_396380;
   reg _396381_396381 ; 
   reg __396381_396381;
   reg _396382_396382 ; 
   reg __396382_396382;
   reg _396383_396383 ; 
   reg __396383_396383;
   reg _396384_396384 ; 
   reg __396384_396384;
   reg _396385_396385 ; 
   reg __396385_396385;
   reg _396386_396386 ; 
   reg __396386_396386;
   reg _396387_396387 ; 
   reg __396387_396387;
   reg _396388_396388 ; 
   reg __396388_396388;
   reg _396389_396389 ; 
   reg __396389_396389;
   reg _396390_396390 ; 
   reg __396390_396390;
   reg _396391_396391 ; 
   reg __396391_396391;
   reg _396392_396392 ; 
   reg __396392_396392;
   reg _396393_396393 ; 
   reg __396393_396393;
   reg _396394_396394 ; 
   reg __396394_396394;
   reg _396395_396395 ; 
   reg __396395_396395;
   reg _396396_396396 ; 
   reg __396396_396396;
   reg _396397_396397 ; 
   reg __396397_396397;
   reg _396398_396398 ; 
   reg __396398_396398;
   reg _396399_396399 ; 
   reg __396399_396399;
   reg _396400_396400 ; 
   reg __396400_396400;
   reg _396401_396401 ; 
   reg __396401_396401;
   reg _396402_396402 ; 
   reg __396402_396402;
   reg _396403_396403 ; 
   reg __396403_396403;
   reg _396404_396404 ; 
   reg __396404_396404;
   reg _396405_396405 ; 
   reg __396405_396405;
   reg _396406_396406 ; 
   reg __396406_396406;
   reg _396407_396407 ; 
   reg __396407_396407;
   reg _396408_396408 ; 
   reg __396408_396408;
   reg _396409_396409 ; 
   reg __396409_396409;
   reg _396410_396410 ; 
   reg __396410_396410;
   reg _396411_396411 ; 
   reg __396411_396411;
   reg _396412_396412 ; 
   reg __396412_396412;
   reg _396413_396413 ; 
   reg __396413_396413;
   reg _396414_396414 ; 
   reg __396414_396414;
   reg _396415_396415 ; 
   reg __396415_396415;
   reg _396416_396416 ; 
   reg __396416_396416;
   reg _396417_396417 ; 
   reg __396417_396417;
   reg _396418_396418 ; 
   reg __396418_396418;
   reg _396419_396419 ; 
   reg __396419_396419;
   reg _396420_396420 ; 
   reg __396420_396420;
   reg _396421_396421 ; 
   reg __396421_396421;
   reg _396422_396422 ; 
   reg __396422_396422;
   reg _396423_396423 ; 
   reg __396423_396423;
   reg _396424_396424 ; 
   reg __396424_396424;
   reg _396425_396425 ; 
   reg __396425_396425;
   reg _396426_396426 ; 
   reg __396426_396426;
   reg _396427_396427 ; 
   reg __396427_396427;
   reg _396428_396428 ; 
   reg __396428_396428;
   reg _396429_396429 ; 
   reg __396429_396429;
   reg _396430_396430 ; 
   reg __396430_396430;
   reg _396431_396431 ; 
   reg __396431_396431;
   reg _396432_396432 ; 
   reg __396432_396432;
   reg _396433_396433 ; 
   reg __396433_396433;
   reg _396434_396434 ; 
   reg __396434_396434;
   reg _396435_396435 ; 
   reg __396435_396435;
   reg _396436_396436 ; 
   reg __396436_396436;
   reg _396437_396437 ; 
   reg __396437_396437;
   reg _396438_396438 ; 
   reg __396438_396438;
   reg _396439_396439 ; 
   reg __396439_396439;
   reg _396440_396440 ; 
   reg __396440_396440;
   reg _396441_396441 ; 
   reg __396441_396441;
   reg _396442_396442 ; 
   reg __396442_396442;
   reg _396443_396443 ; 
   reg __396443_396443;
   reg _396444_396444 ; 
   reg __396444_396444;
   reg _396445_396445 ; 
   reg __396445_396445;
   reg _396446_396446 ; 
   reg __396446_396446;
   reg _396447_396447 ; 
   reg __396447_396447;
   reg _396448_396448 ; 
   reg __396448_396448;
   reg _396449_396449 ; 
   reg __396449_396449;
   reg _396450_396450 ; 
   reg __396450_396450;
   reg _396451_396451 ; 
   reg __396451_396451;
   reg _396452_396452 ; 
   reg __396452_396452;
   reg _396453_396453 ; 
   reg __396453_396453;
   reg _396454_396454 ; 
   reg __396454_396454;
   reg _396455_396455 ; 
   reg __396455_396455;
   reg _396456_396456 ; 
   reg __396456_396456;
   reg _396457_396457 ; 
   reg __396457_396457;
   reg _396458_396458 ; 
   reg __396458_396458;
   reg _396459_396459 ; 
   reg __396459_396459;
   reg _396460_396460 ; 
   reg __396460_396460;
   reg _396461_396461 ; 
   reg __396461_396461;
   reg _396462_396462 ; 
   reg __396462_396462;
   reg _396463_396463 ; 
   reg __396463_396463;
   reg _396464_396464 ; 
   reg __396464_396464;
   reg _396465_396465 ; 
   reg __396465_396465;
   reg _396466_396466 ; 
   reg __396466_396466;
   reg _396467_396467 ; 
   reg __396467_396467;
   reg _396468_396468 ; 
   reg __396468_396468;
   reg _396469_396469 ; 
   reg __396469_396469;
   reg _396470_396470 ; 
   reg __396470_396470;
   reg _396471_396471 ; 
   reg __396471_396471;
   reg _396472_396472 ; 
   reg __396472_396472;
   reg _396473_396473 ; 
   reg __396473_396473;
   reg _396474_396474 ; 
   reg __396474_396474;
   reg _396475_396475 ; 
   reg __396475_396475;
   reg _396476_396476 ; 
   reg __396476_396476;
   reg _396477_396477 ; 
   reg __396477_396477;
   reg _396478_396478 ; 
   reg __396478_396478;
   reg _396479_396479 ; 
   reg __396479_396479;
   reg _396480_396480 ; 
   reg __396480_396480;
   reg _396481_396481 ; 
   reg __396481_396481;
   reg _396482_396482 ; 
   reg __396482_396482;
   reg _396483_396483 ; 
   reg __396483_396483;
   reg _396484_396484 ; 
   reg __396484_396484;
   reg _396485_396485 ; 
   reg __396485_396485;
   reg _396486_396486 ; 
   reg __396486_396486;
   reg _396487_396487 ; 
   reg __396487_396487;
   reg _396488_396488 ; 
   reg __396488_396488;
   reg _396489_396489 ; 
   reg __396489_396489;
   reg _396490_396490 ; 
   reg __396490_396490;
   reg _396491_396491 ; 
   reg __396491_396491;
   reg _396492_396492 ; 
   reg __396492_396492;
   reg _396493_396493 ; 
   reg __396493_396493;
   reg _396494_396494 ; 
   reg __396494_396494;
   reg _396495_396495 ; 
   reg __396495_396495;
   reg _396496_396496 ; 
   reg __396496_396496;
   reg _396497_396497 ; 
   reg __396497_396497;
   reg _396498_396498 ; 
   reg __396498_396498;
   reg _396499_396499 ; 
   reg __396499_396499;
   reg _396500_396500 ; 
   reg __396500_396500;
   reg _396501_396501 ; 
   reg __396501_396501;
   reg _396502_396502 ; 
   reg __396502_396502;
   reg _396503_396503 ; 
   reg __396503_396503;
   reg _396504_396504 ; 
   reg __396504_396504;
   reg _396505_396505 ; 
   reg __396505_396505;
   reg _396506_396506 ; 
   reg __396506_396506;
   reg _396507_396507 ; 
   reg __396507_396507;
   reg _396508_396508 ; 
   reg __396508_396508;
   reg _396509_396509 ; 
   reg __396509_396509;
   reg _396510_396510 ; 
   reg __396510_396510;
   reg _396511_396511 ; 
   reg __396511_396511;
   reg _396512_396512 ; 
   reg __396512_396512;
   reg _396513_396513 ; 
   reg __396513_396513;
   reg _396514_396514 ; 
   reg __396514_396514;
   reg _396515_396515 ; 
   reg __396515_396515;
   reg _396516_396516 ; 
   reg __396516_396516;
   reg _396517_396517 ; 
   reg __396517_396517;
   reg _396518_396518 ; 
   reg __396518_396518;
   reg _396519_396519 ; 
   reg __396519_396519;
   reg _396520_396520 ; 
   reg __396520_396520;
   reg _396521_396521 ; 
   reg __396521_396521;
   reg _396522_396522 ; 
   reg __396522_396522;
   reg _396523_396523 ; 
   reg __396523_396523;
   reg _396524_396524 ; 
   reg __396524_396524;
   reg _396525_396525 ; 
   reg __396525_396525;
   reg _396526_396526 ; 
   reg __396526_396526;
   reg _396527_396527 ; 
   reg __396527_396527;
   reg _396528_396528 ; 
   reg __396528_396528;
   reg _396529_396529 ; 
   reg __396529_396529;
   reg _396530_396530 ; 
   reg __396530_396530;
   reg _396531_396531 ; 
   reg __396531_396531;
   reg _396532_396532 ; 
   reg __396532_396532;
   reg _396533_396533 ; 
   reg __396533_396533;
   reg _396534_396534 ; 
   reg __396534_396534;
   reg _396535_396535 ; 
   reg __396535_396535;
   reg _396536_396536 ; 
   reg __396536_396536;
   reg _396537_396537 ; 
   reg __396537_396537;
   reg _396538_396538 ; 
   reg __396538_396538;
   reg _396539_396539 ; 
   reg __396539_396539;
   reg _396540_396540 ; 
   reg __396540_396540;
   reg _396541_396541 ; 
   reg __396541_396541;
   reg _396542_396542 ; 
   reg __396542_396542;
   reg _396543_396543 ; 
   reg __396543_396543;
   reg _396544_396544 ; 
   reg __396544_396544;
   reg _396545_396545 ; 
   reg __396545_396545;
   reg _396546_396546 ; 
   reg __396546_396546;
   reg _396547_396547 ; 
   reg __396547_396547;
   reg _396548_396548 ; 
   reg __396548_396548;
   reg _396549_396549 ; 
   reg __396549_396549;
   reg _396550_396550 ; 
   reg __396550_396550;
   reg _396551_396551 ; 
   reg __396551_396551;
   reg _396552_396552 ; 
   reg __396552_396552;
   reg _396553_396553 ; 
   reg __396553_396553;
   reg _396554_396554 ; 
   reg __396554_396554;
   reg _396555_396555 ; 
   reg __396555_396555;
   reg _396556_396556 ; 
   reg __396556_396556;
   reg _396557_396557 ; 
   reg __396557_396557;
   reg _396558_396558 ; 
   reg __396558_396558;
   reg _396559_396559 ; 
   reg __396559_396559;
   reg _396560_396560 ; 
   reg __396560_396560;
   reg _396561_396561 ; 
   reg __396561_396561;
   reg _396562_396562 ; 
   reg __396562_396562;
   reg _396563_396563 ; 
   reg __396563_396563;
   reg _396564_396564 ; 
   reg __396564_396564;
   reg _396565_396565 ; 
   reg __396565_396565;
   reg _396566_396566 ; 
   reg __396566_396566;
   reg _396567_396567 ; 
   reg __396567_396567;
   reg _396568_396568 ; 
   reg __396568_396568;
   reg _396569_396569 ; 
   reg __396569_396569;
   reg _396570_396570 ; 
   reg __396570_396570;
   reg _396571_396571 ; 
   reg __396571_396571;
   reg _396572_396572 ; 
   reg __396572_396572;
   reg _396573_396573 ; 
   reg __396573_396573;
   reg _396574_396574 ; 
   reg __396574_396574;
   reg _396575_396575 ; 
   reg __396575_396575;
   reg _396576_396576 ; 
   reg __396576_396576;
   reg _396577_396577 ; 
   reg __396577_396577;
   reg _396578_396578 ; 
   reg __396578_396578;
   reg _396579_396579 ; 
   reg __396579_396579;
   reg _396580_396580 ; 
   reg __396580_396580;
   reg _396581_396581 ; 
   reg __396581_396581;
   reg _396582_396582 ; 
   reg __396582_396582;
   reg _396583_396583 ; 
   reg __396583_396583;
   reg _396584_396584 ; 
   reg __396584_396584;
   reg _396585_396585 ; 
   reg __396585_396585;
   reg _396586_396586 ; 
   reg __396586_396586;
   reg _396587_396587 ; 
   reg __396587_396587;
   reg _396588_396588 ; 
   reg __396588_396588;
   reg _396589_396589 ; 
   reg __396589_396589;
   reg _396590_396590 ; 
   reg __396590_396590;
   reg _396591_396591 ; 
   reg __396591_396591;
   reg _396592_396592 ; 
   reg __396592_396592;
   reg _396593_396593 ; 
   reg __396593_396593;
   reg _396594_396594 ; 
   reg __396594_396594;
   reg _396595_396595 ; 
   reg __396595_396595;
   reg _396596_396596 ; 
   reg __396596_396596;
   reg _396597_396597 ; 
   reg __396597_396597;
   reg _396598_396598 ; 
   reg __396598_396598;
   reg _396599_396599 ; 
   reg __396599_396599;
   reg _396600_396600 ; 
   reg __396600_396600;
   reg _396601_396601 ; 
   reg __396601_396601;
   reg _396602_396602 ; 
   reg __396602_396602;
   reg _396603_396603 ; 
   reg __396603_396603;
   reg _396604_396604 ; 
   reg __396604_396604;
   reg _396605_396605 ; 
   reg __396605_396605;
   reg _396606_396606 ; 
   reg __396606_396606;
   reg _396607_396607 ; 
   reg __396607_396607;
   reg _396608_396608 ; 
   reg __396608_396608;
   reg _396609_396609 ; 
   reg __396609_396609;
   reg _396610_396610 ; 
   reg __396610_396610;
   reg _396611_396611 ; 
   reg __396611_396611;
   reg _396612_396612 ; 
   reg __396612_396612;
   reg _396613_396613 ; 
   reg __396613_396613;
   reg _396614_396614 ; 
   reg __396614_396614;
   reg _396615_396615 ; 
   reg __396615_396615;
   reg _396616_396616 ; 
   reg __396616_396616;
   reg _396617_396617 ; 
   reg __396617_396617;
   reg _396618_396618 ; 
   reg __396618_396618;
   reg _396619_396619 ; 
   reg __396619_396619;
   reg _396620_396620 ; 
   reg __396620_396620;
   reg _396621_396621 ; 
   reg __396621_396621;
   reg _396622_396622 ; 
   reg __396622_396622;
   reg _396623_396623 ; 
   reg __396623_396623;
   reg _396624_396624 ; 
   reg __396624_396624;
   reg _396625_396625 ; 
   reg __396625_396625;
   reg _396626_396626 ; 
   reg __396626_396626;
   reg _396627_396627 ; 
   reg __396627_396627;
   reg _396628_396628 ; 
   reg __396628_396628;
   reg _396629_396629 ; 
   reg __396629_396629;
   reg _396630_396630 ; 
   reg __396630_396630;
   reg _396631_396631 ; 
   reg __396631_396631;
   reg _396632_396632 ; 
   reg __396632_396632;
   reg _396633_396633 ; 
   reg __396633_396633;
   reg _396634_396634 ; 
   reg __396634_396634;
   reg _396635_396635 ; 
   reg __396635_396635;
   reg _396636_396636 ; 
   reg __396636_396636;
   reg _396637_396637 ; 
   reg __396637_396637;
   reg _396638_396638 ; 
   reg __396638_396638;
   reg _396639_396639 ; 
   reg __396639_396639;
   reg _396640_396640 ; 
   reg __396640_396640;
   reg _396641_396641 ; 
   reg __396641_396641;
   reg _396642_396642 ; 
   reg __396642_396642;
   reg _396643_396643 ; 
   reg __396643_396643;
   reg _396644_396644 ; 
   reg __396644_396644;
   reg _396645_396645 ; 
   reg __396645_396645;
   reg _396646_396646 ; 
   reg __396646_396646;
   reg _396647_396647 ; 
   reg __396647_396647;
   reg _396648_396648 ; 
   reg __396648_396648;
   reg _396649_396649 ; 
   reg __396649_396649;
   reg _396650_396650 ; 
   reg __396650_396650;
   reg _396651_396651 ; 
   reg __396651_396651;
   reg _396652_396652 ; 
   reg __396652_396652;
   reg _396653_396653 ; 
   reg __396653_396653;
   reg _396654_396654 ; 
   reg __396654_396654;
   reg _396655_396655 ; 
   reg __396655_396655;
   reg _396656_396656 ; 
   reg __396656_396656;
   reg _396657_396657 ; 
   reg __396657_396657;
   reg _396658_396658 ; 
   reg __396658_396658;
   reg _396659_396659 ; 
   reg __396659_396659;
   reg _396660_396660 ; 
   reg __396660_396660;
   reg _396661_396661 ; 
   reg __396661_396661;
   reg _396662_396662 ; 
   reg __396662_396662;
   reg _396663_396663 ; 
   reg __396663_396663;
   reg _396664_396664 ; 
   reg __396664_396664;
   reg _396665_396665 ; 
   reg __396665_396665;
   reg _396666_396666 ; 
   reg __396666_396666;
   reg _396667_396667 ; 
   reg __396667_396667;
   reg _396668_396668 ; 
   reg __396668_396668;
   reg _396669_396669 ; 
   reg __396669_396669;
   reg _396670_396670 ; 
   reg __396670_396670;
   reg _396671_396671 ; 
   reg __396671_396671;
   reg _396672_396672 ; 
   reg __396672_396672;
   reg _396673_396673 ; 
   reg __396673_396673;
   reg _396674_396674 ; 
   reg __396674_396674;
   reg _396675_396675 ; 
   reg __396675_396675;
   reg _396676_396676 ; 
   reg __396676_396676;
   reg _396677_396677 ; 
   reg __396677_396677;
   reg _396678_396678 ; 
   reg __396678_396678;
   reg _396679_396679 ; 
   reg __396679_396679;
   reg _396680_396680 ; 
   reg __396680_396680;
   reg _396681_396681 ; 
   reg __396681_396681;
   reg _396682_396682 ; 
   reg __396682_396682;
   reg _396683_396683 ; 
   reg __396683_396683;
   reg _396684_396684 ; 
   reg __396684_396684;
   reg _396685_396685 ; 
   reg __396685_396685;
   reg _396686_396686 ; 
   reg __396686_396686;
   reg _396687_396687 ; 
   reg __396687_396687;
   reg _396688_396688 ; 
   reg __396688_396688;
   reg _396689_396689 ; 
   reg __396689_396689;
   reg _396690_396690 ; 
   reg __396690_396690;
   reg _396691_396691 ; 
   reg __396691_396691;
   reg _396692_396692 ; 
   reg __396692_396692;
   reg _396693_396693 ; 
   reg __396693_396693;
   reg _396694_396694 ; 
   reg __396694_396694;
   reg _396695_396695 ; 
   reg __396695_396695;
   reg _396696_396696 ; 
   reg __396696_396696;
   reg _396697_396697 ; 
   reg __396697_396697;
   reg _396698_396698 ; 
   reg __396698_396698;
   reg _396699_396699 ; 
   reg __396699_396699;
   reg _396700_396700 ; 
   reg __396700_396700;
   reg _396701_396701 ; 
   reg __396701_396701;
   reg _396702_396702 ; 
   reg __396702_396702;
   reg _396703_396703 ; 
   reg __396703_396703;
   reg _396704_396704 ; 
   reg __396704_396704;
   reg _396705_396705 ; 
   reg __396705_396705;
   reg _396706_396706 ; 
   reg __396706_396706;
   reg _396707_396707 ; 
   reg __396707_396707;
   reg _396708_396708 ; 
   reg __396708_396708;
   reg _396709_396709 ; 
   reg __396709_396709;
   reg _396710_396710 ; 
   reg __396710_396710;
   reg _396711_396711 ; 
   reg __396711_396711;
   reg _396712_396712 ; 
   reg __396712_396712;
   reg _396713_396713 ; 
   reg __396713_396713;
   reg _396714_396714 ; 
   reg __396714_396714;
   reg _396715_396715 ; 
   reg __396715_396715;
   reg _396716_396716 ; 
   reg __396716_396716;
   reg _396717_396717 ; 
   reg __396717_396717;
   reg _396718_396718 ; 
   reg __396718_396718;
   reg _396719_396719 ; 
   reg __396719_396719;
   reg _396720_396720 ; 
   reg __396720_396720;
   reg _396721_396721 ; 
   reg __396721_396721;
   reg _396722_396722 ; 
   reg __396722_396722;
   reg _396723_396723 ; 
   reg __396723_396723;
   reg _396724_396724 ; 
   reg __396724_396724;
   reg _396725_396725 ; 
   reg __396725_396725;
   reg _396726_396726 ; 
   reg __396726_396726;
   reg _396727_396727 ; 
   reg __396727_396727;
   reg _396728_396728 ; 
   reg __396728_396728;
   reg _396729_396729 ; 
   reg __396729_396729;
   reg _396730_396730 ; 
   reg __396730_396730;
   reg _396731_396731 ; 
   reg __396731_396731;
   reg _396732_396732 ; 
   reg __396732_396732;
   reg _396733_396733 ; 
   reg __396733_396733;
   reg _396734_396734 ; 
   reg __396734_396734;
   reg _396735_396735 ; 
   reg __396735_396735;
   reg _396736_396736 ; 
   reg __396736_396736;
   reg _396737_396737 ; 
   reg __396737_396737;
   reg _396738_396738 ; 
   reg __396738_396738;
   reg _396739_396739 ; 
   reg __396739_396739;
   reg _396740_396740 ; 
   reg __396740_396740;
   reg _396741_396741 ; 
   reg __396741_396741;
   reg _396742_396742 ; 
   reg __396742_396742;
   reg _396743_396743 ; 
   reg __396743_396743;
   reg _396744_396744 ; 
   reg __396744_396744;
   reg _396745_396745 ; 
   reg __396745_396745;
   reg _396746_396746 ; 
   reg __396746_396746;
   reg _396747_396747 ; 
   reg __396747_396747;
   reg _396748_396748 ; 
   reg __396748_396748;
   reg _396749_396749 ; 
   reg __396749_396749;
   reg _396750_396750 ; 
   reg __396750_396750;
   reg _396751_396751 ; 
   reg __396751_396751;
   reg _396752_396752 ; 
   reg __396752_396752;
   reg _396753_396753 ; 
   reg __396753_396753;
   reg _396754_396754 ; 
   reg __396754_396754;
   reg _396755_396755 ; 
   reg __396755_396755;
   reg _396756_396756 ; 
   reg __396756_396756;
   reg _396757_396757 ; 
   reg __396757_396757;
   reg _396758_396758 ; 
   reg __396758_396758;
   reg _396759_396759 ; 
   reg __396759_396759;
   reg _396760_396760 ; 
   reg __396760_396760;
   reg _396761_396761 ; 
   reg __396761_396761;
   reg _396762_396762 ; 
   reg __396762_396762;
   reg _396763_396763 ; 
   reg __396763_396763;
   reg _396764_396764 ; 
   reg __396764_396764;
   reg _396765_396765 ; 
   reg __396765_396765;
   reg _396766_396766 ; 
   reg __396766_396766;
   reg _396767_396767 ; 
   reg __396767_396767;
   reg _396768_396768 ; 
   reg __396768_396768;
   reg _396769_396769 ; 
   reg __396769_396769;
   reg _396770_396770 ; 
   reg __396770_396770;
   reg _396771_396771 ; 
   reg __396771_396771;
   reg _396772_396772 ; 
   reg __396772_396772;
   reg _396773_396773 ; 
   reg __396773_396773;
   reg _396774_396774 ; 
   reg __396774_396774;
   reg _396775_396775 ; 
   reg __396775_396775;
   reg _396776_396776 ; 
   reg __396776_396776;
   reg _396777_396777 ; 
   reg __396777_396777;
   reg _396778_396778 ; 
   reg __396778_396778;
   reg _396779_396779 ; 
   reg __396779_396779;
   reg _396780_396780 ; 
   reg __396780_396780;
   reg _396781_396781 ; 
   reg __396781_396781;
   reg _396782_396782 ; 
   reg __396782_396782;
   reg _396783_396783 ; 
   reg __396783_396783;
   reg _396784_396784 ; 
   reg __396784_396784;
   reg _396785_396785 ; 
   reg __396785_396785;
   reg _396786_396786 ; 
   reg __396786_396786;
   reg _396787_396787 ; 
   reg __396787_396787;
   reg _396788_396788 ; 
   reg __396788_396788;
   reg _396789_396789 ; 
   reg __396789_396789;
   reg _396790_396790 ; 
   reg __396790_396790;
   reg _396791_396791 ; 
   reg __396791_396791;
   reg _396792_396792 ; 
   reg __396792_396792;
   reg _396793_396793 ; 
   reg __396793_396793;
   reg _396794_396794 ; 
   reg __396794_396794;
   reg _396795_396795 ; 
   reg __396795_396795;
   reg _396796_396796 ; 
   reg __396796_396796;
   reg _396797_396797 ; 
   reg __396797_396797;
   reg _396798_396798 ; 
   reg __396798_396798;
   reg _396799_396799 ; 
   reg __396799_396799;
   reg _396800_396800 ; 
   reg __396800_396800;
   reg _396801_396801 ; 
   reg __396801_396801;
   reg _396802_396802 ; 
   reg __396802_396802;
   reg _396803_396803 ; 
   reg __396803_396803;
   reg _396804_396804 ; 
   reg __396804_396804;
   reg _396805_396805 ; 
   reg __396805_396805;
   reg _396806_396806 ; 
   reg __396806_396806;
   reg _396807_396807 ; 
   reg __396807_396807;
   reg _396808_396808 ; 
   reg __396808_396808;
   reg _396809_396809 ; 
   reg __396809_396809;
   reg _396810_396810 ; 
   reg __396810_396810;
   reg _396811_396811 ; 
   reg __396811_396811;
   reg _396812_396812 ; 
   reg __396812_396812;
   reg _396813_396813 ; 
   reg __396813_396813;
   reg _396814_396814 ; 
   reg __396814_396814;
   reg _396815_396815 ; 
   reg __396815_396815;
   reg _396816_396816 ; 
   reg __396816_396816;
   reg _396817_396817 ; 
   reg __396817_396817;
   reg _396818_396818 ; 
   reg __396818_396818;
   reg _396819_396819 ; 
   reg __396819_396819;
   reg _396820_396820 ; 
   reg __396820_396820;
   reg _396821_396821 ; 
   reg __396821_396821;
   reg _396822_396822 ; 
   reg __396822_396822;
   reg _396823_396823 ; 
   reg __396823_396823;
   reg _396824_396824 ; 
   reg __396824_396824;
   reg _396825_396825 ; 
   reg __396825_396825;
   reg _396826_396826 ; 
   reg __396826_396826;
   reg _396827_396827 ; 
   reg __396827_396827;
   reg _396828_396828 ; 
   reg __396828_396828;
   reg _396829_396829 ; 
   reg __396829_396829;
   reg _396830_396830 ; 
   reg __396830_396830;
   reg _396831_396831 ; 
   reg __396831_396831;
   reg _396832_396832 ; 
   reg __396832_396832;
   reg _396833_396833 ; 
   reg __396833_396833;
   reg _396834_396834 ; 
   reg __396834_396834;
   reg _396835_396835 ; 
   reg __396835_396835;
   reg _396836_396836 ; 
   reg __396836_396836;
   reg _396837_396837 ; 
   reg __396837_396837;
   reg _396838_396838 ; 
   reg __396838_396838;
   reg _396839_396839 ; 
   reg __396839_396839;
   reg _396840_396840 ; 
   reg __396840_396840;
   reg _396841_396841 ; 
   reg __396841_396841;
   reg _396842_396842 ; 
   reg __396842_396842;
   reg _396843_396843 ; 
   reg __396843_396843;
   reg _396844_396844 ; 
   reg __396844_396844;
   reg _396845_396845 ; 
   reg __396845_396845;
   reg _396846_396846 ; 
   reg __396846_396846;
   reg _396847_396847 ; 
   reg __396847_396847;
   reg _396848_396848 ; 
   reg __396848_396848;
   reg _396849_396849 ; 
   reg __396849_396849;
   reg _396850_396850 ; 
   reg __396850_396850;
   reg _396851_396851 ; 
   reg __396851_396851;
   reg _396852_396852 ; 
   reg __396852_396852;
   reg _396853_396853 ; 
   reg __396853_396853;
   reg _396854_396854 ; 
   reg __396854_396854;
   reg _396855_396855 ; 
   reg __396855_396855;
   reg _396856_396856 ; 
   reg __396856_396856;
   reg _396857_396857 ; 
   reg __396857_396857;
   reg _396858_396858 ; 
   reg __396858_396858;
   reg _396859_396859 ; 
   reg __396859_396859;
   reg _396860_396860 ; 
   reg __396860_396860;
   reg _396861_396861 ; 
   reg __396861_396861;
   reg _396862_396862 ; 
   reg __396862_396862;
   reg _396863_396863 ; 
   reg __396863_396863;
   reg _396864_396864 ; 
   reg __396864_396864;
   reg _396865_396865 ; 
   reg __396865_396865;
   reg _396866_396866 ; 
   reg __396866_396866;
   reg _396867_396867 ; 
   reg __396867_396867;
   reg _396868_396868 ; 
   reg __396868_396868;
   reg _396869_396869 ; 
   reg __396869_396869;
   reg _396870_396870 ; 
   reg __396870_396870;
   reg _396871_396871 ; 
   reg __396871_396871;
   reg _396872_396872 ; 
   reg __396872_396872;
   reg _396873_396873 ; 
   reg __396873_396873;
   reg _396874_396874 ; 
   reg __396874_396874;
   reg _396875_396875 ; 
   reg __396875_396875;
   reg _396876_396876 ; 
   reg __396876_396876;
   reg _396877_396877 ; 
   reg __396877_396877;
   reg _396878_396878 ; 
   reg __396878_396878;
   reg _396879_396879 ; 
   reg __396879_396879;
   reg _396880_396880 ; 
   reg __396880_396880;
   reg _396881_396881 ; 
   reg __396881_396881;
   reg _396882_396882 ; 
   reg __396882_396882;
   reg _396883_396883 ; 
   reg __396883_396883;
   reg _396884_396884 ; 
   reg __396884_396884;
   reg _396885_396885 ; 
   reg __396885_396885;
   reg _396886_396886 ; 
   reg __396886_396886;
   reg _396887_396887 ; 
   reg __396887_396887;
   reg _396888_396888 ; 
   reg __396888_396888;
   reg _396889_396889 ; 
   reg __396889_396889;
   reg _396890_396890 ; 
   reg __396890_396890;
   reg _396891_396891 ; 
   reg __396891_396891;
   reg _396892_396892 ; 
   reg __396892_396892;
   reg _396893_396893 ; 
   reg __396893_396893;
   reg _396894_396894 ; 
   reg __396894_396894;
   reg _396895_396895 ; 
   reg __396895_396895;
   reg _396896_396896 ; 
   reg __396896_396896;
   reg _396897_396897 ; 
   reg __396897_396897;
   reg _396898_396898 ; 
   reg __396898_396898;
   reg _396899_396899 ; 
   reg __396899_396899;
   reg _396900_396900 ; 
   reg __396900_396900;
   reg _396901_396901 ; 
   reg __396901_396901;
   reg _396902_396902 ; 
   reg __396902_396902;
   reg _396903_396903 ; 
   reg __396903_396903;
   reg _396904_396904 ; 
   reg __396904_396904;
   reg _396905_396905 ; 
   reg __396905_396905;
   reg _396906_396906 ; 
   reg __396906_396906;
   reg _396907_396907 ; 
   reg __396907_396907;
   reg _396908_396908 ; 
   reg __396908_396908;
   reg _396909_396909 ; 
   reg __396909_396909;
   reg _396910_396910 ; 
   reg __396910_396910;
   reg _396911_396911 ; 
   reg __396911_396911;
   reg _396912_396912 ; 
   reg __396912_396912;
   reg _396913_396913 ; 
   reg __396913_396913;
   reg _396914_396914 ; 
   reg __396914_396914;
   reg _396915_396915 ; 
   reg __396915_396915;
   reg _396916_396916 ; 
   reg __396916_396916;
   reg _396917_396917 ; 
   reg __396917_396917;
   reg _396918_396918 ; 
   reg __396918_396918;
   reg _396919_396919 ; 
   reg __396919_396919;
   reg _396920_396920 ; 
   reg __396920_396920;
   reg _396921_396921 ; 
   reg __396921_396921;
   reg _396922_396922 ; 
   reg __396922_396922;
   reg _396923_396923 ; 
   reg __396923_396923;
   reg _396924_396924 ; 
   reg __396924_396924;
   reg _396925_396925 ; 
   reg __396925_396925;
   reg _396926_396926 ; 
   reg __396926_396926;
   reg _396927_396927 ; 
   reg __396927_396927;
   reg _396928_396928 ; 
   reg __396928_396928;
   reg _396929_396929 ; 
   reg __396929_396929;
   reg _396930_396930 ; 
   reg __396930_396930;
   reg _396931_396931 ; 
   reg __396931_396931;
   reg _396932_396932 ; 
   reg __396932_396932;
   reg _396933_396933 ; 
   reg __396933_396933;
   reg _396934_396934 ; 
   reg __396934_396934;
   reg _396935_396935 ; 
   reg __396935_396935;
   reg _396936_396936 ; 
   reg __396936_396936;
   reg _396937_396937 ; 
   reg __396937_396937;
   reg _396938_396938 ; 
   reg __396938_396938;
   reg _396939_396939 ; 
   reg __396939_396939;
   reg _396940_396940 ; 
   reg __396940_396940;
   reg _396941_396941 ; 
   reg __396941_396941;
   reg _396942_396942 ; 
   reg __396942_396942;
   reg _396943_396943 ; 
   reg __396943_396943;
   reg _396944_396944 ; 
   reg __396944_396944;
   reg _396945_396945 ; 
   reg __396945_396945;
   reg _396946_396946 ; 
   reg __396946_396946;
   reg _396947_396947 ; 
   reg __396947_396947;
   reg _396948_396948 ; 
   reg __396948_396948;
   reg _396949_396949 ; 
   reg __396949_396949;
   reg _396950_396950 ; 
   reg __396950_396950;
   reg _396951_396951 ; 
   reg __396951_396951;
   reg _396952_396952 ; 
   reg __396952_396952;
   reg _396953_396953 ; 
   reg __396953_396953;
   reg _396954_396954 ; 
   reg __396954_396954;
   reg _396955_396955 ; 
   reg __396955_396955;
   reg _396956_396956 ; 
   reg __396956_396956;
   reg _396957_396957 ; 
   reg __396957_396957;
   reg _396958_396958 ; 
   reg __396958_396958;
   reg _396959_396959 ; 
   reg __396959_396959;
   reg _396960_396960 ; 
   reg __396960_396960;
   reg _396961_396961 ; 
   reg __396961_396961;
   reg _396962_396962 ; 
   reg __396962_396962;
   reg _396963_396963 ; 
   reg __396963_396963;
   reg _396964_396964 ; 
   reg __396964_396964;
   reg _396965_396965 ; 
   reg __396965_396965;
   reg _396966_396966 ; 
   reg __396966_396966;
   reg _396967_396967 ; 
   reg __396967_396967;
   reg _396968_396968 ; 
   reg __396968_396968;
   reg _396969_396969 ; 
   reg __396969_396969;
   reg _396970_396970 ; 
   reg __396970_396970;
   reg _396971_396971 ; 
   reg __396971_396971;
   reg _396972_396972 ; 
   reg __396972_396972;
   reg _396973_396973 ; 
   reg __396973_396973;
   reg _396974_396974 ; 
   reg __396974_396974;
   reg _396975_396975 ; 
   reg __396975_396975;
   reg _396976_396976 ; 
   reg __396976_396976;
   reg _396977_396977 ; 
   reg __396977_396977;
   reg _396978_396978 ; 
   reg __396978_396978;
   reg _396979_396979 ; 
   reg __396979_396979;
   reg _396980_396980 ; 
   reg __396980_396980;
   reg _396981_396981 ; 
   reg __396981_396981;
   reg _396982_396982 ; 
   reg __396982_396982;
   reg _396983_396983 ; 
   reg __396983_396983;
   reg _396984_396984 ; 
   reg __396984_396984;
   reg _396985_396985 ; 
   reg __396985_396985;
   reg _396986_396986 ; 
   reg __396986_396986;
   reg _396987_396987 ; 
   reg __396987_396987;
   reg _396988_396988 ; 
   reg __396988_396988;
   reg _396989_396989 ; 
   reg __396989_396989;
   reg _396990_396990 ; 
   reg __396990_396990;
   reg _396991_396991 ; 
   reg __396991_396991;
   reg _396992_396992 ; 
   reg __396992_396992;
   reg _396993_396993 ; 
   reg __396993_396993;
   reg _396994_396994 ; 
   reg __396994_396994;
   reg _396995_396995 ; 
   reg __396995_396995;
   reg _396996_396996 ; 
   reg __396996_396996;
   reg _396997_396997 ; 
   reg __396997_396997;
   reg _396998_396998 ; 
   reg __396998_396998;
   reg _396999_396999 ; 
   reg __396999_396999;
   reg _397000_397000 ; 
   reg __397000_397000;
   reg _397001_397001 ; 
   reg __397001_397001;
   reg _397002_397002 ; 
   reg __397002_397002;
   reg _397003_397003 ; 
   reg __397003_397003;
   reg _397004_397004 ; 
   reg __397004_397004;
   reg _397005_397005 ; 
   reg __397005_397005;
   reg _397006_397006 ; 
   reg __397006_397006;
   reg _397007_397007 ; 
   reg __397007_397007;
   reg _397008_397008 ; 
   reg __397008_397008;
   reg _397009_397009 ; 
   reg __397009_397009;
   reg _397010_397010 ; 
   reg __397010_397010;
   reg _397011_397011 ; 
   reg __397011_397011;
   reg _397012_397012 ; 
   reg __397012_397012;
   reg _397013_397013 ; 
   reg __397013_397013;
   reg _397014_397014 ; 
   reg __397014_397014;
   reg _397015_397015 ; 
   reg __397015_397015;
   reg _397016_397016 ; 
   reg __397016_397016;
   reg _397017_397017 ; 
   reg __397017_397017;
   reg _397018_397018 ; 
   reg __397018_397018;
   reg _397019_397019 ; 
   reg __397019_397019;
   reg _397020_397020 ; 
   reg __397020_397020;
   reg _397021_397021 ; 
   reg __397021_397021;
   reg _397022_397022 ; 
   reg __397022_397022;
   reg _397023_397023 ; 
   reg __397023_397023;
   reg _397024_397024 ; 
   reg __397024_397024;
   reg _397025_397025 ; 
   reg __397025_397025;
   reg _397026_397026 ; 
   reg __397026_397026;
   reg _397027_397027 ; 
   reg __397027_397027;
   reg _397028_397028 ; 
   reg __397028_397028;
   reg _397029_397029 ; 
   reg __397029_397029;
   reg _397030_397030 ; 
   reg __397030_397030;
   reg _397031_397031 ; 
   reg __397031_397031;
   reg _397032_397032 ; 
   reg __397032_397032;
   reg _397033_397033 ; 
   reg __397033_397033;
   reg _397034_397034 ; 
   reg __397034_397034;
   reg _397035_397035 ; 
   reg __397035_397035;
   reg _397036_397036 ; 
   reg __397036_397036;
   reg _397037_397037 ; 
   reg __397037_397037;
   reg _397038_397038 ; 
   reg __397038_397038;
   reg _397039_397039 ; 
   reg __397039_397039;
   reg _397040_397040 ; 
   reg __397040_397040;
   reg _397041_397041 ; 
   reg __397041_397041;
   reg _397042_397042 ; 
   reg __397042_397042;
   reg _397043_397043 ; 
   reg __397043_397043;
   reg _397044_397044 ; 
   reg __397044_397044;
   reg _397045_397045 ; 
   reg __397045_397045;
   reg _397046_397046 ; 
   reg __397046_397046;
   reg _397047_397047 ; 
   reg __397047_397047;
   reg _397048_397048 ; 
   reg __397048_397048;
   reg _397049_397049 ; 
   reg __397049_397049;
   reg _397050_397050 ; 
   reg __397050_397050;
   reg _397051_397051 ; 
   reg __397051_397051;
   reg _397052_397052 ; 
   reg __397052_397052;
   reg _397053_397053 ; 
   reg __397053_397053;
   reg _397054_397054 ; 
   reg __397054_397054;
   reg _397055_397055 ; 
   reg __397055_397055;
   reg _397056_397056 ; 
   reg __397056_397056;
   reg _397057_397057 ; 
   reg __397057_397057;
   reg _397058_397058 ; 
   reg __397058_397058;
   reg _397059_397059 ; 
   reg __397059_397059;
   reg _397060_397060 ; 
   reg __397060_397060;
   reg _397061_397061 ; 
   reg __397061_397061;
   reg _397062_397062 ; 
   reg __397062_397062;
   reg _397063_397063 ; 
   reg __397063_397063;
   reg _397064_397064 ; 
   reg __397064_397064;
   reg _397065_397065 ; 
   reg __397065_397065;
   reg _397066_397066 ; 
   reg __397066_397066;
   reg _397067_397067 ; 
   reg __397067_397067;
   reg _397068_397068 ; 
   reg __397068_397068;
   reg _397069_397069 ; 
   reg __397069_397069;
   reg _397070_397070 ; 
   reg __397070_397070;
   reg _397071_397071 ; 
   reg __397071_397071;
   reg _397072_397072 ; 
   reg __397072_397072;
   reg _397073_397073 ; 
   reg __397073_397073;
   reg _397074_397074 ; 
   reg __397074_397074;
   reg _397075_397075 ; 
   reg __397075_397075;
   reg _397076_397076 ; 
   reg __397076_397076;
   reg _397077_397077 ; 
   reg __397077_397077;
   reg _397078_397078 ; 
   reg __397078_397078;
   reg _397079_397079 ; 
   reg __397079_397079;
   reg _397080_397080 ; 
   reg __397080_397080;
   reg _397081_397081 ; 
   reg __397081_397081;
   reg _397082_397082 ; 
   reg __397082_397082;
   reg _397083_397083 ; 
   reg __397083_397083;
   reg _397084_397084 ; 
   reg __397084_397084;
   reg _397085_397085 ; 
   reg __397085_397085;
   reg _397086_397086 ; 
   reg __397086_397086;
   reg _397087_397087 ; 
   reg __397087_397087;
   reg _397088_397088 ; 
   reg __397088_397088;
   reg _397089_397089 ; 
   reg __397089_397089;
   reg _397090_397090 ; 
   reg __397090_397090;
   reg _397091_397091 ; 
   reg __397091_397091;
   reg _397092_397092 ; 
   reg __397092_397092;
   reg _397093_397093 ; 
   reg __397093_397093;
   reg _397094_397094 ; 
   reg __397094_397094;
   reg _397095_397095 ; 
   reg __397095_397095;
   reg _397096_397096 ; 
   reg __397096_397096;
   reg _397097_397097 ; 
   reg __397097_397097;
   reg _397098_397098 ; 
   reg __397098_397098;
   reg _397099_397099 ; 
   reg __397099_397099;
   reg _397100_397100 ; 
   reg __397100_397100;
   reg _397101_397101 ; 
   reg __397101_397101;
   reg _397102_397102 ; 
   reg __397102_397102;
   reg _397103_397103 ; 
   reg __397103_397103;
   reg _397104_397104 ; 
   reg __397104_397104;
   reg _397105_397105 ; 
   reg __397105_397105;
   reg _397106_397106 ; 
   reg __397106_397106;
   reg _397107_397107 ; 
   reg __397107_397107;
   reg _397108_397108 ; 
   reg __397108_397108;
   reg _397109_397109 ; 
   reg __397109_397109;
   reg _397110_397110 ; 
   reg __397110_397110;
   reg _397111_397111 ; 
   reg __397111_397111;
   reg _397112_397112 ; 
   reg __397112_397112;
   reg _397113_397113 ; 
   reg __397113_397113;
   reg _397114_397114 ; 
   reg __397114_397114;
   reg _397115_397115 ; 
   reg __397115_397115;
   reg _397116_397116 ; 
   reg __397116_397116;
   reg _397117_397117 ; 
   reg __397117_397117;
   reg _397118_397118 ; 
   reg __397118_397118;
   reg _397119_397119 ; 
   reg __397119_397119;
   reg _397120_397120 ; 
   reg __397120_397120;
   reg _397121_397121 ; 
   reg __397121_397121;
   reg _397122_397122 ; 
   reg __397122_397122;
   reg _397123_397123 ; 
   reg __397123_397123;
   reg _397124_397124 ; 
   reg __397124_397124;
   reg _397125_397125 ; 
   reg __397125_397125;
   reg _397126_397126 ; 
   reg __397126_397126;
   reg _397127_397127 ; 
   reg __397127_397127;
   reg _397128_397128 ; 
   reg __397128_397128;
   reg _397129_397129 ; 
   reg __397129_397129;
   reg _397130_397130 ; 
   reg __397130_397130;
   reg _397131_397131 ; 
   reg __397131_397131;
   reg _397132_397132 ; 
   reg __397132_397132;
   reg _397133_397133 ; 
   reg __397133_397133;
   reg _397134_397134 ; 
   reg __397134_397134;
   reg _397135_397135 ; 
   reg __397135_397135;
   reg _397136_397136 ; 
   reg __397136_397136;
   reg _397137_397137 ; 
   reg __397137_397137;
   reg _397138_397138 ; 
   reg __397138_397138;
   reg _397139_397139 ; 
   reg __397139_397139;
   reg _397140_397140 ; 
   reg __397140_397140;
   reg _397141_397141 ; 
   reg __397141_397141;
   reg _397142_397142 ; 
   reg __397142_397142;
   reg _397143_397143 ; 
   reg __397143_397143;
   reg _397144_397144 ; 
   reg __397144_397144;
   reg _397145_397145 ; 
   reg __397145_397145;
   reg _397146_397146 ; 
   reg __397146_397146;
   reg _397147_397147 ; 
   reg __397147_397147;
   reg _397148_397148 ; 
   reg __397148_397148;
   reg _397149_397149 ; 
   reg __397149_397149;
   reg _397150_397150 ; 
   reg __397150_397150;
   reg _397151_397151 ; 
   reg __397151_397151;
   reg _397152_397152 ; 
   reg __397152_397152;
   reg _397153_397153 ; 
   reg __397153_397153;
   reg _397154_397154 ; 
   reg __397154_397154;
   reg _397155_397155 ; 
   reg __397155_397155;
   reg _397156_397156 ; 
   reg __397156_397156;
   reg _397157_397157 ; 
   reg __397157_397157;
   reg _397158_397158 ; 
   reg __397158_397158;
   reg _397159_397159 ; 
   reg __397159_397159;
   reg _397160_397160 ; 
   reg __397160_397160;
   reg _397161_397161 ; 
   reg __397161_397161;
   reg _397162_397162 ; 
   reg __397162_397162;
   reg _397163_397163 ; 
   reg __397163_397163;
   reg _397164_397164 ; 
   reg __397164_397164;
   reg _397165_397165 ; 
   reg __397165_397165;
   reg _397166_397166 ; 
   reg __397166_397166;
   reg _397167_397167 ; 
   reg __397167_397167;
   reg _397168_397168 ; 
   reg __397168_397168;
   reg _397169_397169 ; 
   reg __397169_397169;
   reg _397170_397170 ; 
   reg __397170_397170;
   reg _397171_397171 ; 
   reg __397171_397171;
   reg _397172_397172 ; 
   reg __397172_397172;
   reg _397173_397173 ; 
   reg __397173_397173;
   reg _397174_397174 ; 
   reg __397174_397174;
   reg _397175_397175 ; 
   reg __397175_397175;
   reg _397176_397176 ; 
   reg __397176_397176;
   reg _397177_397177 ; 
   reg __397177_397177;
   reg _397178_397178 ; 
   reg __397178_397178;
   reg _397179_397179 ; 
   reg __397179_397179;
   reg _397180_397180 ; 
   reg __397180_397180;
   reg _397181_397181 ; 
   reg __397181_397181;
   reg _397182_397182 ; 
   reg __397182_397182;
   reg _397183_397183 ; 
   reg __397183_397183;
   reg _397184_397184 ; 
   reg __397184_397184;
   reg _397185_397185 ; 
   reg __397185_397185;
   reg _397186_397186 ; 
   reg __397186_397186;
   reg _397187_397187 ; 
   reg __397187_397187;
   reg _397188_397188 ; 
   reg __397188_397188;
   reg _397189_397189 ; 
   reg __397189_397189;
   reg _397190_397190 ; 
   reg __397190_397190;
   reg _397191_397191 ; 
   reg __397191_397191;
   reg _397192_397192 ; 
   reg __397192_397192;
   reg _397193_397193 ; 
   reg __397193_397193;
   reg _397194_397194 ; 
   reg __397194_397194;
   reg _397195_397195 ; 
   reg __397195_397195;
   reg _397196_397196 ; 
   reg __397196_397196;
   reg _397197_397197 ; 
   reg __397197_397197;
   reg _397198_397198 ; 
   reg __397198_397198;
   reg _397199_397199 ; 
   reg __397199_397199;
   reg _397200_397200 ; 
   reg __397200_397200;
   reg _397201_397201 ; 
   reg __397201_397201;
   reg _397202_397202 ; 
   reg __397202_397202;
   reg _397203_397203 ; 
   reg __397203_397203;
   reg _397204_397204 ; 
   reg __397204_397204;
   reg _397205_397205 ; 
   reg __397205_397205;
   reg _397206_397206 ; 
   reg __397206_397206;
   reg _397207_397207 ; 
   reg __397207_397207;
   reg _397208_397208 ; 
   reg __397208_397208;
   reg _397209_397209 ; 
   reg __397209_397209;
   reg _397210_397210 ; 
   reg __397210_397210;
   reg _397211_397211 ; 
   reg __397211_397211;
   reg _397212_397212 ; 
   reg __397212_397212;
   reg _397213_397213 ; 
   reg __397213_397213;
   reg _397214_397214 ; 
   reg __397214_397214;
   reg _397215_397215 ; 
   reg __397215_397215;
   reg _397216_397216 ; 
   reg __397216_397216;
   reg _397217_397217 ; 
   reg __397217_397217;
   reg _397218_397218 ; 
   reg __397218_397218;
   reg _397219_397219 ; 
   reg __397219_397219;
   reg _397220_397220 ; 
   reg __397220_397220;
   reg _397221_397221 ; 
   reg __397221_397221;
   reg _397222_397222 ; 
   reg __397222_397222;
   reg _397223_397223 ; 
   reg __397223_397223;
   reg _397224_397224 ; 
   reg __397224_397224;
   reg _397225_397225 ; 
   reg __397225_397225;
   reg _397226_397226 ; 
   reg __397226_397226;
   reg _397227_397227 ; 
   reg __397227_397227;
   reg _397228_397228 ; 
   reg __397228_397228;
   reg _397229_397229 ; 
   reg __397229_397229;
   reg _397230_397230 ; 
   reg __397230_397230;
   reg _397231_397231 ; 
   reg __397231_397231;
   reg _397232_397232 ; 
   reg __397232_397232;
   reg _397233_397233 ; 
   reg __397233_397233;
   reg _397234_397234 ; 
   reg __397234_397234;
   reg _397235_397235 ; 
   reg __397235_397235;
   reg _397236_397236 ; 
   reg __397236_397236;
   reg _397237_397237 ; 
   reg __397237_397237;
   reg _397238_397238 ; 
   reg __397238_397238;
   reg _397239_397239 ; 
   reg __397239_397239;
   reg _397240_397240 ; 
   reg __397240_397240;
   reg _397241_397241 ; 
   reg __397241_397241;
   reg _397242_397242 ; 
   reg __397242_397242;
   reg _397243_397243 ; 
   reg __397243_397243;
   reg _397244_397244 ; 
   reg __397244_397244;
   reg _397245_397245 ; 
   reg __397245_397245;
   reg _397246_397246 ; 
   reg __397246_397246;
   reg _397247_397247 ; 
   reg __397247_397247;
   reg _397248_397248 ; 
   reg __397248_397248;
   reg _397249_397249 ; 
   reg __397249_397249;
   reg _397250_397250 ; 
   reg __397250_397250;
   reg _397251_397251 ; 
   reg __397251_397251;
   reg _397252_397252 ; 
   reg __397252_397252;
   reg _397253_397253 ; 
   reg __397253_397253;
   reg _397254_397254 ; 
   reg __397254_397254;
   reg _397255_397255 ; 
   reg __397255_397255;
   reg _397256_397256 ; 
   reg __397256_397256;
   reg _397257_397257 ; 
   reg __397257_397257;
   reg _397258_397258 ; 
   reg __397258_397258;
   reg _397259_397259 ; 
   reg __397259_397259;
   reg _397260_397260 ; 
   reg __397260_397260;
   reg _397261_397261 ; 
   reg __397261_397261;
   reg _397262_397262 ; 
   reg __397262_397262;
   reg _397263_397263 ; 
   reg __397263_397263;
   reg _397264_397264 ; 
   reg __397264_397264;
   reg _397265_397265 ; 
   reg __397265_397265;
   reg _397266_397266 ; 
   reg __397266_397266;
   reg _397267_397267 ; 
   reg __397267_397267;
   reg _397268_397268 ; 
   reg __397268_397268;
   reg _397269_397269 ; 
   reg __397269_397269;
   reg _397270_397270 ; 
   reg __397270_397270;
   reg _397271_397271 ; 
   reg __397271_397271;
   reg _397272_397272 ; 
   reg __397272_397272;
   reg _397273_397273 ; 
   reg __397273_397273;
   reg _397274_397274 ; 
   reg __397274_397274;
   reg _397275_397275 ; 
   reg __397275_397275;
   reg _397276_397276 ; 
   reg __397276_397276;
   reg _397277_397277 ; 
   reg __397277_397277;
   reg _397278_397278 ; 
   reg __397278_397278;
   reg _397279_397279 ; 
   reg __397279_397279;
   reg _397280_397280 ; 
   reg __397280_397280;
   reg _397281_397281 ; 
   reg __397281_397281;
   reg _397282_397282 ; 
   reg __397282_397282;
   reg _397283_397283 ; 
   reg __397283_397283;
   reg _397284_397284 ; 
   reg __397284_397284;
   reg _397285_397285 ; 
   reg __397285_397285;
   reg _397286_397286 ; 
   reg __397286_397286;
   reg _397287_397287 ; 
   reg __397287_397287;
   reg _397288_397288 ; 
   reg __397288_397288;
   reg _397289_397289 ; 
   reg __397289_397289;
   reg _397290_397290 ; 
   reg __397290_397290;
   reg _397291_397291 ; 
   reg __397291_397291;
   reg _397292_397292 ; 
   reg __397292_397292;
   reg _397293_397293 ; 
   reg __397293_397293;
   reg _397294_397294 ; 
   reg __397294_397294;
   reg _397295_397295 ; 
   reg __397295_397295;
   reg _397296_397296 ; 
   reg __397296_397296;
   reg _397297_397297 ; 
   reg __397297_397297;
   reg _397298_397298 ; 
   reg __397298_397298;
   reg _397299_397299 ; 
   reg __397299_397299;
   reg _397300_397300 ; 
   reg __397300_397300;
   reg _397301_397301 ; 
   reg __397301_397301;
   reg _397302_397302 ; 
   reg __397302_397302;
   reg _397303_397303 ; 
   reg __397303_397303;
   reg _397304_397304 ; 
   reg __397304_397304;
   reg _397305_397305 ; 
   reg __397305_397305;
   reg _397306_397306 ; 
   reg __397306_397306;
   reg _397307_397307 ; 
   reg __397307_397307;
   reg _397308_397308 ; 
   reg __397308_397308;
   reg _397309_397309 ; 
   reg __397309_397309;
   reg _397310_397310 ; 
   reg __397310_397310;
   reg _397311_397311 ; 
   reg __397311_397311;
   reg _397312_397312 ; 
   reg __397312_397312;
   reg _397313_397313 ; 
   reg __397313_397313;
   reg _397314_397314 ; 
   reg __397314_397314;
   reg _397315_397315 ; 
   reg __397315_397315;
   reg _397316_397316 ; 
   reg __397316_397316;
   reg _397317_397317 ; 
   reg __397317_397317;
   reg _397318_397318 ; 
   reg __397318_397318;
   reg _397319_397319 ; 
   reg __397319_397319;
   reg _397320_397320 ; 
   reg __397320_397320;
   reg _397321_397321 ; 
   reg __397321_397321;
   reg _397322_397322 ; 
   reg __397322_397322;
   reg _397323_397323 ; 
   reg __397323_397323;
   reg _397324_397324 ; 
   reg __397324_397324;
   reg _397325_397325 ; 
   reg __397325_397325;
   reg _397326_397326 ; 
   reg __397326_397326;
   reg _397327_397327 ; 
   reg __397327_397327;
   reg _397328_397328 ; 
   reg __397328_397328;
   reg _397329_397329 ; 
   reg __397329_397329;
   reg _397330_397330 ; 
   reg __397330_397330;
   reg _397331_397331 ; 
   reg __397331_397331;
   reg _397332_397332 ; 
   reg __397332_397332;
   reg _397333_397333 ; 
   reg __397333_397333;
   reg _397334_397334 ; 
   reg __397334_397334;
   reg _397335_397335 ; 
   reg __397335_397335;
   reg _397336_397336 ; 
   reg __397336_397336;
   reg _397337_397337 ; 
   reg __397337_397337;
   reg _397338_397338 ; 
   reg __397338_397338;
   reg _397339_397339 ; 
   reg __397339_397339;
   reg _397340_397340 ; 
   reg __397340_397340;
   reg _397341_397341 ; 
   reg __397341_397341;
   reg _397342_397342 ; 
   reg __397342_397342;
   reg _397343_397343 ; 
   reg __397343_397343;
   reg _397344_397344 ; 
   reg __397344_397344;
   reg _397345_397345 ; 
   reg __397345_397345;
   reg _397346_397346 ; 
   reg __397346_397346;
   reg _397347_397347 ; 
   reg __397347_397347;
   reg _397348_397348 ; 
   reg __397348_397348;
   reg _397349_397349 ; 
   reg __397349_397349;
   reg _397350_397350 ; 
   reg __397350_397350;
   reg _397351_397351 ; 
   reg __397351_397351;
   reg _397352_397352 ; 
   reg __397352_397352;
   reg _397353_397353 ; 
   reg __397353_397353;
   reg _397354_397354 ; 
   reg __397354_397354;
   reg _397355_397355 ; 
   reg __397355_397355;
   reg _397356_397356 ; 
   reg __397356_397356;
   reg _397357_397357 ; 
   reg __397357_397357;
   reg _397358_397358 ; 
   reg __397358_397358;
   reg _397359_397359 ; 
   reg __397359_397359;
   reg _397360_397360 ; 
   reg __397360_397360;
   reg _397361_397361 ; 
   reg __397361_397361;
   reg _397362_397362 ; 
   reg __397362_397362;
   reg _397363_397363 ; 
   reg __397363_397363;
   reg _397364_397364 ; 
   reg __397364_397364;
   reg _397365_397365 ; 
   reg __397365_397365;
   reg _397366_397366 ; 
   reg __397366_397366;
   reg _397367_397367 ; 
   reg __397367_397367;
   reg _397368_397368 ; 
   reg __397368_397368;
   reg _397369_397369 ; 
   reg __397369_397369;
   reg _397370_397370 ; 
   reg __397370_397370;
   reg _397371_397371 ; 
   reg __397371_397371;
   reg _397372_397372 ; 
   reg __397372_397372;
   reg _397373_397373 ; 
   reg __397373_397373;
   reg _397374_397374 ; 
   reg __397374_397374;
   reg _397375_397375 ; 
   reg __397375_397375;
   reg _397376_397376 ; 
   reg __397376_397376;
   reg _397377_397377 ; 
   reg __397377_397377;
   reg _397378_397378 ; 
   reg __397378_397378;
   reg _397379_397379 ; 
   reg __397379_397379;
   reg _397380_397380 ; 
   reg __397380_397380;
   reg _397381_397381 ; 
   reg __397381_397381;
   reg _397382_397382 ; 
   reg __397382_397382;
   reg _397383_397383 ; 
   reg __397383_397383;
   reg _397384_397384 ; 
   reg __397384_397384;
   reg _397385_397385 ; 
   reg __397385_397385;
   reg _397386_397386 ; 
   reg __397386_397386;
   reg _397387_397387 ; 
   reg __397387_397387;
   reg _397388_397388 ; 
   reg __397388_397388;
   reg _397389_397389 ; 
   reg __397389_397389;
   reg _397390_397390 ; 
   reg __397390_397390;
   reg _397391_397391 ; 
   reg __397391_397391;
   reg _397392_397392 ; 
   reg __397392_397392;
   reg _397393_397393 ; 
   reg __397393_397393;
   reg _397394_397394 ; 
   reg __397394_397394;
   reg _397395_397395 ; 
   reg __397395_397395;
   reg _397396_397396 ; 
   reg __397396_397396;
   reg _397397_397397 ; 
   reg __397397_397397;
   reg _397398_397398 ; 
   reg __397398_397398;
   reg _397399_397399 ; 
   reg __397399_397399;
   reg _397400_397400 ; 
   reg __397400_397400;
   reg _397401_397401 ; 
   reg __397401_397401;
   reg _397402_397402 ; 
   reg __397402_397402;
   reg _397403_397403 ; 
   reg __397403_397403;
   reg _397404_397404 ; 
   reg __397404_397404;
   reg _397405_397405 ; 
   reg __397405_397405;
   reg _397406_397406 ; 
   reg __397406_397406;
   reg _397407_397407 ; 
   reg __397407_397407;
   reg _397408_397408 ; 
   reg __397408_397408;
   reg _397409_397409 ; 
   reg __397409_397409;
   reg _397410_397410 ; 
   reg __397410_397410;
   reg _397411_397411 ; 
   reg __397411_397411;
   reg _397412_397412 ; 
   reg __397412_397412;
   reg _397413_397413 ; 
   reg __397413_397413;
   reg _397414_397414 ; 
   reg __397414_397414;
   reg _397415_397415 ; 
   reg __397415_397415;
   reg _397416_397416 ; 
   reg __397416_397416;
   reg _397417_397417 ; 
   reg __397417_397417;
   reg _397418_397418 ; 
   reg __397418_397418;
   reg _397419_397419 ; 
   reg __397419_397419;
   reg _397420_397420 ; 
   reg __397420_397420;
   reg _397421_397421 ; 
   reg __397421_397421;
   reg _397422_397422 ; 
   reg __397422_397422;
   reg _397423_397423 ; 
   reg __397423_397423;
   reg _397424_397424 ; 
   reg __397424_397424;
   reg _397425_397425 ; 
   reg __397425_397425;
   reg _397426_397426 ; 
   reg __397426_397426;
   reg _397427_397427 ; 
   reg __397427_397427;
   reg _397428_397428 ; 
   reg __397428_397428;
   reg _397429_397429 ; 
   reg __397429_397429;
   reg _397430_397430 ; 
   reg __397430_397430;
   reg _397431_397431 ; 
   reg __397431_397431;
   reg _397432_397432 ; 
   reg __397432_397432;
   reg _397433_397433 ; 
   reg __397433_397433;
   reg _397434_397434 ; 
   reg __397434_397434;
   reg _397435_397435 ; 
   reg __397435_397435;
   reg _397436_397436 ; 
   reg __397436_397436;
   reg _397437_397437 ; 
   reg __397437_397437;
   reg _397438_397438 ; 
   reg __397438_397438;
   reg _397439_397439 ; 
   reg __397439_397439;
   reg _397440_397440 ; 
   reg __397440_397440;
   reg _397441_397441 ; 
   reg __397441_397441;
   reg _397442_397442 ; 
   reg __397442_397442;
   reg _397443_397443 ; 
   reg __397443_397443;
   reg _397444_397444 ; 
   reg __397444_397444;
   reg _397445_397445 ; 
   reg __397445_397445;
   reg _397446_397446 ; 
   reg __397446_397446;
   reg _397447_397447 ; 
   reg __397447_397447;
   reg _397448_397448 ; 
   reg __397448_397448;
   reg _397449_397449 ; 
   reg __397449_397449;
   reg _397450_397450 ; 
   reg __397450_397450;
   reg _397451_397451 ; 
   reg __397451_397451;
   reg _397452_397452 ; 
   reg __397452_397452;
   reg _397453_397453 ; 
   reg __397453_397453;
   reg _397454_397454 ; 
   reg __397454_397454;
   reg _397455_397455 ; 
   reg __397455_397455;
   reg _397456_397456 ; 
   reg __397456_397456;
   reg _397457_397457 ; 
   reg __397457_397457;
   reg _397458_397458 ; 
   reg __397458_397458;
   reg _397459_397459 ; 
   reg __397459_397459;
   reg _397460_397460 ; 
   reg __397460_397460;
   reg _397461_397461 ; 
   reg __397461_397461;
   reg _397462_397462 ; 
   reg __397462_397462;
   reg _397463_397463 ; 
   reg __397463_397463;
   reg _397464_397464 ; 
   reg __397464_397464;
   reg _397465_397465 ; 
   reg __397465_397465;
   reg _397466_397466 ; 
   reg __397466_397466;
   reg _397467_397467 ; 
   reg __397467_397467;
   reg _397468_397468 ; 
   reg __397468_397468;
   reg _397469_397469 ; 
   reg __397469_397469;
   reg _397470_397470 ; 
   reg __397470_397470;
   reg _397471_397471 ; 
   reg __397471_397471;
   reg _397472_397472 ; 
   reg __397472_397472;
   reg _397473_397473 ; 
   reg __397473_397473;
   reg _397474_397474 ; 
   reg __397474_397474;
   reg _397475_397475 ; 
   reg __397475_397475;
   reg _397476_397476 ; 
   reg __397476_397476;
   reg _397477_397477 ; 
   reg __397477_397477;
   reg _397478_397478 ; 
   reg __397478_397478;
   reg _397479_397479 ; 
   reg __397479_397479;
   reg _397480_397480 ; 
   reg __397480_397480;
   reg _397481_397481 ; 
   reg __397481_397481;
   reg _397482_397482 ; 
   reg __397482_397482;
   reg _397483_397483 ; 
   reg __397483_397483;
   reg _397484_397484 ; 
   reg __397484_397484;
   reg _397485_397485 ; 
   reg __397485_397485;
   reg _397486_397486 ; 
   reg __397486_397486;
   reg _397487_397487 ; 
   reg __397487_397487;
   reg _397488_397488 ; 
   reg __397488_397488;
   reg _397489_397489 ; 
   reg __397489_397489;
   reg _397490_397490 ; 
   reg __397490_397490;
   reg _397491_397491 ; 
   reg __397491_397491;
   reg _397492_397492 ; 
   reg __397492_397492;
   reg _397493_397493 ; 
   reg __397493_397493;
   reg _397494_397494 ; 
   reg __397494_397494;
   reg _397495_397495 ; 
   reg __397495_397495;
   reg _397496_397496 ; 
   reg __397496_397496;
   reg _397497_397497 ; 
   reg __397497_397497;
   reg _397498_397498 ; 
   reg __397498_397498;
   reg _397499_397499 ; 
   reg __397499_397499;
   reg _397500_397500 ; 
   reg __397500_397500;
   reg _397501_397501 ; 
   reg __397501_397501;
   reg _397502_397502 ; 
   reg __397502_397502;
   reg _397503_397503 ; 
   reg __397503_397503;
   reg _397504_397504 ; 
   reg __397504_397504;
   reg _397505_397505 ; 
   reg __397505_397505;
   reg _397506_397506 ; 
   reg __397506_397506;
   reg _397507_397507 ; 
   reg __397507_397507;
   reg _397508_397508 ; 
   reg __397508_397508;
   reg _397509_397509 ; 
   reg __397509_397509;
   reg _397510_397510 ; 
   reg __397510_397510;
   reg _397511_397511 ; 
   reg __397511_397511;
   reg _397512_397512 ; 
   reg __397512_397512;
   reg _397513_397513 ; 
   reg __397513_397513;
   reg _397514_397514 ; 
   reg __397514_397514;
   reg _397515_397515 ; 
   reg __397515_397515;
   reg _397516_397516 ; 
   reg __397516_397516;
   reg _397517_397517 ; 
   reg __397517_397517;
   reg _397518_397518 ; 
   reg __397518_397518;
   reg _397519_397519 ; 
   reg __397519_397519;
   reg _397520_397520 ; 
   reg __397520_397520;
   reg _397521_397521 ; 
   reg __397521_397521;
   reg _397522_397522 ; 
   reg __397522_397522;
   reg _397523_397523 ; 
   reg __397523_397523;
   reg _397524_397524 ; 
   reg __397524_397524;
   reg _397525_397525 ; 
   reg __397525_397525;
   reg _397526_397526 ; 
   reg __397526_397526;
   reg _397527_397527 ; 
   reg __397527_397527;
   reg _397528_397528 ; 
   reg __397528_397528;
   reg _397529_397529 ; 
   reg __397529_397529;
   reg _397530_397530 ; 
   reg __397530_397530;
   reg _397531_397531 ; 
   reg __397531_397531;
   reg _397532_397532 ; 
   reg __397532_397532;
   reg _397533_397533 ; 
   reg __397533_397533;
   reg _397534_397534 ; 
   reg __397534_397534;
   reg _397535_397535 ; 
   reg __397535_397535;
   reg _397536_397536 ; 
   reg __397536_397536;
   reg _397537_397537 ; 
   reg __397537_397537;
   reg _397538_397538 ; 
   reg __397538_397538;
   reg _397539_397539 ; 
   reg __397539_397539;
   reg _397540_397540 ; 
   reg __397540_397540;
   reg _397541_397541 ; 
   reg __397541_397541;
   reg _397542_397542 ; 
   reg __397542_397542;
   reg _397543_397543 ; 
   reg __397543_397543;
   reg _397544_397544 ; 
   reg __397544_397544;
   reg _397545_397545 ; 
   reg __397545_397545;
   reg _397546_397546 ; 
   reg __397546_397546;
   reg _397547_397547 ; 
   reg __397547_397547;
   reg _397548_397548 ; 
   reg __397548_397548;
   reg _397549_397549 ; 
   reg __397549_397549;
   reg _397550_397550 ; 
   reg __397550_397550;
   reg _397551_397551 ; 
   reg __397551_397551;
   reg _397552_397552 ; 
   reg __397552_397552;
   reg _397553_397553 ; 
   reg __397553_397553;
   reg _397554_397554 ; 
   reg __397554_397554;
   reg _397555_397555 ; 
   reg __397555_397555;
   reg _397556_397556 ; 
   reg __397556_397556;
   reg _397557_397557 ; 
   reg __397557_397557;
   reg _397558_397558 ; 
   reg __397558_397558;
   reg _397559_397559 ; 
   reg __397559_397559;
   reg _397560_397560 ; 
   reg __397560_397560;
   reg _397561_397561 ; 
   reg __397561_397561;
   reg _397562_397562 ; 
   reg __397562_397562;
   reg _397563_397563 ; 
   reg __397563_397563;
   reg _397564_397564 ; 
   reg __397564_397564;
   reg _397565_397565 ; 
   reg __397565_397565;
   reg _397566_397566 ; 
   reg __397566_397566;
   reg _397567_397567 ; 
   reg __397567_397567;
   reg _397568_397568 ; 
   reg __397568_397568;
   reg _397569_397569 ; 
   reg __397569_397569;
   reg _397570_397570 ; 
   reg __397570_397570;
   reg _397571_397571 ; 
   reg __397571_397571;
   reg _397572_397572 ; 
   reg __397572_397572;
   reg _397573_397573 ; 
   reg __397573_397573;
   reg _397574_397574 ; 
   reg __397574_397574;
   reg _397575_397575 ; 
   reg __397575_397575;
   reg _397576_397576 ; 
   reg __397576_397576;
   reg _397577_397577 ; 
   reg __397577_397577;
   reg _397578_397578 ; 
   reg __397578_397578;
   reg _397579_397579 ; 
   reg __397579_397579;
   reg _397580_397580 ; 
   reg __397580_397580;
   reg _397581_397581 ; 
   reg __397581_397581;
   reg _397582_397582 ; 
   reg __397582_397582;
   reg _397583_397583 ; 
   reg __397583_397583;
   reg _397584_397584 ; 
   reg __397584_397584;
   reg _397585_397585 ; 
   reg __397585_397585;
   reg _397586_397586 ; 
   reg __397586_397586;
   reg _397587_397587 ; 
   reg __397587_397587;
   reg _397588_397588 ; 
   reg __397588_397588;
   reg _397589_397589 ; 
   reg __397589_397589;
   reg _397590_397590 ; 
   reg __397590_397590;
   reg _397591_397591 ; 
   reg __397591_397591;
   reg _397592_397592 ; 
   reg __397592_397592;
   reg _397593_397593 ; 
   reg __397593_397593;
   reg _397594_397594 ; 
   reg __397594_397594;
   reg _397595_397595 ; 
   reg __397595_397595;
   reg _397596_397596 ; 
   reg __397596_397596;
   reg _397597_397597 ; 
   reg __397597_397597;
   reg _397598_397598 ; 
   reg __397598_397598;
   reg _397599_397599 ; 
   reg __397599_397599;
   reg _397600_397600 ; 
   reg __397600_397600;
   reg _397601_397601 ; 
   reg __397601_397601;
   reg _397602_397602 ; 
   reg __397602_397602;
   reg _397603_397603 ; 
   reg __397603_397603;
   reg _397604_397604 ; 
   reg __397604_397604;
   reg _397605_397605 ; 
   reg __397605_397605;
   reg _397606_397606 ; 
   reg __397606_397606;
   reg _397607_397607 ; 
   reg __397607_397607;
   reg _397608_397608 ; 
   reg __397608_397608;
   reg _397609_397609 ; 
   reg __397609_397609;
   reg _397610_397610 ; 
   reg __397610_397610;
   reg _397611_397611 ; 
   reg __397611_397611;
   reg _397612_397612 ; 
   reg __397612_397612;
   reg _397613_397613 ; 
   reg __397613_397613;
   reg _397614_397614 ; 
   reg __397614_397614;
   reg _397615_397615 ; 
   reg __397615_397615;
   reg _397616_397616 ; 
   reg __397616_397616;
   reg _397617_397617 ; 
   reg __397617_397617;
   reg _397618_397618 ; 
   reg __397618_397618;
   reg _397619_397619 ; 
   reg __397619_397619;
   reg _397620_397620 ; 
   reg __397620_397620;
   reg _397621_397621 ; 
   reg __397621_397621;
   reg _397622_397622 ; 
   reg __397622_397622;
   reg _397623_397623 ; 
   reg __397623_397623;
   reg _397624_397624 ; 
   reg __397624_397624;
   reg _397625_397625 ; 
   reg __397625_397625;
   reg _397626_397626 ; 
   reg __397626_397626;
   reg _397627_397627 ; 
   reg __397627_397627;
   reg _397628_397628 ; 
   reg __397628_397628;
   reg _397629_397629 ; 
   reg __397629_397629;
   reg _397630_397630 ; 
   reg __397630_397630;
   reg _397631_397631 ; 
   reg __397631_397631;
   reg _397632_397632 ; 
   reg __397632_397632;
   reg _397633_397633 ; 
   reg __397633_397633;
   reg _397634_397634 ; 
   reg __397634_397634;
   reg _397635_397635 ; 
   reg __397635_397635;
   reg _397636_397636 ; 
   reg __397636_397636;
   reg _397637_397637 ; 
   reg __397637_397637;
   reg _397638_397638 ; 
   reg __397638_397638;
   reg _397639_397639 ; 
   reg __397639_397639;
   reg _397640_397640 ; 
   reg __397640_397640;
   reg _397641_397641 ; 
   reg __397641_397641;
   reg _397642_397642 ; 
   reg __397642_397642;
   reg _397643_397643 ; 
   reg __397643_397643;
   reg _397644_397644 ; 
   reg __397644_397644;
   reg _397645_397645 ; 
   reg __397645_397645;
   reg _397646_397646 ; 
   reg __397646_397646;
   reg _397647_397647 ; 
   reg __397647_397647;
   reg _397648_397648 ; 
   reg __397648_397648;
   reg _397649_397649 ; 
   reg __397649_397649;
   reg _397650_397650 ; 
   reg __397650_397650;
   reg _397651_397651 ; 
   reg __397651_397651;
   reg _397652_397652 ; 
   reg __397652_397652;
   reg _397653_397653 ; 
   reg __397653_397653;
   reg _397654_397654 ; 
   reg __397654_397654;
   reg _397655_397655 ; 
   reg __397655_397655;
   reg _397656_397656 ; 
   reg __397656_397656;
   reg _397657_397657 ; 
   reg __397657_397657;
   reg _397658_397658 ; 
   reg __397658_397658;
   reg _397659_397659 ; 
   reg __397659_397659;
   reg _397660_397660 ; 
   reg __397660_397660;
   reg _397661_397661 ; 
   reg __397661_397661;
   reg _397662_397662 ; 
   reg __397662_397662;
   reg _397663_397663 ; 
   reg __397663_397663;
   reg _397664_397664 ; 
   reg __397664_397664;
   reg _397665_397665 ; 
   reg __397665_397665;
   reg _397666_397666 ; 
   reg __397666_397666;
   reg _397667_397667 ; 
   reg __397667_397667;
   reg _397668_397668 ; 
   reg __397668_397668;
   reg _397669_397669 ; 
   reg __397669_397669;
   reg _397670_397670 ; 
   reg __397670_397670;
   reg _397671_397671 ; 
   reg __397671_397671;
   reg _397672_397672 ; 
   reg __397672_397672;
   reg _397673_397673 ; 
   reg __397673_397673;
   reg _397674_397674 ; 
   reg __397674_397674;
   reg _397675_397675 ; 
   reg __397675_397675;
   reg _397676_397676 ; 
   reg __397676_397676;
   reg _397677_397677 ; 
   reg __397677_397677;
   reg _397678_397678 ; 
   reg __397678_397678;
   reg _397679_397679 ; 
   reg __397679_397679;
   reg _397680_397680 ; 
   reg __397680_397680;
   reg _397681_397681 ; 
   reg __397681_397681;
   reg _397682_397682 ; 
   reg __397682_397682;
   reg _397683_397683 ; 
   reg __397683_397683;
   reg _397684_397684 ; 
   reg __397684_397684;
   reg _397685_397685 ; 
   reg __397685_397685;
   reg _397686_397686 ; 
   reg __397686_397686;
   reg _397687_397687 ; 
   reg __397687_397687;
   reg _397688_397688 ; 
   reg __397688_397688;
   reg _397689_397689 ; 
   reg __397689_397689;
   reg _397690_397690 ; 
   reg __397690_397690;
   reg _397691_397691 ; 
   reg __397691_397691;
   reg _397692_397692 ; 
   reg __397692_397692;
   reg _397693_397693 ; 
   reg __397693_397693;
   reg _397694_397694 ; 
   reg __397694_397694;
   reg _397695_397695 ; 
   reg __397695_397695;
   reg _397696_397696 ; 
   reg __397696_397696;
   reg _397697_397697 ; 
   reg __397697_397697;
   reg _397698_397698 ; 
   reg __397698_397698;
   reg _397699_397699 ; 
   reg __397699_397699;
   reg _397700_397700 ; 
   reg __397700_397700;
   reg _397701_397701 ; 
   reg __397701_397701;
   reg _397702_397702 ; 
   reg __397702_397702;
   reg _397703_397703 ; 
   reg __397703_397703;
   reg _397704_397704 ; 
   reg __397704_397704;
   reg _397705_397705 ; 
   reg __397705_397705;
   reg _397706_397706 ; 
   reg __397706_397706;
   reg _397707_397707 ; 
   reg __397707_397707;
   reg _397708_397708 ; 
   reg __397708_397708;
   reg _397709_397709 ; 
   reg __397709_397709;
   reg _397710_397710 ; 
   reg __397710_397710;
   reg _397711_397711 ; 
   reg __397711_397711;
   reg _397712_397712 ; 
   reg __397712_397712;
   reg _397713_397713 ; 
   reg __397713_397713;
   reg _397714_397714 ; 
   reg __397714_397714;
   reg _397715_397715 ; 
   reg __397715_397715;
   reg _397716_397716 ; 
   reg __397716_397716;
   reg _397717_397717 ; 
   reg __397717_397717;
   reg _397718_397718 ; 
   reg __397718_397718;
   reg _397719_397719 ; 
   reg __397719_397719;
   reg _397720_397720 ; 
   reg __397720_397720;
   reg _397721_397721 ; 
   reg __397721_397721;
   reg _397722_397722 ; 
   reg __397722_397722;
   reg _397723_397723 ; 
   reg __397723_397723;
   reg _397724_397724 ; 
   reg __397724_397724;
   reg _397725_397725 ; 
   reg __397725_397725;
   reg _397726_397726 ; 
   reg __397726_397726;
   reg _397727_397727 ; 
   reg __397727_397727;
   reg _397728_397728 ; 
   reg __397728_397728;
   reg _397729_397729 ; 
   reg __397729_397729;
   reg _397730_397730 ; 
   reg __397730_397730;
   reg _397731_397731 ; 
   reg __397731_397731;
   reg _397732_397732 ; 
   reg __397732_397732;
   reg _397733_397733 ; 
   reg __397733_397733;
   reg _397734_397734 ; 
   reg __397734_397734;
   reg _397735_397735 ; 
   reg __397735_397735;
   reg _397736_397736 ; 
   reg __397736_397736;
   reg _397737_397737 ; 
   reg __397737_397737;
   reg _397738_397738 ; 
   reg __397738_397738;
   reg _397739_397739 ; 
   reg __397739_397739;
   reg _397740_397740 ; 
   reg __397740_397740;
   reg _397741_397741 ; 
   reg __397741_397741;
   reg _397742_397742 ; 
   reg __397742_397742;
   reg _397743_397743 ; 
   reg __397743_397743;
   reg _397744_397744 ; 
   reg __397744_397744;
   reg _397745_397745 ; 
   reg __397745_397745;
   reg _397746_397746 ; 
   reg __397746_397746;
   reg _397747_397747 ; 
   reg __397747_397747;
   reg _397748_397748 ; 
   reg __397748_397748;
   reg _397749_397749 ; 
   reg __397749_397749;
   reg _397750_397750 ; 
   reg __397750_397750;
   reg _397751_397751 ; 
   reg __397751_397751;
   reg _397752_397752 ; 
   reg __397752_397752;
   reg _397753_397753 ; 
   reg __397753_397753;
   reg _397754_397754 ; 
   reg __397754_397754;
   reg _397755_397755 ; 
   reg __397755_397755;
   reg _397756_397756 ; 
   reg __397756_397756;
   reg _397757_397757 ; 
   reg __397757_397757;
   reg _397758_397758 ; 
   reg __397758_397758;
   reg _397759_397759 ; 
   reg __397759_397759;
   reg _397760_397760 ; 
   reg __397760_397760;
   reg _397761_397761 ; 
   reg __397761_397761;
   reg _397762_397762 ; 
   reg __397762_397762;
   reg _397763_397763 ; 
   reg __397763_397763;
   reg _397764_397764 ; 
   reg __397764_397764;
   reg _397765_397765 ; 
   reg __397765_397765;
   reg _397766_397766 ; 
   reg __397766_397766;
   reg _397767_397767 ; 
   reg __397767_397767;
   reg _397768_397768 ; 
   reg __397768_397768;
   reg _397769_397769 ; 
   reg __397769_397769;
   reg _397770_397770 ; 
   reg __397770_397770;
   reg _397771_397771 ; 
   reg __397771_397771;
   reg _397772_397772 ; 
   reg __397772_397772;
   reg _397773_397773 ; 
   reg __397773_397773;
   reg _397774_397774 ; 
   reg __397774_397774;
   reg _397775_397775 ; 
   reg __397775_397775;
   reg _397776_397776 ; 
   reg __397776_397776;
   reg _397777_397777 ; 
   reg __397777_397777;
   reg _397778_397778 ; 
   reg __397778_397778;
   reg _397779_397779 ; 
   reg __397779_397779;
   reg _397780_397780 ; 
   reg __397780_397780;
   reg _397781_397781 ; 
   reg __397781_397781;
   reg _397782_397782 ; 
   reg __397782_397782;
   reg _397783_397783 ; 
   reg __397783_397783;
   reg _397784_397784 ; 
   reg __397784_397784;
   reg _397785_397785 ; 
   reg __397785_397785;
   reg _397786_397786 ; 
   reg __397786_397786;
   reg _397787_397787 ; 
   reg __397787_397787;
   reg _397788_397788 ; 
   reg __397788_397788;
   reg _397789_397789 ; 
   reg __397789_397789;
   reg _397790_397790 ; 
   reg __397790_397790;
   reg _397791_397791 ; 
   reg __397791_397791;
   reg _397792_397792 ; 
   reg __397792_397792;
   reg _397793_397793 ; 
   reg __397793_397793;
   reg _397794_397794 ; 
   reg __397794_397794;
   reg _397795_397795 ; 
   reg __397795_397795;
   reg _397796_397796 ; 
   reg __397796_397796;
   reg _397797_397797 ; 
   reg __397797_397797;
   reg _397798_397798 ; 
   reg __397798_397798;
   reg _397799_397799 ; 
   reg __397799_397799;
   reg _397800_397800 ; 
   reg __397800_397800;
   reg _397801_397801 ; 
   reg __397801_397801;
   reg _397802_397802 ; 
   reg __397802_397802;
   reg _397803_397803 ; 
   reg __397803_397803;
   reg _397804_397804 ; 
   reg __397804_397804;
   reg _397805_397805 ; 
   reg __397805_397805;
   reg _397806_397806 ; 
   reg __397806_397806;
   reg _397807_397807 ; 
   reg __397807_397807;
   reg _397808_397808 ; 
   reg __397808_397808;
   reg _397809_397809 ; 
   reg __397809_397809;
   reg _397810_397810 ; 
   reg __397810_397810;
   reg _397811_397811 ; 
   reg __397811_397811;
   reg _397812_397812 ; 
   reg __397812_397812;
   reg _397813_397813 ; 
   reg __397813_397813;
   reg _397814_397814 ; 
   reg __397814_397814;
   reg _397815_397815 ; 
   reg __397815_397815;
   reg _397816_397816 ; 
   reg __397816_397816;
   reg _397817_397817 ; 
   reg __397817_397817;
   reg _397818_397818 ; 
   reg __397818_397818;
   reg _397819_397819 ; 
   reg __397819_397819;
   reg _397820_397820 ; 
   reg __397820_397820;
   reg _397821_397821 ; 
   reg __397821_397821;
   reg _397822_397822 ; 
   reg __397822_397822;
   reg _397823_397823 ; 
   reg __397823_397823;
   reg _397824_397824 ; 
   reg __397824_397824;
   reg _397825_397825 ; 
   reg __397825_397825;
   reg _397826_397826 ; 
   reg __397826_397826;
   reg _397827_397827 ; 
   reg __397827_397827;
   reg _397828_397828 ; 
   reg __397828_397828;
   reg _397829_397829 ; 
   reg __397829_397829;
   reg _397830_397830 ; 
   reg __397830_397830;
   reg _397831_397831 ; 
   reg __397831_397831;
   reg _397832_397832 ; 
   reg __397832_397832;
   reg _397833_397833 ; 
   reg __397833_397833;
   reg _397834_397834 ; 
   reg __397834_397834;
   reg _397835_397835 ; 
   reg __397835_397835;
   reg _397836_397836 ; 
   reg __397836_397836;
   reg _397837_397837 ; 
   reg __397837_397837;
   reg _397838_397838 ; 
   reg __397838_397838;
   reg _397839_397839 ; 
   reg __397839_397839;
   reg _397840_397840 ; 
   reg __397840_397840;
   reg _397841_397841 ; 
   reg __397841_397841;
   reg _397842_397842 ; 
   reg __397842_397842;
   reg _397843_397843 ; 
   reg __397843_397843;
   reg _397844_397844 ; 
   reg __397844_397844;
   reg _397845_397845 ; 
   reg __397845_397845;
   reg _397846_397846 ; 
   reg __397846_397846;
   reg _397847_397847 ; 
   reg __397847_397847;
   reg _397848_397848 ; 
   reg __397848_397848;
   reg _397849_397849 ; 
   reg __397849_397849;
   reg _397850_397850 ; 
   reg __397850_397850;
   reg _397851_397851 ; 
   reg __397851_397851;
   reg _397852_397852 ; 
   reg __397852_397852;
   reg _397853_397853 ; 
   reg __397853_397853;
   reg _397854_397854 ; 
   reg __397854_397854;
   reg _397855_397855 ; 
   reg __397855_397855;
   reg _397856_397856 ; 
   reg __397856_397856;
   reg _397857_397857 ; 
   reg __397857_397857;
   reg _397858_397858 ; 
   reg __397858_397858;
   reg _397859_397859 ; 
   reg __397859_397859;
   reg _397860_397860 ; 
   reg __397860_397860;
   reg _397861_397861 ; 
   reg __397861_397861;
   reg _397862_397862 ; 
   reg __397862_397862;
   reg _397863_397863 ; 
   reg __397863_397863;
   reg _397864_397864 ; 
   reg __397864_397864;
   reg _397865_397865 ; 
   reg __397865_397865;
   reg _397866_397866 ; 
   reg __397866_397866;
   reg _397867_397867 ; 
   reg __397867_397867;
   reg _397868_397868 ; 
   reg __397868_397868;
   reg _397869_397869 ; 
   reg __397869_397869;
   reg _397870_397870 ; 
   reg __397870_397870;
   reg _397871_397871 ; 
   reg __397871_397871;
   reg _397872_397872 ; 
   reg __397872_397872;
   reg _397873_397873 ; 
   reg __397873_397873;
   reg _397874_397874 ; 
   reg __397874_397874;
   reg _397875_397875 ; 
   reg __397875_397875;
   reg _397876_397876 ; 
   reg __397876_397876;
   reg _397877_397877 ; 
   reg __397877_397877;
   reg _397878_397878 ; 
   reg __397878_397878;
   reg _397879_397879 ; 
   reg __397879_397879;
   reg _397880_397880 ; 
   reg __397880_397880;
   reg _397881_397881 ; 
   reg __397881_397881;
   reg _397882_397882 ; 
   reg __397882_397882;
   reg _397883_397883 ; 
   reg __397883_397883;
   reg _397884_397884 ; 
   reg __397884_397884;
   reg _397885_397885 ; 
   reg __397885_397885;
   reg _397886_397886 ; 
   reg __397886_397886;
   reg _397887_397887 ; 
   reg __397887_397887;
   reg _397888_397888 ; 
   reg __397888_397888;
   reg _397889_397889 ; 
   reg __397889_397889;
   reg _397890_397890 ; 
   reg __397890_397890;
   reg _397891_397891 ; 
   reg __397891_397891;
   reg _397892_397892 ; 
   reg __397892_397892;
   reg _397893_397893 ; 
   reg __397893_397893;
   reg _397894_397894 ; 
   reg __397894_397894;
   reg _397895_397895 ; 
   reg __397895_397895;
   reg _397896_397896 ; 
   reg __397896_397896;
   reg _397897_397897 ; 
   reg __397897_397897;
   reg _397898_397898 ; 
   reg __397898_397898;
   reg _397899_397899 ; 
   reg __397899_397899;
   reg _397900_397900 ; 
   reg __397900_397900;
   reg _397901_397901 ; 
   reg __397901_397901;
   reg _397902_397902 ; 
   reg __397902_397902;
   reg _397903_397903 ; 
   reg __397903_397903;
   reg _397904_397904 ; 
   reg __397904_397904;
   reg _397905_397905 ; 
   reg __397905_397905;
   reg _397906_397906 ; 
   reg __397906_397906;
   reg _397907_397907 ; 
   reg __397907_397907;
   reg _397908_397908 ; 
   reg __397908_397908;
   reg _397909_397909 ; 
   reg __397909_397909;
   reg _397910_397910 ; 
   reg __397910_397910;
   reg _397911_397911 ; 
   reg __397911_397911;
   reg _397912_397912 ; 
   reg __397912_397912;
   reg _397913_397913 ; 
   reg __397913_397913;
   reg _397914_397914 ; 
   reg __397914_397914;
   reg _397915_397915 ; 
   reg __397915_397915;
   reg _397916_397916 ; 
   reg __397916_397916;
   reg _397917_397917 ; 
   reg __397917_397917;
   reg _397918_397918 ; 
   reg __397918_397918;
   reg _397919_397919 ; 
   reg __397919_397919;
   reg _397920_397920 ; 
   reg __397920_397920;
   reg _397921_397921 ; 
   reg __397921_397921;
   reg _397922_397922 ; 
   reg __397922_397922;
   reg _397923_397923 ; 
   reg __397923_397923;
   reg _397924_397924 ; 
   reg __397924_397924;
   reg _397925_397925 ; 
   reg __397925_397925;
   reg _397926_397926 ; 
   reg __397926_397926;
   reg _397927_397927 ; 
   reg __397927_397927;
   reg _397928_397928 ; 
   reg __397928_397928;
   reg _397929_397929 ; 
   reg __397929_397929;
   reg _397930_397930 ; 
   reg __397930_397930;
   reg _397931_397931 ; 
   reg __397931_397931;
   reg _397932_397932 ; 
   reg __397932_397932;
   reg _397933_397933 ; 
   reg __397933_397933;
   reg _397934_397934 ; 
   reg __397934_397934;
   reg _397935_397935 ; 
   reg __397935_397935;
   reg _397936_397936 ; 
   reg __397936_397936;
   reg _397937_397937 ; 
   reg __397937_397937;
   reg _397938_397938 ; 
   reg __397938_397938;
   reg _397939_397939 ; 
   reg __397939_397939;
   reg _397940_397940 ; 
   reg __397940_397940;
   reg _397941_397941 ; 
   reg __397941_397941;
   reg _397942_397942 ; 
   reg __397942_397942;
   reg _397943_397943 ; 
   reg __397943_397943;
   reg _397944_397944 ; 
   reg __397944_397944;
   reg _397945_397945 ; 
   reg __397945_397945;
   reg _397946_397946 ; 
   reg __397946_397946;
   reg _397947_397947 ; 
   reg __397947_397947;
   reg _397948_397948 ; 
   reg __397948_397948;
   reg _397949_397949 ; 
   reg __397949_397949;
   reg _397950_397950 ; 
   reg __397950_397950;
   reg _397951_397951 ; 
   reg __397951_397951;
   reg _397952_397952 ; 
   reg __397952_397952;
   reg _397953_397953 ; 
   reg __397953_397953;
   reg _397954_397954 ; 
   reg __397954_397954;
   reg _397955_397955 ; 
   reg __397955_397955;
   reg _397956_397956 ; 
   reg __397956_397956;
   reg _397957_397957 ; 
   reg __397957_397957;
   reg _397958_397958 ; 
   reg __397958_397958;
   reg _397959_397959 ; 
   reg __397959_397959;
   reg _397960_397960 ; 
   reg __397960_397960;
   reg _397961_397961 ; 
   reg __397961_397961;
   reg _397962_397962 ; 
   reg __397962_397962;
   reg _397963_397963 ; 
   reg __397963_397963;
   reg _397964_397964 ; 
   reg __397964_397964;
   reg _397965_397965 ; 
   reg __397965_397965;
   reg _397966_397966 ; 
   reg __397966_397966;
   reg _397967_397967 ; 
   reg __397967_397967;
   reg _397968_397968 ; 
   reg __397968_397968;
   reg _397969_397969 ; 
   reg __397969_397969;
   reg _397970_397970 ; 
   reg __397970_397970;
   reg _397971_397971 ; 
   reg __397971_397971;
   reg _397972_397972 ; 
   reg __397972_397972;
   reg _397973_397973 ; 
   reg __397973_397973;
   reg _397974_397974 ; 
   reg __397974_397974;
   reg _397975_397975 ; 
   reg __397975_397975;
   reg _397976_397976 ; 
   reg __397976_397976;
   reg _397977_397977 ; 
   reg __397977_397977;
   reg _397978_397978 ; 
   reg __397978_397978;
   reg _397979_397979 ; 
   reg __397979_397979;
   reg _397980_397980 ; 
   reg __397980_397980;
   reg _397981_397981 ; 
   reg __397981_397981;
   reg _397982_397982 ; 
   reg __397982_397982;
   reg _397983_397983 ; 
   reg __397983_397983;
   reg _397984_397984 ; 
   reg __397984_397984;
   reg _397985_397985 ; 
   reg __397985_397985;
   reg _397986_397986 ; 
   reg __397986_397986;
   reg _397987_397987 ; 
   reg __397987_397987;
   reg _397988_397988 ; 
   reg __397988_397988;
   reg _397989_397989 ; 
   reg __397989_397989;
   reg _397990_397990 ; 
   reg __397990_397990;
   reg _397991_397991 ; 
   reg __397991_397991;
   reg _397992_397992 ; 
   reg __397992_397992;
   reg _397993_397993 ; 
   reg __397993_397993;
   reg _397994_397994 ; 
   reg __397994_397994;
   reg _397995_397995 ; 
   reg __397995_397995;
   reg _397996_397996 ; 
   reg __397996_397996;
   reg _397997_397997 ; 
   reg __397997_397997;
   reg _397998_397998 ; 
   reg __397998_397998;
   reg _397999_397999 ; 
   reg __397999_397999;
   reg _398000_398000 ; 
   reg __398000_398000;
   reg _398001_398001 ; 
   reg __398001_398001;
   reg _398002_398002 ; 
   reg __398002_398002;
   reg _398003_398003 ; 
   reg __398003_398003;
   reg _398004_398004 ; 
   reg __398004_398004;
   reg _398005_398005 ; 
   reg __398005_398005;
   reg _398006_398006 ; 
   reg __398006_398006;
   reg _398007_398007 ; 
   reg __398007_398007;
   reg _398008_398008 ; 
   reg __398008_398008;
   reg _398009_398009 ; 
   reg __398009_398009;
   reg _398010_398010 ; 
   reg __398010_398010;
   reg _398011_398011 ; 
   reg __398011_398011;
   reg _398012_398012 ; 
   reg __398012_398012;
   reg _398013_398013 ; 
   reg __398013_398013;
   reg _398014_398014 ; 
   reg __398014_398014;
   reg _398015_398015 ; 
   reg __398015_398015;
   reg _398016_398016 ; 
   reg __398016_398016;
   reg _398017_398017 ; 
   reg __398017_398017;
   reg _398018_398018 ; 
   reg __398018_398018;
   reg _398019_398019 ; 
   reg __398019_398019;
   reg _398020_398020 ; 
   reg __398020_398020;
   reg _398021_398021 ; 
   reg __398021_398021;
   reg _398022_398022 ; 
   reg __398022_398022;
   reg _398023_398023 ; 
   reg __398023_398023;
   reg _398024_398024 ; 
   reg __398024_398024;
   reg _398025_398025 ; 
   reg __398025_398025;
   reg _398026_398026 ; 
   reg __398026_398026;
   reg _398027_398027 ; 
   reg __398027_398027;
   reg _398028_398028 ; 
   reg __398028_398028;
   reg _398029_398029 ; 
   reg __398029_398029;
   reg _398030_398030 ; 
   reg __398030_398030;
   reg _398031_398031 ; 
   reg __398031_398031;
   reg _398032_398032 ; 
   reg __398032_398032;
   reg _398033_398033 ; 
   reg __398033_398033;
   reg _398034_398034 ; 
   reg __398034_398034;
   reg _398035_398035 ; 
   reg __398035_398035;
   reg _398036_398036 ; 
   reg __398036_398036;
   reg _398037_398037 ; 
   reg __398037_398037;
   reg _398038_398038 ; 
   reg __398038_398038;
   reg _398039_398039 ; 
   reg __398039_398039;
   reg _398040_398040 ; 
   reg __398040_398040;
   reg _398041_398041 ; 
   reg __398041_398041;
   reg _398042_398042 ; 
   reg __398042_398042;
   reg _398043_398043 ; 
   reg __398043_398043;
   reg _398044_398044 ; 
   reg __398044_398044;
   reg _398045_398045 ; 
   reg __398045_398045;
   reg _398046_398046 ; 
   reg __398046_398046;
   reg _398047_398047 ; 
   reg __398047_398047;
   reg _398048_398048 ; 
   reg __398048_398048;
   reg _398049_398049 ; 
   reg __398049_398049;
   reg _398050_398050 ; 
   reg __398050_398050;
   reg _398051_398051 ; 
   reg __398051_398051;
   reg _398052_398052 ; 
   reg __398052_398052;
   reg _398053_398053 ; 
   reg __398053_398053;
   reg _398054_398054 ; 
   reg __398054_398054;
   reg _398055_398055 ; 
   reg __398055_398055;
   reg _398056_398056 ; 
   reg __398056_398056;
   reg _398057_398057 ; 
   reg __398057_398057;
   reg _398058_398058 ; 
   reg __398058_398058;
   reg _398059_398059 ; 
   reg __398059_398059;
   reg _398060_398060 ; 
   reg __398060_398060;
   reg _398061_398061 ; 
   reg __398061_398061;
   reg _398062_398062 ; 
   reg __398062_398062;
   reg _398063_398063 ; 
   reg __398063_398063;
   reg _398064_398064 ; 
   reg __398064_398064;
   reg _398065_398065 ; 
   reg __398065_398065;
   reg _398066_398066 ; 
   reg __398066_398066;
   reg _398067_398067 ; 
   reg __398067_398067;
   reg _398068_398068 ; 
   reg __398068_398068;
   reg _398069_398069 ; 
   reg __398069_398069;
   reg _398070_398070 ; 
   reg __398070_398070;
   reg _398071_398071 ; 
   reg __398071_398071;
   reg _398072_398072 ; 
   reg __398072_398072;
   reg _398073_398073 ; 
   reg __398073_398073;
   reg _398074_398074 ; 
   reg __398074_398074;
   reg _398075_398075 ; 
   reg __398075_398075;
   reg _398076_398076 ; 
   reg __398076_398076;
   reg _398077_398077 ; 
   reg __398077_398077;
   reg _398078_398078 ; 
   reg __398078_398078;
   reg _398079_398079 ; 
   reg __398079_398079;
   reg _398080_398080 ; 
   reg __398080_398080;
   reg _398081_398081 ; 
   reg __398081_398081;
   reg _398082_398082 ; 
   reg __398082_398082;
   reg _398083_398083 ; 
   reg __398083_398083;
   reg _398084_398084 ; 
   reg __398084_398084;
   reg _398085_398085 ; 
   reg __398085_398085;
   reg _398086_398086 ; 
   reg __398086_398086;
   reg _398087_398087 ; 
   reg __398087_398087;
   reg _398088_398088 ; 
   reg __398088_398088;
   reg _398089_398089 ; 
   reg __398089_398089;
   reg _398090_398090 ; 
   reg __398090_398090;
   reg _398091_398091 ; 
   reg __398091_398091;
   reg _398092_398092 ; 
   reg __398092_398092;
   reg _398093_398093 ; 
   reg __398093_398093;
   reg _398094_398094 ; 
   reg __398094_398094;
   reg _398095_398095 ; 
   reg __398095_398095;
   reg _398096_398096 ; 
   reg __398096_398096;
   reg _398097_398097 ; 
   reg __398097_398097;
   reg _398098_398098 ; 
   reg __398098_398098;
   reg _398099_398099 ; 
   reg __398099_398099;
   reg _398100_398100 ; 
   reg __398100_398100;
   reg _398101_398101 ; 
   reg __398101_398101;
   reg _398102_398102 ; 
   reg __398102_398102;
   reg _398103_398103 ; 
   reg __398103_398103;
   reg _398104_398104 ; 
   reg __398104_398104;
   reg _398105_398105 ; 
   reg __398105_398105;
   reg _398106_398106 ; 
   reg __398106_398106;
   reg _398107_398107 ; 
   reg __398107_398107;
   reg _398108_398108 ; 
   reg __398108_398108;
   reg _398109_398109 ; 
   reg __398109_398109;
   reg _398110_398110 ; 
   reg __398110_398110;
   reg _398111_398111 ; 
   reg __398111_398111;
   reg _398112_398112 ; 
   reg __398112_398112;
   reg _398113_398113 ; 
   reg __398113_398113;
   reg _398114_398114 ; 
   reg __398114_398114;
   reg _398115_398115 ; 
   reg __398115_398115;
   reg _398116_398116 ; 
   reg __398116_398116;
   reg _398117_398117 ; 
   reg __398117_398117;
   reg _398118_398118 ; 
   reg __398118_398118;
   reg _398119_398119 ; 
   reg __398119_398119;
   reg _398120_398120 ; 
   reg __398120_398120;
   reg _398121_398121 ; 
   reg __398121_398121;
   reg _398122_398122 ; 
   reg __398122_398122;
   reg _398123_398123 ; 
   reg __398123_398123;
   reg _398124_398124 ; 
   reg __398124_398124;
   reg _398125_398125 ; 
   reg __398125_398125;
   reg _398126_398126 ; 
   reg __398126_398126;
   reg _398127_398127 ; 
   reg __398127_398127;
   reg _398128_398128 ; 
   reg __398128_398128;
   reg _398129_398129 ; 
   reg __398129_398129;
   reg _398130_398130 ; 
   reg __398130_398130;
   reg _398131_398131 ; 
   reg __398131_398131;
   reg _398132_398132 ; 
   reg __398132_398132;
   reg _398133_398133 ; 
   reg __398133_398133;
   reg _398134_398134 ; 
   reg __398134_398134;
   reg _398135_398135 ; 
   reg __398135_398135;
   reg _398136_398136 ; 
   reg __398136_398136;
   reg _398137_398137 ; 
   reg __398137_398137;
   reg _398138_398138 ; 
   reg __398138_398138;
   reg _398139_398139 ; 
   reg __398139_398139;
   reg _398140_398140 ; 
   reg __398140_398140;
   reg _398141_398141 ; 
   reg __398141_398141;
   reg _398142_398142 ; 
   reg __398142_398142;
   reg _398143_398143 ; 
   reg __398143_398143;
   reg _398144_398144 ; 
   reg __398144_398144;
   reg _398145_398145 ; 
   reg __398145_398145;
   reg _398146_398146 ; 
   reg __398146_398146;
   reg _398147_398147 ; 
   reg __398147_398147;
   reg _398148_398148 ; 
   reg __398148_398148;
   reg _398149_398149 ; 
   reg __398149_398149;
   reg _398150_398150 ; 
   reg __398150_398150;
   reg _398151_398151 ; 
   reg __398151_398151;
   reg _398152_398152 ; 
   reg __398152_398152;
   reg _398153_398153 ; 
   reg __398153_398153;
   reg _398154_398154 ; 
   reg __398154_398154;
   reg _398155_398155 ; 
   reg __398155_398155;
   reg _398156_398156 ; 
   reg __398156_398156;
   reg _398157_398157 ; 
   reg __398157_398157;
   reg _398158_398158 ; 
   reg __398158_398158;
   reg _398159_398159 ; 
   reg __398159_398159;
   reg _398160_398160 ; 
   reg __398160_398160;
   reg _398161_398161 ; 
   reg __398161_398161;
   reg _398162_398162 ; 
   reg __398162_398162;
   reg _398163_398163 ; 
   reg __398163_398163;
   reg _398164_398164 ; 
   reg __398164_398164;
   reg _398165_398165 ; 
   reg __398165_398165;
   reg _398166_398166 ; 
   reg __398166_398166;
   reg _398167_398167 ; 
   reg __398167_398167;
   reg _398168_398168 ; 
   reg __398168_398168;
   reg _398169_398169 ; 
   reg __398169_398169;
   reg _398170_398170 ; 
   reg __398170_398170;
   reg _398171_398171 ; 
   reg __398171_398171;
   reg _398172_398172 ; 
   reg __398172_398172;
   reg _398173_398173 ; 
   reg __398173_398173;
   reg _398174_398174 ; 
   reg __398174_398174;
   reg _398175_398175 ; 
   reg __398175_398175;
   reg _398176_398176 ; 
   reg __398176_398176;
   reg _398177_398177 ; 
   reg __398177_398177;
   reg _398178_398178 ; 
   reg __398178_398178;
   reg _398179_398179 ; 
   reg __398179_398179;
   reg _398180_398180 ; 
   reg __398180_398180;
   reg _398181_398181 ; 
   reg __398181_398181;
   reg _398182_398182 ; 
   reg __398182_398182;
   reg _398183_398183 ; 
   reg __398183_398183;
   reg _398184_398184 ; 
   reg __398184_398184;
   reg _398185_398185 ; 
   reg __398185_398185;
   reg _398186_398186 ; 
   reg __398186_398186;
   reg _398187_398187 ; 
   reg __398187_398187;
   reg _398188_398188 ; 
   reg __398188_398188;
   reg _398189_398189 ; 
   reg __398189_398189;
   reg _398190_398190 ; 
   reg __398190_398190;
   reg _398191_398191 ; 
   reg __398191_398191;
   reg _398192_398192 ; 
   reg __398192_398192;
   reg _398193_398193 ; 
   reg __398193_398193;
   reg _398194_398194 ; 
   reg __398194_398194;
   reg _398195_398195 ; 
   reg __398195_398195;
   reg _398196_398196 ; 
   reg __398196_398196;
   reg _398197_398197 ; 
   reg __398197_398197;
   reg _398198_398198 ; 
   reg __398198_398198;
   reg _398199_398199 ; 
   reg __398199_398199;
   reg _398200_398200 ; 
   reg __398200_398200;
   reg _398201_398201 ; 
   reg __398201_398201;
   reg _398202_398202 ; 
   reg __398202_398202;
   reg _398203_398203 ; 
   reg __398203_398203;
   reg _398204_398204 ; 
   reg __398204_398204;
   reg _398205_398205 ; 
   reg __398205_398205;
   reg _398206_398206 ; 
   reg __398206_398206;
   reg _398207_398207 ; 
   reg __398207_398207;
   reg _398208_398208 ; 
   reg __398208_398208;
   reg _398209_398209 ; 
   reg __398209_398209;
   reg _398210_398210 ; 
   reg __398210_398210;
   reg _398211_398211 ; 
   reg __398211_398211;
   reg _398212_398212 ; 
   reg __398212_398212;
   reg _398213_398213 ; 
   reg __398213_398213;
   reg _398214_398214 ; 
   reg __398214_398214;
   reg _398215_398215 ; 
   reg __398215_398215;
   reg _398216_398216 ; 
   reg __398216_398216;
   reg _398217_398217 ; 
   reg __398217_398217;
   reg _398218_398218 ; 
   reg __398218_398218;
   reg _398219_398219 ; 
   reg __398219_398219;
   reg _398220_398220 ; 
   reg __398220_398220;
   reg _398221_398221 ; 
   reg __398221_398221;
   reg _398222_398222 ; 
   reg __398222_398222;
   reg _398223_398223 ; 
   reg __398223_398223;
   reg _398224_398224 ; 
   reg __398224_398224;
   reg _398225_398225 ; 
   reg __398225_398225;
   reg _398226_398226 ; 
   reg __398226_398226;
   reg _398227_398227 ; 
   reg __398227_398227;
   reg _398228_398228 ; 
   reg __398228_398228;
   reg _398229_398229 ; 
   reg __398229_398229;
   reg _398230_398230 ; 
   reg __398230_398230;
   reg _398231_398231 ; 
   reg __398231_398231;
   reg _398232_398232 ; 
   reg __398232_398232;
   reg _398233_398233 ; 
   reg __398233_398233;
   reg _398234_398234 ; 
   reg __398234_398234;
   reg _398235_398235 ; 
   reg __398235_398235;
   reg _398236_398236 ; 
   reg __398236_398236;
   reg _398237_398237 ; 
   reg __398237_398237;
   reg _398238_398238 ; 
   reg __398238_398238;
   reg _398239_398239 ; 
   reg __398239_398239;
   reg _398240_398240 ; 
   reg __398240_398240;
   reg _398241_398241 ; 
   reg __398241_398241;
   reg _398242_398242 ; 
   reg __398242_398242;
   reg _398243_398243 ; 
   reg __398243_398243;
   reg _398244_398244 ; 
   reg __398244_398244;
   reg _398245_398245 ; 
   reg __398245_398245;
   reg _398246_398246 ; 
   reg __398246_398246;
   reg _398247_398247 ; 
   reg __398247_398247;
   reg _398248_398248 ; 
   reg __398248_398248;
   reg _398249_398249 ; 
   reg __398249_398249;
   reg _398250_398250 ; 
   reg __398250_398250;
   reg _398251_398251 ; 
   reg __398251_398251;
   reg _398252_398252 ; 
   reg __398252_398252;
   reg _398253_398253 ; 
   reg __398253_398253;
   reg _398254_398254 ; 
   reg __398254_398254;
   reg _398255_398255 ; 
   reg __398255_398255;
   reg _398256_398256 ; 
   reg __398256_398256;
   reg _398257_398257 ; 
   reg __398257_398257;
   reg _398258_398258 ; 
   reg __398258_398258;
   reg _398259_398259 ; 
   reg __398259_398259;
   reg _398260_398260 ; 
   reg __398260_398260;
   reg _398261_398261 ; 
   reg __398261_398261;
   reg _398262_398262 ; 
   reg __398262_398262;
   reg _398263_398263 ; 
   reg __398263_398263;
   reg _398264_398264 ; 
   reg __398264_398264;
   reg _398265_398265 ; 
   reg __398265_398265;
   reg _398266_398266 ; 
   reg __398266_398266;
   reg _398267_398267 ; 
   reg __398267_398267;
   reg _398268_398268 ; 
   reg __398268_398268;
   reg _398269_398269 ; 
   reg __398269_398269;
   reg _398270_398270 ; 
   reg __398270_398270;
   reg _398271_398271 ; 
   reg __398271_398271;
   reg _398272_398272 ; 
   reg __398272_398272;
   reg _398273_398273 ; 
   reg __398273_398273;
   reg _398274_398274 ; 
   reg __398274_398274;
   reg _398275_398275 ; 
   reg __398275_398275;
   reg _398276_398276 ; 
   reg __398276_398276;
   reg _398277_398277 ; 
   reg __398277_398277;
   reg _398278_398278 ; 
   reg __398278_398278;
   reg _398279_398279 ; 
   reg __398279_398279;
   reg _398280_398280 ; 
   reg __398280_398280;
   reg _398281_398281 ; 
   reg __398281_398281;
   reg _398282_398282 ; 
   reg __398282_398282;
   reg _398283_398283 ; 
   reg __398283_398283;
   reg _398284_398284 ; 
   reg __398284_398284;
   reg _398285_398285 ; 
   reg __398285_398285;
   reg _398286_398286 ; 
   reg __398286_398286;
   reg _398287_398287 ; 
   reg __398287_398287;
   reg _398288_398288 ; 
   reg __398288_398288;
   reg _398289_398289 ; 
   reg __398289_398289;
   reg _398290_398290 ; 
   reg __398290_398290;
   reg _398291_398291 ; 
   reg __398291_398291;
   reg _398292_398292 ; 
   reg __398292_398292;
   reg _398293_398293 ; 
   reg __398293_398293;
   reg _398294_398294 ; 
   reg __398294_398294;
   reg _398295_398295 ; 
   reg __398295_398295;
   reg _398296_398296 ; 
   reg __398296_398296;
   reg _398297_398297 ; 
   reg __398297_398297;
   reg _398298_398298 ; 
   reg __398298_398298;
   reg _398299_398299 ; 
   reg __398299_398299;
   reg _398300_398300 ; 
   reg __398300_398300;
   reg _398301_398301 ; 
   reg __398301_398301;
   reg _398302_398302 ; 
   reg __398302_398302;
   reg _398303_398303 ; 
   reg __398303_398303;
   reg _398304_398304 ; 
   reg __398304_398304;
   reg _398305_398305 ; 
   reg __398305_398305;
   reg _398306_398306 ; 
   reg __398306_398306;
   reg _398307_398307 ; 
   reg __398307_398307;
   reg _398308_398308 ; 
   reg __398308_398308;
   reg _398309_398309 ; 
   reg __398309_398309;
   reg _398310_398310 ; 
   reg __398310_398310;
   reg _398311_398311 ; 
   reg __398311_398311;
   reg _398312_398312 ; 
   reg __398312_398312;
   reg _398313_398313 ; 
   reg __398313_398313;
   reg _398314_398314 ; 
   reg __398314_398314;
   reg _398315_398315 ; 
   reg __398315_398315;
   reg _398316_398316 ; 
   reg __398316_398316;
   reg _398317_398317 ; 
   reg __398317_398317;
   reg _398318_398318 ; 
   reg __398318_398318;
   reg _398319_398319 ; 
   reg __398319_398319;
   reg _398320_398320 ; 
   reg __398320_398320;
   reg _398321_398321 ; 
   reg __398321_398321;
   reg _398322_398322 ; 
   reg __398322_398322;
   reg _398323_398323 ; 
   reg __398323_398323;
   reg _398324_398324 ; 
   reg __398324_398324;
   reg _398325_398325 ; 
   reg __398325_398325;
   reg _398326_398326 ; 
   reg __398326_398326;
   reg _398327_398327 ; 
   reg __398327_398327;
   reg _398328_398328 ; 
   reg __398328_398328;
   reg _398329_398329 ; 
   reg __398329_398329;
   reg _398330_398330 ; 
   reg __398330_398330;
   reg _398331_398331 ; 
   reg __398331_398331;
   reg _398332_398332 ; 
   reg __398332_398332;
   reg _398333_398333 ; 
   reg __398333_398333;
   reg _398334_398334 ; 
   reg __398334_398334;
   reg _398335_398335 ; 
   reg __398335_398335;
   reg _398336_398336 ; 
   reg __398336_398336;
   reg _398337_398337 ; 
   reg __398337_398337;
   reg _398338_398338 ; 
   reg __398338_398338;
   reg _398339_398339 ; 
   reg __398339_398339;
   reg _398340_398340 ; 
   reg __398340_398340;
   reg _398341_398341 ; 
   reg __398341_398341;
   reg _398342_398342 ; 
   reg __398342_398342;
   reg _398343_398343 ; 
   reg __398343_398343;
   reg _398344_398344 ; 
   reg __398344_398344;
   reg _398345_398345 ; 
   reg __398345_398345;
   reg _398346_398346 ; 
   reg __398346_398346;
   reg _398347_398347 ; 
   reg __398347_398347;
   reg _398348_398348 ; 
   reg __398348_398348;
   reg _398349_398349 ; 
   reg __398349_398349;
   reg _398350_398350 ; 
   reg __398350_398350;
   reg _398351_398351 ; 
   reg __398351_398351;
   reg _398352_398352 ; 
   reg __398352_398352;
   reg _398353_398353 ; 
   reg __398353_398353;
   reg _398354_398354 ; 
   reg __398354_398354;
   reg _398355_398355 ; 
   reg __398355_398355;
   reg _398356_398356 ; 
   reg __398356_398356;
   reg _398357_398357 ; 
   reg __398357_398357;
   reg _398358_398358 ; 
   reg __398358_398358;
   reg _398359_398359 ; 
   reg __398359_398359;
   reg _398360_398360 ; 
   reg __398360_398360;
   reg _398361_398361 ; 
   reg __398361_398361;
   reg _398362_398362 ; 
   reg __398362_398362;
   reg _398363_398363 ; 
   reg __398363_398363;
   reg _398364_398364 ; 
   reg __398364_398364;
   reg _398365_398365 ; 
   reg __398365_398365;
   reg _398366_398366 ; 
   reg __398366_398366;
   reg _398367_398367 ; 
   reg __398367_398367;
   reg _398368_398368 ; 
   reg __398368_398368;
   reg _398369_398369 ; 
   reg __398369_398369;
   reg _398370_398370 ; 
   reg __398370_398370;
   reg _398371_398371 ; 
   reg __398371_398371;
   reg _398372_398372 ; 
   reg __398372_398372;
   reg _398373_398373 ; 
   reg __398373_398373;
   reg _398374_398374 ; 
   reg __398374_398374;
   reg _398375_398375 ; 
   reg __398375_398375;
   reg _398376_398376 ; 
   reg __398376_398376;
   reg _398377_398377 ; 
   reg __398377_398377;
   reg _398378_398378 ; 
   reg __398378_398378;
   reg _398379_398379 ; 
   reg __398379_398379;
   reg _398380_398380 ; 
   reg __398380_398380;
   reg _398381_398381 ; 
   reg __398381_398381;
   reg _398382_398382 ; 
   reg __398382_398382;
   reg _398383_398383 ; 
   reg __398383_398383;
   reg _398384_398384 ; 
   reg __398384_398384;
   reg _398385_398385 ; 
   reg __398385_398385;
   reg _398386_398386 ; 
   reg __398386_398386;
   reg _398387_398387 ; 
   reg __398387_398387;
   reg _398388_398388 ; 
   reg __398388_398388;
   reg _398389_398389 ; 
   reg __398389_398389;
   reg _398390_398390 ; 
   reg __398390_398390;
   reg _398391_398391 ; 
   reg __398391_398391;
   reg _398392_398392 ; 
   reg __398392_398392;
   reg _398393_398393 ; 
   reg __398393_398393;
   reg _398394_398394 ; 
   reg __398394_398394;
   reg _398395_398395 ; 
   reg __398395_398395;
   reg _398396_398396 ; 
   reg __398396_398396;
   reg _398397_398397 ; 
   reg __398397_398397;
   reg _398398_398398 ; 
   reg __398398_398398;
   reg _398399_398399 ; 
   reg __398399_398399;
   reg _398400_398400 ; 
   reg __398400_398400;
   reg _398401_398401 ; 
   reg __398401_398401;
   reg _398402_398402 ; 
   reg __398402_398402;
   reg _398403_398403 ; 
   reg __398403_398403;
   reg _398404_398404 ; 
   reg __398404_398404;
   reg _398405_398405 ; 
   reg __398405_398405;
   reg _398406_398406 ; 
   reg __398406_398406;
   reg _398407_398407 ; 
   reg __398407_398407;
   reg _398408_398408 ; 
   reg __398408_398408;
   reg _398409_398409 ; 
   reg __398409_398409;
   reg _398410_398410 ; 
   reg __398410_398410;
   reg _398411_398411 ; 
   reg __398411_398411;
   reg _398412_398412 ; 
   reg __398412_398412;
   reg _398413_398413 ; 
   reg __398413_398413;
   reg _398414_398414 ; 
   reg __398414_398414;
   reg _398415_398415 ; 
   reg __398415_398415;
   reg _398416_398416 ; 
   reg __398416_398416;
   reg _398417_398417 ; 
   reg __398417_398417;
   reg _398418_398418 ; 
   reg __398418_398418;
   reg _398419_398419 ; 
   reg __398419_398419;
   reg _398420_398420 ; 
   reg __398420_398420;
   reg _398421_398421 ; 
   reg __398421_398421;
   reg _398422_398422 ; 
   reg __398422_398422;
   reg _398423_398423 ; 
   reg __398423_398423;
   reg _398424_398424 ; 
   reg __398424_398424;
   reg _398425_398425 ; 
   reg __398425_398425;
   reg _398426_398426 ; 
   reg __398426_398426;
   reg _398427_398427 ; 
   reg __398427_398427;
   reg _398428_398428 ; 
   reg __398428_398428;
   reg _398429_398429 ; 
   reg __398429_398429;
   reg _398430_398430 ; 
   reg __398430_398430;
   reg _398431_398431 ; 
   reg __398431_398431;
   reg _398432_398432 ; 
   reg __398432_398432;
   reg _398433_398433 ; 
   reg __398433_398433;
   reg _398434_398434 ; 
   reg __398434_398434;
   reg _398435_398435 ; 
   reg __398435_398435;
   reg _398436_398436 ; 
   reg __398436_398436;
   reg _398437_398437 ; 
   reg __398437_398437;
   reg _398438_398438 ; 
   reg __398438_398438;
   reg _398439_398439 ; 
   reg __398439_398439;
   reg _398440_398440 ; 
   reg __398440_398440;
   reg _398441_398441 ; 
   reg __398441_398441;
   reg _398442_398442 ; 
   reg __398442_398442;
   reg _398443_398443 ; 
   reg __398443_398443;
   reg _398444_398444 ; 
   reg __398444_398444;
   reg _398445_398445 ; 
   reg __398445_398445;
   reg _398446_398446 ; 
   reg __398446_398446;
   reg _398447_398447 ; 
   reg __398447_398447;
   reg _398448_398448 ; 
   reg __398448_398448;
   reg _398449_398449 ; 
   reg __398449_398449;
   reg _398450_398450 ; 
   reg __398450_398450;
   reg _398451_398451 ; 
   reg __398451_398451;
   reg _398452_398452 ; 
   reg __398452_398452;
   reg _398453_398453 ; 
   reg __398453_398453;
   reg _398454_398454 ; 
   reg __398454_398454;
   reg _398455_398455 ; 
   reg __398455_398455;
   reg _398456_398456 ; 
   reg __398456_398456;
   reg _398457_398457 ; 
   reg __398457_398457;
   reg _398458_398458 ; 
   reg __398458_398458;
   reg _398459_398459 ; 
   reg __398459_398459;
   reg _398460_398460 ; 
   reg __398460_398460;
   reg _398461_398461 ; 
   reg __398461_398461;
   reg _398462_398462 ; 
   reg __398462_398462;
   reg _398463_398463 ; 
   reg __398463_398463;
   reg _398464_398464 ; 
   reg __398464_398464;
   reg _398465_398465 ; 
   reg __398465_398465;
   reg _398466_398466 ; 
   reg __398466_398466;
   reg _398467_398467 ; 
   reg __398467_398467;
   reg _398468_398468 ; 
   reg __398468_398468;
   reg _398469_398469 ; 
   reg __398469_398469;
   reg _398470_398470 ; 
   reg __398470_398470;
   reg _398471_398471 ; 
   reg __398471_398471;
   reg _398472_398472 ; 
   reg __398472_398472;
   reg _398473_398473 ; 
   reg __398473_398473;
   reg _398474_398474 ; 
   reg __398474_398474;
   reg _398475_398475 ; 
   reg __398475_398475;
   reg _398476_398476 ; 
   reg __398476_398476;
   reg _398477_398477 ; 
   reg __398477_398477;
   reg _398478_398478 ; 
   reg __398478_398478;
   reg _398479_398479 ; 
   reg __398479_398479;
   reg _398480_398480 ; 
   reg __398480_398480;
   reg _398481_398481 ; 
   reg __398481_398481;
   reg _398482_398482 ; 
   reg __398482_398482;
   reg _398483_398483 ; 
   reg __398483_398483;
   reg _398484_398484 ; 
   reg __398484_398484;
   reg _398485_398485 ; 
   reg __398485_398485;
   reg _398486_398486 ; 
   reg __398486_398486;
   reg _398487_398487 ; 
   reg __398487_398487;
   reg _398488_398488 ; 
   reg __398488_398488;
   reg _398489_398489 ; 
   reg __398489_398489;
   reg _398490_398490 ; 
   reg __398490_398490;
   reg _398491_398491 ; 
   reg __398491_398491;
   reg _398492_398492 ; 
   reg __398492_398492;
   reg _398493_398493 ; 
   reg __398493_398493;
   reg _398494_398494 ; 
   reg __398494_398494;
   reg _398495_398495 ; 
   reg __398495_398495;
   reg _398496_398496 ; 
   reg __398496_398496;
   reg _398497_398497 ; 
   reg __398497_398497;
   reg _398498_398498 ; 
   reg __398498_398498;
   reg _398499_398499 ; 
   reg __398499_398499;
   reg _398500_398500 ; 
   reg __398500_398500;
   reg _398501_398501 ; 
   reg __398501_398501;
   reg _398502_398502 ; 
   reg __398502_398502;
   reg _398503_398503 ; 
   reg __398503_398503;
   reg _398504_398504 ; 
   reg __398504_398504;
   reg _398505_398505 ; 
   reg __398505_398505;
   reg _398506_398506 ; 
   reg __398506_398506;
   reg _398507_398507 ; 
   reg __398507_398507;
   reg _398508_398508 ; 
   reg __398508_398508;
   reg _398509_398509 ; 
   reg __398509_398509;
   reg _398510_398510 ; 
   reg __398510_398510;
   reg _398511_398511 ; 
   reg __398511_398511;
   reg _398512_398512 ; 
   reg __398512_398512;
   reg _398513_398513 ; 
   reg __398513_398513;
   reg _398514_398514 ; 
   reg __398514_398514;
   reg _398515_398515 ; 
   reg __398515_398515;
   reg _398516_398516 ; 
   reg __398516_398516;
   reg _398517_398517 ; 
   reg __398517_398517;
   reg _398518_398518 ; 
   reg __398518_398518;
   reg _398519_398519 ; 
   reg __398519_398519;
   reg _398520_398520 ; 
   reg __398520_398520;
   reg _398521_398521 ; 
   reg __398521_398521;
   reg _398522_398522 ; 
   reg __398522_398522;
   reg _398523_398523 ; 
   reg __398523_398523;
   reg _398524_398524 ; 
   reg __398524_398524;
   reg _398525_398525 ; 
   reg __398525_398525;
   reg _398526_398526 ; 
   reg __398526_398526;
   reg _398527_398527 ; 
   reg __398527_398527;
   reg _398528_398528 ; 
   reg __398528_398528;
   reg _398529_398529 ; 
   reg __398529_398529;
   reg _398530_398530 ; 
   reg __398530_398530;
   reg _398531_398531 ; 
   reg __398531_398531;
   reg _398532_398532 ; 
   reg __398532_398532;
   reg _398533_398533 ; 
   reg __398533_398533;
   reg _398534_398534 ; 
   reg __398534_398534;
   reg _398535_398535 ; 
   reg __398535_398535;
   reg _398536_398536 ; 
   reg __398536_398536;
   reg _398537_398537 ; 
   reg __398537_398537;
   reg _398538_398538 ; 
   reg __398538_398538;
   reg _398539_398539 ; 
   reg __398539_398539;
   reg _398540_398540 ; 
   reg __398540_398540;
   reg _398541_398541 ; 
   reg __398541_398541;
   reg _398542_398542 ; 
   reg __398542_398542;
   reg _398543_398543 ; 
   reg __398543_398543;
   reg _398544_398544 ; 
   reg __398544_398544;
   reg _398545_398545 ; 
   reg __398545_398545;
   reg _398546_398546 ; 
   reg __398546_398546;
   reg _398547_398547 ; 
   reg __398547_398547;
   reg _398548_398548 ; 
   reg __398548_398548;
   reg _398549_398549 ; 
   reg __398549_398549;
   reg _398550_398550 ; 
   reg __398550_398550;
   reg _398551_398551 ; 
   reg __398551_398551;
   reg _398552_398552 ; 
   reg __398552_398552;
   reg _398553_398553 ; 
   reg __398553_398553;
   reg _398554_398554 ; 
   reg __398554_398554;
   reg _398555_398555 ; 
   reg __398555_398555;
   reg _398556_398556 ; 
   reg __398556_398556;
   reg _398557_398557 ; 
   reg __398557_398557;
   reg _398558_398558 ; 
   reg __398558_398558;
   reg _398559_398559 ; 
   reg __398559_398559;
   reg _398560_398560 ; 
   reg __398560_398560;
   reg _398561_398561 ; 
   reg __398561_398561;
   reg _398562_398562 ; 
   reg __398562_398562;
   reg _398563_398563 ; 
   reg __398563_398563;
   reg _398564_398564 ; 
   reg __398564_398564;
   reg _398565_398565 ; 
   reg __398565_398565;
   reg _398566_398566 ; 
   reg __398566_398566;
   reg _398567_398567 ; 
   reg __398567_398567;
   reg _398568_398568 ; 
   reg __398568_398568;
   reg _398569_398569 ; 
   reg __398569_398569;
   reg _398570_398570 ; 
   reg __398570_398570;
   reg _398571_398571 ; 
   reg __398571_398571;
   reg _398572_398572 ; 
   reg __398572_398572;
   reg _398573_398573 ; 
   reg __398573_398573;
   reg _398574_398574 ; 
   reg __398574_398574;
   reg _398575_398575 ; 
   reg __398575_398575;
   reg _398576_398576 ; 
   reg __398576_398576;
   reg _398577_398577 ; 
   reg __398577_398577;
   reg _398578_398578 ; 
   reg __398578_398578;
   reg _398579_398579 ; 
   reg __398579_398579;
   reg _398580_398580 ; 
   reg __398580_398580;
   reg _398581_398581 ; 
   reg __398581_398581;
   reg _398582_398582 ; 
   reg __398582_398582;
   reg _398583_398583 ; 
   reg __398583_398583;
   reg _398584_398584 ; 
   reg __398584_398584;
   reg _398585_398585 ; 
   reg __398585_398585;
   reg _398586_398586 ; 
   reg __398586_398586;
   reg _398587_398587 ; 
   reg __398587_398587;
   reg _398588_398588 ; 
   reg __398588_398588;
   reg _398589_398589 ; 
   reg __398589_398589;
   reg _398590_398590 ; 
   reg __398590_398590;
   reg _398591_398591 ; 
   reg __398591_398591;
   reg _398592_398592 ; 
   reg __398592_398592;
   reg _398593_398593 ; 
   reg __398593_398593;
   reg _398594_398594 ; 
   reg __398594_398594;
   reg _398595_398595 ; 
   reg __398595_398595;
   reg _398596_398596 ; 
   reg __398596_398596;
   reg _398597_398597 ; 
   reg __398597_398597;
   reg _398598_398598 ; 
   reg __398598_398598;
   reg _398599_398599 ; 
   reg __398599_398599;
   reg _398600_398600 ; 
   reg __398600_398600;
   reg _398601_398601 ; 
   reg __398601_398601;
   reg _398602_398602 ; 
   reg __398602_398602;
   reg _398603_398603 ; 
   reg __398603_398603;
   reg _398604_398604 ; 
   reg __398604_398604;
   reg _398605_398605 ; 
   reg __398605_398605;
   reg _398606_398606 ; 
   reg __398606_398606;
   reg _398607_398607 ; 
   reg __398607_398607;
   reg _398608_398608 ; 
   reg __398608_398608;
   reg _398609_398609 ; 
   reg __398609_398609;
   reg _398610_398610 ; 
   reg __398610_398610;
   reg _398611_398611 ; 
   reg __398611_398611;
   reg _398612_398612 ; 
   reg __398612_398612;
   reg _398613_398613 ; 
   reg __398613_398613;
   reg _398614_398614 ; 
   reg __398614_398614;
   reg _398615_398615 ; 
   reg __398615_398615;
   reg _398616_398616 ; 
   reg __398616_398616;
   reg _398617_398617 ; 
   reg __398617_398617;
   reg _398618_398618 ; 
   reg __398618_398618;
   reg _398619_398619 ; 
   reg __398619_398619;
   reg _398620_398620 ; 
   reg __398620_398620;
   reg _398621_398621 ; 
   reg __398621_398621;
   reg _398622_398622 ; 
   reg __398622_398622;
   reg _398623_398623 ; 
   reg __398623_398623;
   reg _398624_398624 ; 
   reg __398624_398624;
   reg _398625_398625 ; 
   reg __398625_398625;
   reg _398626_398626 ; 
   reg __398626_398626;
   reg _398627_398627 ; 
   reg __398627_398627;
   reg _398628_398628 ; 
   reg __398628_398628;
   reg _398629_398629 ; 
   reg __398629_398629;
   reg _398630_398630 ; 
   reg __398630_398630;
   reg _398631_398631 ; 
   reg __398631_398631;
   reg _398632_398632 ; 
   reg __398632_398632;
   reg _398633_398633 ; 
   reg __398633_398633;
   reg _398634_398634 ; 
   reg __398634_398634;
   reg _398635_398635 ; 
   reg __398635_398635;
   reg _398636_398636 ; 
   reg __398636_398636;
   reg _398637_398637 ; 
   reg __398637_398637;
   reg _398638_398638 ; 
   reg __398638_398638;
   reg _398639_398639 ; 
   reg __398639_398639;
   reg _398640_398640 ; 
   reg __398640_398640;
   reg _398641_398641 ; 
   reg __398641_398641;
   reg _398642_398642 ; 
   reg __398642_398642;
   reg _398643_398643 ; 
   reg __398643_398643;
   reg _398644_398644 ; 
   reg __398644_398644;
   reg _398645_398645 ; 
   reg __398645_398645;
   reg _398646_398646 ; 
   reg __398646_398646;
   reg _398647_398647 ; 
   reg __398647_398647;
   reg _398648_398648 ; 
   reg __398648_398648;
   reg _398649_398649 ; 
   reg __398649_398649;
   reg _398650_398650 ; 
   reg __398650_398650;
   reg _398651_398651 ; 
   reg __398651_398651;
   reg _398652_398652 ; 
   reg __398652_398652;
   reg _398653_398653 ; 
   reg __398653_398653;
   reg _398654_398654 ; 
   reg __398654_398654;
   reg _398655_398655 ; 
   reg __398655_398655;
   reg _398656_398656 ; 
   reg __398656_398656;
   reg _398657_398657 ; 
   reg __398657_398657;
   reg _398658_398658 ; 
   reg __398658_398658;
   reg _398659_398659 ; 
   reg __398659_398659;
   reg _398660_398660 ; 
   reg __398660_398660;
   reg _398661_398661 ; 
   reg __398661_398661;
   reg _398662_398662 ; 
   reg __398662_398662;
   reg _398663_398663 ; 
   reg __398663_398663;
   reg _398664_398664 ; 
   reg __398664_398664;
   reg _398665_398665 ; 
   reg __398665_398665;
   reg _398666_398666 ; 
   reg __398666_398666;
   reg _398667_398667 ; 
   reg __398667_398667;
   reg _398668_398668 ; 
   reg __398668_398668;
   reg _398669_398669 ; 
   reg __398669_398669;
   reg _398670_398670 ; 
   reg __398670_398670;
   reg _398671_398671 ; 
   reg __398671_398671;
   reg _398672_398672 ; 
   reg __398672_398672;
   reg _398673_398673 ; 
   reg __398673_398673;
   reg _398674_398674 ; 
   reg __398674_398674;
   reg _398675_398675 ; 
   reg __398675_398675;
   reg _398676_398676 ; 
   reg __398676_398676;
   reg _398677_398677 ; 
   reg __398677_398677;
   reg _398678_398678 ; 
   reg __398678_398678;
   reg _398679_398679 ; 
   reg __398679_398679;
   reg _398680_398680 ; 
   reg __398680_398680;
   reg _398681_398681 ; 
   reg __398681_398681;
   reg _398682_398682 ; 
   reg __398682_398682;
   reg _398683_398683 ; 
   reg __398683_398683;
   reg _398684_398684 ; 
   reg __398684_398684;
   reg _398685_398685 ; 
   reg __398685_398685;
   reg _398686_398686 ; 
   reg __398686_398686;
   reg _398687_398687 ; 
   reg __398687_398687;
   reg _398688_398688 ; 
   reg __398688_398688;
   reg _398689_398689 ; 
   reg __398689_398689;
   reg _398690_398690 ; 
   reg __398690_398690;
   reg _398691_398691 ; 
   reg __398691_398691;
   reg _398692_398692 ; 
   reg __398692_398692;
   reg _398693_398693 ; 
   reg __398693_398693;
   reg _398694_398694 ; 
   reg __398694_398694;
   reg _398695_398695 ; 
   reg __398695_398695;
   reg _398696_398696 ; 
   reg __398696_398696;
   reg _398697_398697 ; 
   reg __398697_398697;
   reg _398698_398698 ; 
   reg __398698_398698;
   reg _398699_398699 ; 
   reg __398699_398699;
   reg _398700_398700 ; 
   reg __398700_398700;
   reg _398701_398701 ; 
   reg __398701_398701;
   reg _398702_398702 ; 
   reg __398702_398702;
   reg _398703_398703 ; 
   reg __398703_398703;
   reg _398704_398704 ; 
   reg __398704_398704;
   reg _398705_398705 ; 
   reg __398705_398705;
   reg _398706_398706 ; 
   reg __398706_398706;
   reg _398707_398707 ; 
   reg __398707_398707;
   reg _398708_398708 ; 
   reg __398708_398708;
   reg _398709_398709 ; 
   reg __398709_398709;
   reg _398710_398710 ; 
   reg __398710_398710;
   reg _398711_398711 ; 
   reg __398711_398711;
   reg _398712_398712 ; 
   reg __398712_398712;
   reg _398713_398713 ; 
   reg __398713_398713;
   reg _398714_398714 ; 
   reg __398714_398714;
   reg _398715_398715 ; 
   reg __398715_398715;
   reg _398716_398716 ; 
   reg __398716_398716;
   reg _398717_398717 ; 
   reg __398717_398717;
   reg _398718_398718 ; 
   reg __398718_398718;
   reg _398719_398719 ; 
   reg __398719_398719;
   reg _398720_398720 ; 
   reg __398720_398720;
   reg _398721_398721 ; 
   reg __398721_398721;
   reg _398722_398722 ; 
   reg __398722_398722;
   reg _398723_398723 ; 
   reg __398723_398723;
   reg _398724_398724 ; 
   reg __398724_398724;
   reg _398725_398725 ; 
   reg __398725_398725;
   reg _398726_398726 ; 
   reg __398726_398726;
   reg _398727_398727 ; 
   reg __398727_398727;
   reg _398728_398728 ; 
   reg __398728_398728;
   reg _398729_398729 ; 
   reg __398729_398729;
   reg _398730_398730 ; 
   reg __398730_398730;
   reg _398731_398731 ; 
   reg __398731_398731;
   reg _398732_398732 ; 
   reg __398732_398732;
   reg _398733_398733 ; 
   reg __398733_398733;
   reg _398734_398734 ; 
   reg __398734_398734;
   reg _398735_398735 ; 
   reg __398735_398735;
   reg _398736_398736 ; 
   reg __398736_398736;
   reg _398737_398737 ; 
   reg __398737_398737;
   reg _398738_398738 ; 
   reg __398738_398738;
   reg _398739_398739 ; 
   reg __398739_398739;
   reg _398740_398740 ; 
   reg __398740_398740;
   reg _398741_398741 ; 
   reg __398741_398741;
   reg _398742_398742 ; 
   reg __398742_398742;
   reg _398743_398743 ; 
   reg __398743_398743;
   reg _398744_398744 ; 
   reg __398744_398744;
   reg _398745_398745 ; 
   reg __398745_398745;
   reg _398746_398746 ; 
   reg __398746_398746;
   reg _398747_398747 ; 
   reg __398747_398747;
   reg _398748_398748 ; 
   reg __398748_398748;
   reg _398749_398749 ; 
   reg __398749_398749;
   reg _398750_398750 ; 
   reg __398750_398750;
   reg _398751_398751 ; 
   reg __398751_398751;
   reg _398752_398752 ; 
   reg __398752_398752;
   reg _398753_398753 ; 
   reg __398753_398753;
   reg _398754_398754 ; 
   reg __398754_398754;
   reg _398755_398755 ; 
   reg __398755_398755;
   reg _398756_398756 ; 
   reg __398756_398756;
   reg _398757_398757 ; 
   reg __398757_398757;
   reg _398758_398758 ; 
   reg __398758_398758;
   reg _398759_398759 ; 
   reg __398759_398759;
   reg _398760_398760 ; 
   reg __398760_398760;
   reg _398761_398761 ; 
   reg __398761_398761;
   reg _398762_398762 ; 
   reg __398762_398762;
   reg _398763_398763 ; 
   reg __398763_398763;
   reg _398764_398764 ; 
   reg __398764_398764;
   reg _398765_398765 ; 
   reg __398765_398765;
   reg _398766_398766 ; 
   reg __398766_398766;
   reg _398767_398767 ; 
   reg __398767_398767;
   reg _398768_398768 ; 
   reg __398768_398768;
   reg _398769_398769 ; 
   reg __398769_398769;
   reg _398770_398770 ; 
   reg __398770_398770;
   reg _398771_398771 ; 
   reg __398771_398771;
   reg _398772_398772 ; 
   reg __398772_398772;
   reg _398773_398773 ; 
   reg __398773_398773;
   reg _398774_398774 ; 
   reg __398774_398774;
   reg _398775_398775 ; 
   reg __398775_398775;
   reg _398776_398776 ; 
   reg __398776_398776;
   reg _398777_398777 ; 
   reg __398777_398777;
   reg _398778_398778 ; 
   reg __398778_398778;
   reg _398779_398779 ; 
   reg __398779_398779;
   reg _398780_398780 ; 
   reg __398780_398780;
   reg _398781_398781 ; 
   reg __398781_398781;
   reg _398782_398782 ; 
   reg __398782_398782;
   reg _398783_398783 ; 
   reg __398783_398783;
   reg _398784_398784 ; 
   reg __398784_398784;
   reg _398785_398785 ; 
   reg __398785_398785;
   reg _398786_398786 ; 
   reg __398786_398786;
   reg _398787_398787 ; 
   reg __398787_398787;
   reg _398788_398788 ; 
   reg __398788_398788;
   reg _398789_398789 ; 
   reg __398789_398789;
   reg _398790_398790 ; 
   reg __398790_398790;
   reg _398791_398791 ; 
   reg __398791_398791;
   reg _398792_398792 ; 
   reg __398792_398792;
   reg _398793_398793 ; 
   reg __398793_398793;
   reg _398794_398794 ; 
   reg __398794_398794;
   reg _398795_398795 ; 
   reg __398795_398795;
   reg _398796_398796 ; 
   reg __398796_398796;
   reg _398797_398797 ; 
   reg __398797_398797;
   reg _398798_398798 ; 
   reg __398798_398798;
   reg _398799_398799 ; 
   reg __398799_398799;
   reg _398800_398800 ; 
   reg __398800_398800;
   reg _398801_398801 ; 
   reg __398801_398801;
   reg _398802_398802 ; 
   reg __398802_398802;
   reg _398803_398803 ; 
   reg __398803_398803;
   reg _398804_398804 ; 
   reg __398804_398804;
   reg _398805_398805 ; 
   reg __398805_398805;
   reg _398806_398806 ; 
   reg __398806_398806;
   reg _398807_398807 ; 
   reg __398807_398807;
   reg _398808_398808 ; 
   reg __398808_398808;
   reg _398809_398809 ; 
   reg __398809_398809;
   reg _398810_398810 ; 
   reg __398810_398810;
   reg _398811_398811 ; 
   reg __398811_398811;
   reg _398812_398812 ; 
   reg __398812_398812;
   reg _398813_398813 ; 
   reg __398813_398813;
   reg _398814_398814 ; 
   reg __398814_398814;
   reg _398815_398815 ; 
   reg __398815_398815;
   reg _398816_398816 ; 
   reg __398816_398816;
   reg _398817_398817 ; 
   reg __398817_398817;
   reg _398818_398818 ; 
   reg __398818_398818;
   reg _398819_398819 ; 
   reg __398819_398819;
   reg _398820_398820 ; 
   reg __398820_398820;
   reg _398821_398821 ; 
   reg __398821_398821;
   reg _398822_398822 ; 
   reg __398822_398822;
   reg _398823_398823 ; 
   reg __398823_398823;
   reg _398824_398824 ; 
   reg __398824_398824;
   reg _398825_398825 ; 
   reg __398825_398825;
   reg _398826_398826 ; 
   reg __398826_398826;
   reg _398827_398827 ; 
   reg __398827_398827;
   reg _398828_398828 ; 
   reg __398828_398828;
   reg _398829_398829 ; 
   reg __398829_398829;
   reg _398830_398830 ; 
   reg __398830_398830;
   reg _398831_398831 ; 
   reg __398831_398831;
   reg _398832_398832 ; 
   reg __398832_398832;
   reg _398833_398833 ; 
   reg __398833_398833;
   reg _398834_398834 ; 
   reg __398834_398834;
   reg _398835_398835 ; 
   reg __398835_398835;
   reg _398836_398836 ; 
   reg __398836_398836;
   reg _398837_398837 ; 
   reg __398837_398837;
   reg _398838_398838 ; 
   reg __398838_398838;
   reg _398839_398839 ; 
   reg __398839_398839;
   reg _398840_398840 ; 
   reg __398840_398840;
   reg _398841_398841 ; 
   reg __398841_398841;
   reg _398842_398842 ; 
   reg __398842_398842;
   reg _398843_398843 ; 
   reg __398843_398843;
   reg _398844_398844 ; 
   reg __398844_398844;
   reg _398845_398845 ; 
   reg __398845_398845;
   reg _398846_398846 ; 
   reg __398846_398846;
   reg _398847_398847 ; 
   reg __398847_398847;
   reg _398848_398848 ; 
   reg __398848_398848;
   reg _398849_398849 ; 
   reg __398849_398849;
   reg _398850_398850 ; 
   reg __398850_398850;
   reg _398851_398851 ; 
   reg __398851_398851;
   reg _398852_398852 ; 
   reg __398852_398852;
   reg _398853_398853 ; 
   reg __398853_398853;
   reg _398854_398854 ; 
   reg __398854_398854;
   reg _398855_398855 ; 
   reg __398855_398855;
   reg _398856_398856 ; 
   reg __398856_398856;
   reg _398857_398857 ; 
   reg __398857_398857;
   reg _398858_398858 ; 
   reg __398858_398858;
   reg _398859_398859 ; 
   reg __398859_398859;
   reg _398860_398860 ; 
   reg __398860_398860;
   reg _398861_398861 ; 
   reg __398861_398861;
   reg _398862_398862 ; 
   reg __398862_398862;
   reg _398863_398863 ; 
   reg __398863_398863;
   reg _398864_398864 ; 
   reg __398864_398864;
   reg _398865_398865 ; 
   reg __398865_398865;
   reg _398866_398866 ; 
   reg __398866_398866;
   reg _398867_398867 ; 
   reg __398867_398867;
   reg _398868_398868 ; 
   reg __398868_398868;
   reg _398869_398869 ; 
   reg __398869_398869;
   reg _398870_398870 ; 
   reg __398870_398870;
   reg _398871_398871 ; 
   reg __398871_398871;
   reg _398872_398872 ; 
   reg __398872_398872;
   reg _398873_398873 ; 
   reg __398873_398873;
   reg _398874_398874 ; 
   reg __398874_398874;
   reg _398875_398875 ; 
   reg __398875_398875;
   reg _398876_398876 ; 
   reg __398876_398876;
   reg _398877_398877 ; 
   reg __398877_398877;
   reg _398878_398878 ; 
   reg __398878_398878;
   reg _398879_398879 ; 
   reg __398879_398879;
   reg _398880_398880 ; 
   reg __398880_398880;
   reg _398881_398881 ; 
   reg __398881_398881;
   reg _398882_398882 ; 
   reg __398882_398882;
   reg _398883_398883 ; 
   reg __398883_398883;
   reg _398884_398884 ; 
   reg __398884_398884;
   reg _398885_398885 ; 
   reg __398885_398885;
   reg _398886_398886 ; 
   reg __398886_398886;
   reg _398887_398887 ; 
   reg __398887_398887;
   reg _398888_398888 ; 
   reg __398888_398888;
   reg _398889_398889 ; 
   reg __398889_398889;
   reg _398890_398890 ; 
   reg __398890_398890;
   reg _398891_398891 ; 
   reg __398891_398891;
   reg _398892_398892 ; 
   reg __398892_398892;
   reg _398893_398893 ; 
   reg __398893_398893;
   reg _398894_398894 ; 
   reg __398894_398894;
   reg _398895_398895 ; 
   reg __398895_398895;
   reg _398896_398896 ; 
   reg __398896_398896;
   reg _398897_398897 ; 
   reg __398897_398897;
   reg _398898_398898 ; 
   reg __398898_398898;
   reg _398899_398899 ; 
   reg __398899_398899;
   reg _398900_398900 ; 
   reg __398900_398900;
   reg _398901_398901 ; 
   reg __398901_398901;
   reg _398902_398902 ; 
   reg __398902_398902;
   reg _398903_398903 ; 
   reg __398903_398903;
   reg _398904_398904 ; 
   reg __398904_398904;
   reg _398905_398905 ; 
   reg __398905_398905;
   reg _398906_398906 ; 
   reg __398906_398906;
   reg _398907_398907 ; 
   reg __398907_398907;
   reg _398908_398908 ; 
   reg __398908_398908;
   reg _398909_398909 ; 
   reg __398909_398909;
   reg _398910_398910 ; 
   reg __398910_398910;
   reg _398911_398911 ; 
   reg __398911_398911;
   reg _398912_398912 ; 
   reg __398912_398912;
   reg _398913_398913 ; 
   reg __398913_398913;
   reg _398914_398914 ; 
   reg __398914_398914;
   reg _398915_398915 ; 
   reg __398915_398915;
   reg _398916_398916 ; 
   reg __398916_398916;
   reg _398917_398917 ; 
   reg __398917_398917;
   reg _398918_398918 ; 
   reg __398918_398918;
   reg _398919_398919 ; 
   reg __398919_398919;
   reg _398920_398920 ; 
   reg __398920_398920;
   reg _398921_398921 ; 
   reg __398921_398921;
   reg _398922_398922 ; 
   reg __398922_398922;
   reg _398923_398923 ; 
   reg __398923_398923;
   reg _398924_398924 ; 
   reg __398924_398924;
   reg _398925_398925 ; 
   reg __398925_398925;
   reg _398926_398926 ; 
   reg __398926_398926;
   reg _398927_398927 ; 
   reg __398927_398927;
   reg _398928_398928 ; 
   reg __398928_398928;
   reg _398929_398929 ; 
   reg __398929_398929;
   reg _398930_398930 ; 
   reg __398930_398930;
   reg _398931_398931 ; 
   reg __398931_398931;
   reg _398932_398932 ; 
   reg __398932_398932;
   reg _398933_398933 ; 
   reg __398933_398933;
   reg _398934_398934 ; 
   reg __398934_398934;
   reg _398935_398935 ; 
   reg __398935_398935;
   reg _398936_398936 ; 
   reg __398936_398936;
   reg _398937_398937 ; 
   reg __398937_398937;
   reg _398938_398938 ; 
   reg __398938_398938;
   reg _398939_398939 ; 
   reg __398939_398939;
   reg _398940_398940 ; 
   reg __398940_398940;
   reg _398941_398941 ; 
   reg __398941_398941;
   reg _398942_398942 ; 
   reg __398942_398942;
   reg _398943_398943 ; 
   reg __398943_398943;
   reg _398944_398944 ; 
   reg __398944_398944;
   reg _398945_398945 ; 
   reg __398945_398945;
   reg _398946_398946 ; 
   reg __398946_398946;
   reg _398947_398947 ; 
   reg __398947_398947;
   reg _398948_398948 ; 
   reg __398948_398948;
   reg _398949_398949 ; 
   reg __398949_398949;
   reg _398950_398950 ; 
   reg __398950_398950;
   reg _398951_398951 ; 
   reg __398951_398951;
   reg _398952_398952 ; 
   reg __398952_398952;
   reg _398953_398953 ; 
   reg __398953_398953;
   reg _398954_398954 ; 
   reg __398954_398954;
   reg _398955_398955 ; 
   reg __398955_398955;
   reg _398956_398956 ; 
   reg __398956_398956;
   reg _398957_398957 ; 
   reg __398957_398957;
   reg _398958_398958 ; 
   reg __398958_398958;
   reg _398959_398959 ; 
   reg __398959_398959;
   reg _398960_398960 ; 
   reg __398960_398960;
   reg _398961_398961 ; 
   reg __398961_398961;
   reg _398962_398962 ; 
   reg __398962_398962;
   reg _398963_398963 ; 
   reg __398963_398963;
   reg _398964_398964 ; 
   reg __398964_398964;
   reg _398965_398965 ; 
   reg __398965_398965;
   reg _398966_398966 ; 
   reg __398966_398966;
   reg _398967_398967 ; 
   reg __398967_398967;
   reg _398968_398968 ; 
   reg __398968_398968;
   reg _398969_398969 ; 
   reg __398969_398969;
   reg _398970_398970 ; 
   reg __398970_398970;
   reg _398971_398971 ; 
   reg __398971_398971;
   reg _398972_398972 ; 
   reg __398972_398972;
   reg _398973_398973 ; 
   reg __398973_398973;
   reg _398974_398974 ; 
   reg __398974_398974;
   reg _398975_398975 ; 
   reg __398975_398975;
   reg _398976_398976 ; 
   reg __398976_398976;
   reg _398977_398977 ; 
   reg __398977_398977;
   reg _398978_398978 ; 
   reg __398978_398978;
   reg _398979_398979 ; 
   reg __398979_398979;
   reg _398980_398980 ; 
   reg __398980_398980;
   reg _398981_398981 ; 
   reg __398981_398981;
   reg _398982_398982 ; 
   reg __398982_398982;
   reg _398983_398983 ; 
   reg __398983_398983;
   reg _398984_398984 ; 
   reg __398984_398984;
   reg _398985_398985 ; 
   reg __398985_398985;
   reg _398986_398986 ; 
   reg __398986_398986;
   reg _398987_398987 ; 
   reg __398987_398987;
   reg _398988_398988 ; 
   reg __398988_398988;
   reg _398989_398989 ; 
   reg __398989_398989;
   reg _398990_398990 ; 
   reg __398990_398990;
   reg _398991_398991 ; 
   reg __398991_398991;
   reg _398992_398992 ; 
   reg __398992_398992;
   reg _398993_398993 ; 
   reg __398993_398993;
   reg _398994_398994 ; 
   reg __398994_398994;
   reg _398995_398995 ; 
   reg __398995_398995;
   reg _398996_398996 ; 
   reg __398996_398996;
   reg _398997_398997 ; 
   reg __398997_398997;
   reg _398998_398998 ; 
   reg __398998_398998;
   reg _398999_398999 ; 
   reg __398999_398999;
   reg _399000_399000 ; 
   reg __399000_399000;
   reg _399001_399001 ; 
   reg __399001_399001;
   reg _399002_399002 ; 
   reg __399002_399002;
   reg _399003_399003 ; 
   reg __399003_399003;
   reg _399004_399004 ; 
   reg __399004_399004;
   reg _399005_399005 ; 
   reg __399005_399005;
   reg _399006_399006 ; 
   reg __399006_399006;
   reg _399007_399007 ; 
   reg __399007_399007;
   reg _399008_399008 ; 
   reg __399008_399008;
   reg _399009_399009 ; 
   reg __399009_399009;
   reg _399010_399010 ; 
   reg __399010_399010;
   reg _399011_399011 ; 
   reg __399011_399011;
   reg _399012_399012 ; 
   reg __399012_399012;
   reg _399013_399013 ; 
   reg __399013_399013;
   reg _399014_399014 ; 
   reg __399014_399014;
   reg _399015_399015 ; 
   reg __399015_399015;
   reg _399016_399016 ; 
   reg __399016_399016;
   reg _399017_399017 ; 
   reg __399017_399017;
   reg _399018_399018 ; 
   reg __399018_399018;
   reg _399019_399019 ; 
   reg __399019_399019;
   reg _399020_399020 ; 
   reg __399020_399020;
   reg _399021_399021 ; 
   reg __399021_399021;
   reg _399022_399022 ; 
   reg __399022_399022;
   reg _399023_399023 ; 
   reg __399023_399023;
   reg _399024_399024 ; 
   reg __399024_399024;
   reg _399025_399025 ; 
   reg __399025_399025;
   reg _399026_399026 ; 
   reg __399026_399026;
   reg _399027_399027 ; 
   reg __399027_399027;
   reg _399028_399028 ; 
   reg __399028_399028;
   reg _399029_399029 ; 
   reg __399029_399029;
   reg _399030_399030 ; 
   reg __399030_399030;
   reg _399031_399031 ; 
   reg __399031_399031;
   reg _399032_399032 ; 
   reg __399032_399032;
   reg _399033_399033 ; 
   reg __399033_399033;
   reg _399034_399034 ; 
   reg __399034_399034;
   reg _399035_399035 ; 
   reg __399035_399035;
   reg _399036_399036 ; 
   reg __399036_399036;
   reg _399037_399037 ; 
   reg __399037_399037;
   reg _399038_399038 ; 
   reg __399038_399038;
   reg _399039_399039 ; 
   reg __399039_399039;
   reg _399040_399040 ; 
   reg __399040_399040;
   reg _399041_399041 ; 
   reg __399041_399041;
   reg _399042_399042 ; 
   reg __399042_399042;
   reg _399043_399043 ; 
   reg __399043_399043;
   reg _399044_399044 ; 
   reg __399044_399044;
   reg _399045_399045 ; 
   reg __399045_399045;
   reg _399046_399046 ; 
   reg __399046_399046;
   reg _399047_399047 ; 
   reg __399047_399047;
   reg _399048_399048 ; 
   reg __399048_399048;
   reg _399049_399049 ; 
   reg __399049_399049;
   reg _399050_399050 ; 
   reg __399050_399050;
   reg _399051_399051 ; 
   reg __399051_399051;
   reg _399052_399052 ; 
   reg __399052_399052;
   reg _399053_399053 ; 
   reg __399053_399053;
   reg _399054_399054 ; 
   reg __399054_399054;
   reg _399055_399055 ; 
   reg __399055_399055;
   reg _399056_399056 ; 
   reg __399056_399056;
   reg _399057_399057 ; 
   reg __399057_399057;
   reg _399058_399058 ; 
   reg __399058_399058;
   reg _399059_399059 ; 
   reg __399059_399059;
   reg _399060_399060 ; 
   reg __399060_399060;
   reg _399061_399061 ; 
   reg __399061_399061;
   reg _399062_399062 ; 
   reg __399062_399062;
   reg _399063_399063 ; 
   reg __399063_399063;
   reg _399064_399064 ; 
   reg __399064_399064;
   reg _399065_399065 ; 
   reg __399065_399065;
   reg _399066_399066 ; 
   reg __399066_399066;
   reg _399067_399067 ; 
   reg __399067_399067;
   reg _399068_399068 ; 
   reg __399068_399068;
   reg _399069_399069 ; 
   reg __399069_399069;
   reg _399070_399070 ; 
   reg __399070_399070;
   reg _399071_399071 ; 
   reg __399071_399071;
   reg _399072_399072 ; 
   reg __399072_399072;
   reg _399073_399073 ; 
   reg __399073_399073;
   reg _399074_399074 ; 
   reg __399074_399074;
   reg _399075_399075 ; 
   reg __399075_399075;
   reg _399076_399076 ; 
   reg __399076_399076;
   reg _399077_399077 ; 
   reg __399077_399077;
   reg _399078_399078 ; 
   reg __399078_399078;
   reg _399079_399079 ; 
   reg __399079_399079;
   reg _399080_399080 ; 
   reg __399080_399080;
   reg _399081_399081 ; 
   reg __399081_399081;
   reg _399082_399082 ; 
   reg __399082_399082;
   reg _399083_399083 ; 
   reg __399083_399083;
   reg _399084_399084 ; 
   reg __399084_399084;
   reg _399085_399085 ; 
   reg __399085_399085;
   reg _399086_399086 ; 
   reg __399086_399086;
   reg _399087_399087 ; 
   reg __399087_399087;
   reg _399088_399088 ; 
   reg __399088_399088;
   reg _399089_399089 ; 
   reg __399089_399089;
   reg _399090_399090 ; 
   reg __399090_399090;
   reg _399091_399091 ; 
   reg __399091_399091;
   reg _399092_399092 ; 
   reg __399092_399092;
   reg _399093_399093 ; 
   reg __399093_399093;
   reg _399094_399094 ; 
   reg __399094_399094;
   reg _399095_399095 ; 
   reg __399095_399095;
   reg _399096_399096 ; 
   reg __399096_399096;
   reg _399097_399097 ; 
   reg __399097_399097;
   reg _399098_399098 ; 
   reg __399098_399098;
   reg _399099_399099 ; 
   reg __399099_399099;
   reg _399100_399100 ; 
   reg __399100_399100;
   reg _399101_399101 ; 
   reg __399101_399101;
   reg _399102_399102 ; 
   reg __399102_399102;
   reg _399103_399103 ; 
   reg __399103_399103;
   reg _399104_399104 ; 
   reg __399104_399104;
   reg _399105_399105 ; 
   reg __399105_399105;
   reg _399106_399106 ; 
   reg __399106_399106;
   reg _399107_399107 ; 
   reg __399107_399107;
   reg _399108_399108 ; 
   reg __399108_399108;
   reg _399109_399109 ; 
   reg __399109_399109;
   reg _399110_399110 ; 
   reg __399110_399110;
   reg _399111_399111 ; 
   reg __399111_399111;
   reg _399112_399112 ; 
   reg __399112_399112;
   reg _399113_399113 ; 
   reg __399113_399113;
   reg _399114_399114 ; 
   reg __399114_399114;
   reg _399115_399115 ; 
   reg __399115_399115;
   reg _399116_399116 ; 
   reg __399116_399116;
   reg _399117_399117 ; 
   reg __399117_399117;
   reg _399118_399118 ; 
   reg __399118_399118;
   reg _399119_399119 ; 
   reg __399119_399119;
   reg _399120_399120 ; 
   reg __399120_399120;
   reg _399121_399121 ; 
   reg __399121_399121;
   reg _399122_399122 ; 
   reg __399122_399122;
   reg _399123_399123 ; 
   reg __399123_399123;
   reg _399124_399124 ; 
   reg __399124_399124;
   reg _399125_399125 ; 
   reg __399125_399125;
   reg _399126_399126 ; 
   reg __399126_399126;
   reg _399127_399127 ; 
   reg __399127_399127;
   reg _399128_399128 ; 
   reg __399128_399128;
   reg _399129_399129 ; 
   reg __399129_399129;
   reg _399130_399130 ; 
   reg __399130_399130;
   reg _399131_399131 ; 
   reg __399131_399131;
   reg _399132_399132 ; 
   reg __399132_399132;
   reg _399133_399133 ; 
   reg __399133_399133;
   reg _399134_399134 ; 
   reg __399134_399134;
   reg _399135_399135 ; 
   reg __399135_399135;
   reg _399136_399136 ; 
   reg __399136_399136;
   reg _399137_399137 ; 
   reg __399137_399137;
   reg _399138_399138 ; 
   reg __399138_399138;
   reg _399139_399139 ; 
   reg __399139_399139;
   reg _399140_399140 ; 
   reg __399140_399140;
   reg _399141_399141 ; 
   reg __399141_399141;
   reg _399142_399142 ; 
   reg __399142_399142;
   reg _399143_399143 ; 
   reg __399143_399143;
   reg _399144_399144 ; 
   reg __399144_399144;
   reg _399145_399145 ; 
   reg __399145_399145;
   reg _399146_399146 ; 
   reg __399146_399146;
   reg _399147_399147 ; 
   reg __399147_399147;
   reg _399148_399148 ; 
   reg __399148_399148;
   reg _399149_399149 ; 
   reg __399149_399149;
   reg _399150_399150 ; 
   reg __399150_399150;
   reg _399151_399151 ; 
   reg __399151_399151;
   reg _399152_399152 ; 
   reg __399152_399152;
   reg _399153_399153 ; 
   reg __399153_399153;
   reg _399154_399154 ; 
   reg __399154_399154;
   reg _399155_399155 ; 
   reg __399155_399155;
   reg _399156_399156 ; 
   reg __399156_399156;
   reg _399157_399157 ; 
   reg __399157_399157;
   reg _399158_399158 ; 
   reg __399158_399158;
   reg _399159_399159 ; 
   reg __399159_399159;
   reg _399160_399160 ; 
   reg __399160_399160;
   reg _399161_399161 ; 
   reg __399161_399161;
   reg _399162_399162 ; 
   reg __399162_399162;
   reg _399163_399163 ; 
   reg __399163_399163;
   reg _399164_399164 ; 
   reg __399164_399164;
   reg _399165_399165 ; 
   reg __399165_399165;
   reg _399166_399166 ; 
   reg __399166_399166;
   reg _399167_399167 ; 
   reg __399167_399167;
   reg _399168_399168 ; 
   reg __399168_399168;
   reg _399169_399169 ; 
   reg __399169_399169;
   reg _399170_399170 ; 
   reg __399170_399170;
   reg _399171_399171 ; 
   reg __399171_399171;
   reg _399172_399172 ; 
   reg __399172_399172;
   reg _399173_399173 ; 
   reg __399173_399173;
   reg _399174_399174 ; 
   reg __399174_399174;
   reg _399175_399175 ; 
   reg __399175_399175;
   reg _399176_399176 ; 
   reg __399176_399176;
   reg _399177_399177 ; 
   reg __399177_399177;
   reg _399178_399178 ; 
   reg __399178_399178;
   reg _399179_399179 ; 
   reg __399179_399179;
   reg _399180_399180 ; 
   reg __399180_399180;
   reg _399181_399181 ; 
   reg __399181_399181;
   reg _399182_399182 ; 
   reg __399182_399182;
   reg _399183_399183 ; 
   reg __399183_399183;
   reg _399184_399184 ; 
   reg __399184_399184;
   reg _399185_399185 ; 
   reg __399185_399185;
   reg _399186_399186 ; 
   reg __399186_399186;
   reg _399187_399187 ; 
   reg __399187_399187;
   reg _399188_399188 ; 
   reg __399188_399188;
   reg _399189_399189 ; 
   reg __399189_399189;
   reg _399190_399190 ; 
   reg __399190_399190;
   reg _399191_399191 ; 
   reg __399191_399191;
   reg _399192_399192 ; 
   reg __399192_399192;
   reg _399193_399193 ; 
   reg __399193_399193;
   reg _399194_399194 ; 
   reg __399194_399194;
   reg _399195_399195 ; 
   reg __399195_399195;
   reg _399196_399196 ; 
   reg __399196_399196;
   reg _399197_399197 ; 
   reg __399197_399197;
   reg _399198_399198 ; 
   reg __399198_399198;
   reg _399199_399199 ; 
   reg __399199_399199;
   reg _399200_399200 ; 
   reg __399200_399200;
   reg _399201_399201 ; 
   reg __399201_399201;
   reg _399202_399202 ; 
   reg __399202_399202;
   reg _399203_399203 ; 
   reg __399203_399203;
   reg _399204_399204 ; 
   reg __399204_399204;
   reg _399205_399205 ; 
   reg __399205_399205;
   reg _399206_399206 ; 
   reg __399206_399206;
   reg _399207_399207 ; 
   reg __399207_399207;
   reg _399208_399208 ; 
   reg __399208_399208;
   reg _399209_399209 ; 
   reg __399209_399209;
   reg _399210_399210 ; 
   reg __399210_399210;
   reg _399211_399211 ; 
   reg __399211_399211;
   reg _399212_399212 ; 
   reg __399212_399212;
   reg _399213_399213 ; 
   reg __399213_399213;
   reg _399214_399214 ; 
   reg __399214_399214;
   reg _399215_399215 ; 
   reg __399215_399215;
   reg _399216_399216 ; 
   reg __399216_399216;
   reg _399217_399217 ; 
   reg __399217_399217;
   reg _399218_399218 ; 
   reg __399218_399218;
   reg _399219_399219 ; 
   reg __399219_399219;
   reg _399220_399220 ; 
   reg __399220_399220;
   reg _399221_399221 ; 
   reg __399221_399221;
   reg _399222_399222 ; 
   reg __399222_399222;
   reg _399223_399223 ; 
   reg __399223_399223;
   reg _399224_399224 ; 
   reg __399224_399224;
   reg _399225_399225 ; 
   reg __399225_399225;
   reg _399226_399226 ; 
   reg __399226_399226;
   reg _399227_399227 ; 
   reg __399227_399227;
   reg _399228_399228 ; 
   reg __399228_399228;
   reg _399229_399229 ; 
   reg __399229_399229;
   reg _399230_399230 ; 
   reg __399230_399230;
   reg _399231_399231 ; 
   reg __399231_399231;
   reg _399232_399232 ; 
   reg __399232_399232;
   reg _399233_399233 ; 
   reg __399233_399233;
   reg _399234_399234 ; 
   reg __399234_399234;
   reg _399235_399235 ; 
   reg __399235_399235;
   reg _399236_399236 ; 
   reg __399236_399236;
   reg _399237_399237 ; 
   reg __399237_399237;
   reg _399238_399238 ; 
   reg __399238_399238;
   reg _399239_399239 ; 
   reg __399239_399239;
   reg _399240_399240 ; 
   reg __399240_399240;
   reg _399241_399241 ; 
   reg __399241_399241;
   reg _399242_399242 ; 
   reg __399242_399242;
   reg _399243_399243 ; 
   reg __399243_399243;
   reg _399244_399244 ; 
   reg __399244_399244;
   reg _399245_399245 ; 
   reg __399245_399245;
   reg _399246_399246 ; 
   reg __399246_399246;
   reg _399247_399247 ; 
   reg __399247_399247;
   reg _399248_399248 ; 
   reg __399248_399248;
   reg _399249_399249 ; 
   reg __399249_399249;
   reg _399250_399250 ; 
   reg __399250_399250;
   reg _399251_399251 ; 
   reg __399251_399251;
   reg _399252_399252 ; 
   reg __399252_399252;
   reg _399253_399253 ; 
   reg __399253_399253;
   reg _399254_399254 ; 
   reg __399254_399254;
   reg _399255_399255 ; 
   reg __399255_399255;
   reg _399256_399256 ; 
   reg __399256_399256;
   reg _399257_399257 ; 
   reg __399257_399257;
   reg _399258_399258 ; 
   reg __399258_399258;
   reg _399259_399259 ; 
   reg __399259_399259;
   reg _399260_399260 ; 
   reg __399260_399260;
   reg _399261_399261 ; 
   reg __399261_399261;
   reg _399262_399262 ; 
   reg __399262_399262;
   reg _399263_399263 ; 
   reg __399263_399263;
   reg _399264_399264 ; 
   reg __399264_399264;
   reg _399265_399265 ; 
   reg __399265_399265;
   reg _399266_399266 ; 
   reg __399266_399266;
   reg _399267_399267 ; 
   reg __399267_399267;
   reg _399268_399268 ; 
   reg __399268_399268;
   reg _399269_399269 ; 
   reg __399269_399269;
   reg _399270_399270 ; 
   reg __399270_399270;
   reg _399271_399271 ; 
   reg __399271_399271;
   reg _399272_399272 ; 
   reg __399272_399272;
   reg _399273_399273 ; 
   reg __399273_399273;
   reg _399274_399274 ; 
   reg __399274_399274;
   reg _399275_399275 ; 
   reg __399275_399275;
   reg _399276_399276 ; 
   reg __399276_399276;
   reg _399277_399277 ; 
   reg __399277_399277;
   reg _399278_399278 ; 
   reg __399278_399278;
   reg _399279_399279 ; 
   reg __399279_399279;
   reg _399280_399280 ; 
   reg __399280_399280;
   reg _399281_399281 ; 
   reg __399281_399281;
   reg _399282_399282 ; 
   reg __399282_399282;
   reg _399283_399283 ; 
   reg __399283_399283;
   reg _399284_399284 ; 
   reg __399284_399284;
   reg _399285_399285 ; 
   reg __399285_399285;
   reg _399286_399286 ; 
   reg __399286_399286;
   reg _399287_399287 ; 
   reg __399287_399287;
   reg _399288_399288 ; 
   reg __399288_399288;
   reg _399289_399289 ; 
   reg __399289_399289;
   reg _399290_399290 ; 
   reg __399290_399290;
   reg _399291_399291 ; 
   reg __399291_399291;
   reg _399292_399292 ; 
   reg __399292_399292;
   reg _399293_399293 ; 
   reg __399293_399293;
   reg _399294_399294 ; 
   reg __399294_399294;
   reg _399295_399295 ; 
   reg __399295_399295;
   reg _399296_399296 ; 
   reg __399296_399296;
   reg _399297_399297 ; 
   reg __399297_399297;
   reg _399298_399298 ; 
   reg __399298_399298;
   reg _399299_399299 ; 
   reg __399299_399299;
   reg _399300_399300 ; 
   reg __399300_399300;
   reg _399301_399301 ; 
   reg __399301_399301;
   reg _399302_399302 ; 
   reg __399302_399302;
   reg _399303_399303 ; 
   reg __399303_399303;
   reg _399304_399304 ; 
   reg __399304_399304;
   reg _399305_399305 ; 
   reg __399305_399305;
   reg _399306_399306 ; 
   reg __399306_399306;
   reg _399307_399307 ; 
   reg __399307_399307;
   reg _399308_399308 ; 
   reg __399308_399308;
   reg _399309_399309 ; 
   reg __399309_399309;
   reg _399310_399310 ; 
   reg __399310_399310;
   reg _399311_399311 ; 
   reg __399311_399311;
   reg _399312_399312 ; 
   reg __399312_399312;
   reg _399313_399313 ; 
   reg __399313_399313;
   reg _399314_399314 ; 
   reg __399314_399314;
   reg _399315_399315 ; 
   reg __399315_399315;
   reg _399316_399316 ; 
   reg __399316_399316;
   reg _399317_399317 ; 
   reg __399317_399317;
   reg _399318_399318 ; 
   reg __399318_399318;
   reg _399319_399319 ; 
   reg __399319_399319;
   reg _399320_399320 ; 
   reg __399320_399320;
   reg _399321_399321 ; 
   reg __399321_399321;
   reg _399322_399322 ; 
   reg __399322_399322;
   reg _399323_399323 ; 
   reg __399323_399323;
   reg _399324_399324 ; 
   reg __399324_399324;
   reg _399325_399325 ; 
   reg __399325_399325;
   reg _399326_399326 ; 
   reg __399326_399326;
   reg _399327_399327 ; 
   reg __399327_399327;
   reg _399328_399328 ; 
   reg __399328_399328;
   reg _399329_399329 ; 
   reg __399329_399329;
   reg _399330_399330 ; 
   reg __399330_399330;
   reg _399331_399331 ; 
   reg __399331_399331;
   reg _399332_399332 ; 
   reg __399332_399332;
   reg _399333_399333 ; 
   reg __399333_399333;
   reg _399334_399334 ; 
   reg __399334_399334;
   reg _399335_399335 ; 
   reg __399335_399335;
   reg _399336_399336 ; 
   reg __399336_399336;
   reg _399337_399337 ; 
   reg __399337_399337;
   reg _399338_399338 ; 
   reg __399338_399338;
   reg _399339_399339 ; 
   reg __399339_399339;
   reg _399340_399340 ; 
   reg __399340_399340;
   reg _399341_399341 ; 
   reg __399341_399341;
   reg _399342_399342 ; 
   reg __399342_399342;
   reg _399343_399343 ; 
   reg __399343_399343;
   reg _399344_399344 ; 
   reg __399344_399344;
   reg _399345_399345 ; 
   reg __399345_399345;
   reg _399346_399346 ; 
   reg __399346_399346;
   reg _399347_399347 ; 
   reg __399347_399347;
   reg _399348_399348 ; 
   reg __399348_399348;
   reg _399349_399349 ; 
   reg __399349_399349;
   reg _399350_399350 ; 
   reg __399350_399350;
   reg _399351_399351 ; 
   reg __399351_399351;
   reg _399352_399352 ; 
   reg __399352_399352;
   reg _399353_399353 ; 
   reg __399353_399353;
   reg _399354_399354 ; 
   reg __399354_399354;
   reg _399355_399355 ; 
   reg __399355_399355;
   reg _399356_399356 ; 
   reg __399356_399356;
   reg _399357_399357 ; 
   reg __399357_399357;
   reg _399358_399358 ; 
   reg __399358_399358;
   reg _399359_399359 ; 
   reg __399359_399359;
   reg _399360_399360 ; 
   reg __399360_399360;
   reg _399361_399361 ; 
   reg __399361_399361;
   reg _399362_399362 ; 
   reg __399362_399362;
   reg _399363_399363 ; 
   reg __399363_399363;
   reg _399364_399364 ; 
   reg __399364_399364;
   reg _399365_399365 ; 
   reg __399365_399365;
   reg _399366_399366 ; 
   reg __399366_399366;
   reg _399367_399367 ; 
   reg __399367_399367;
   reg _399368_399368 ; 
   reg __399368_399368;
   reg _399369_399369 ; 
   reg __399369_399369;
   reg _399370_399370 ; 
   reg __399370_399370;
   reg _399371_399371 ; 
   reg __399371_399371;
   reg _399372_399372 ; 
   reg __399372_399372;
   reg _399373_399373 ; 
   reg __399373_399373;
   reg _399374_399374 ; 
   reg __399374_399374;
   reg _399375_399375 ; 
   reg __399375_399375;
   reg _399376_399376 ; 
   reg __399376_399376;
   reg _399377_399377 ; 
   reg __399377_399377;
   reg _399378_399378 ; 
   reg __399378_399378;
   reg _399379_399379 ; 
   reg __399379_399379;
   reg _399380_399380 ; 
   reg __399380_399380;
   reg _399381_399381 ; 
   reg __399381_399381;
   reg _399382_399382 ; 
   reg __399382_399382;
   reg _399383_399383 ; 
   reg __399383_399383;
   reg _399384_399384 ; 
   reg __399384_399384;
   reg _399385_399385 ; 
   reg __399385_399385;
   reg _399386_399386 ; 
   reg __399386_399386;
   reg _399387_399387 ; 
   reg __399387_399387;
   reg _399388_399388 ; 
   reg __399388_399388;
   reg _399389_399389 ; 
   reg __399389_399389;
   reg _399390_399390 ; 
   reg __399390_399390;
   reg _399391_399391 ; 
   reg __399391_399391;
   reg _399392_399392 ; 
   reg __399392_399392;
   reg _399393_399393 ; 
   reg __399393_399393;
   reg _399394_399394 ; 
   reg __399394_399394;
   reg _399395_399395 ; 
   reg __399395_399395;
   reg _399396_399396 ; 
   reg __399396_399396;
   reg _399397_399397 ; 
   reg __399397_399397;
   reg _399398_399398 ; 
   reg __399398_399398;
   reg _399399_399399 ; 
   reg __399399_399399;
   reg _399400_399400 ; 
   reg __399400_399400;
   reg _399401_399401 ; 
   reg __399401_399401;
   reg _399402_399402 ; 
   reg __399402_399402;
   reg _399403_399403 ; 
   reg __399403_399403;
   reg _399404_399404 ; 
   reg __399404_399404;
   reg _399405_399405 ; 
   reg __399405_399405;
   reg _399406_399406 ; 
   reg __399406_399406;
   reg _399407_399407 ; 
   reg __399407_399407;
   reg _399408_399408 ; 
   reg __399408_399408;
   reg _399409_399409 ; 
   reg __399409_399409;
   reg _399410_399410 ; 
   reg __399410_399410;
   reg _399411_399411 ; 
   reg __399411_399411;
   reg _399412_399412 ; 
   reg __399412_399412;
   reg _399413_399413 ; 
   reg __399413_399413;
   reg _399414_399414 ; 
   reg __399414_399414;
   reg _399415_399415 ; 
   reg __399415_399415;
   reg _399416_399416 ; 
   reg __399416_399416;
   reg _399417_399417 ; 
   reg __399417_399417;
   reg _399418_399418 ; 
   reg __399418_399418;
   reg _399419_399419 ; 
   reg __399419_399419;
   reg _399420_399420 ; 
   reg __399420_399420;
   reg _399421_399421 ; 
   reg __399421_399421;
   reg _399422_399422 ; 
   reg __399422_399422;
   reg _399423_399423 ; 
   reg __399423_399423;
   reg _399424_399424 ; 
   reg __399424_399424;
   reg _399425_399425 ; 
   reg __399425_399425;
   reg _399426_399426 ; 
   reg __399426_399426;
   reg _399427_399427 ; 
   reg __399427_399427;
   reg _399428_399428 ; 
   reg __399428_399428;
   reg _399429_399429 ; 
   reg __399429_399429;
   reg _399430_399430 ; 
   reg __399430_399430;
   reg _399431_399431 ; 
   reg __399431_399431;
   reg _399432_399432 ; 
   reg __399432_399432;
   reg _399433_399433 ; 
   reg __399433_399433;
   reg _399434_399434 ; 
   reg __399434_399434;
   reg _399435_399435 ; 
   reg __399435_399435;
   reg _399436_399436 ; 
   reg __399436_399436;
   reg _399437_399437 ; 
   reg __399437_399437;
   reg _399438_399438 ; 
   reg __399438_399438;
   reg _399439_399439 ; 
   reg __399439_399439;
   reg _399440_399440 ; 
   reg __399440_399440;
   reg _399441_399441 ; 
   reg __399441_399441;
   reg _399442_399442 ; 
   reg __399442_399442;
   reg _399443_399443 ; 
   reg __399443_399443;
   reg _399444_399444 ; 
   reg __399444_399444;
   reg _399445_399445 ; 
   reg __399445_399445;
   reg _399446_399446 ; 
   reg __399446_399446;
   reg _399447_399447 ; 
   reg __399447_399447;
   reg _399448_399448 ; 
   reg __399448_399448;
   reg _399449_399449 ; 
   reg __399449_399449;
   reg _399450_399450 ; 
   reg __399450_399450;
   reg _399451_399451 ; 
   reg __399451_399451;
   reg _399452_399452 ; 
   reg __399452_399452;
   reg _399453_399453 ; 
   reg __399453_399453;
   reg _399454_399454 ; 
   reg __399454_399454;
   reg _399455_399455 ; 
   reg __399455_399455;
   reg _399456_399456 ; 
   reg __399456_399456;
   reg _399457_399457 ; 
   reg __399457_399457;
   reg _399458_399458 ; 
   reg __399458_399458;
   reg _399459_399459 ; 
   reg __399459_399459;
   reg _399460_399460 ; 
   reg __399460_399460;
   reg _399461_399461 ; 
   reg __399461_399461;
   reg _399462_399462 ; 
   reg __399462_399462;
   reg _399463_399463 ; 
   reg __399463_399463;
   reg _399464_399464 ; 
   reg __399464_399464;
   reg _399465_399465 ; 
   reg __399465_399465;
   reg _399466_399466 ; 
   reg __399466_399466;
   reg _399467_399467 ; 
   reg __399467_399467;
   reg _399468_399468 ; 
   reg __399468_399468;
   reg _399469_399469 ; 
   reg __399469_399469;
   reg _399470_399470 ; 
   reg __399470_399470;
   reg _399471_399471 ; 
   reg __399471_399471;
   reg _399472_399472 ; 
   reg __399472_399472;
   reg _399473_399473 ; 
   reg __399473_399473;
   reg _399474_399474 ; 
   reg __399474_399474;
   reg _399475_399475 ; 
   reg __399475_399475;
   reg _399476_399476 ; 
   reg __399476_399476;
   reg _399477_399477 ; 
   reg __399477_399477;
   reg _399478_399478 ; 
   reg __399478_399478;
   reg _399479_399479 ; 
   reg __399479_399479;
   reg _399480_399480 ; 
   reg __399480_399480;
   reg _399481_399481 ; 
   reg __399481_399481;
   reg _399482_399482 ; 
   reg __399482_399482;
   reg _399483_399483 ; 
   reg __399483_399483;
   reg _399484_399484 ; 
   reg __399484_399484;
   reg _399485_399485 ; 
   reg __399485_399485;
   reg _399486_399486 ; 
   reg __399486_399486;
   reg _399487_399487 ; 
   reg __399487_399487;
   reg _399488_399488 ; 
   reg __399488_399488;
   reg _399489_399489 ; 
   reg __399489_399489;
   reg _399490_399490 ; 
   reg __399490_399490;
   reg _399491_399491 ; 
   reg __399491_399491;
   reg _399492_399492 ; 
   reg __399492_399492;
   reg _399493_399493 ; 
   reg __399493_399493;
   reg _399494_399494 ; 
   reg __399494_399494;
   reg _399495_399495 ; 
   reg __399495_399495;
   reg _399496_399496 ; 
   reg __399496_399496;
   reg _399497_399497 ; 
   reg __399497_399497;
   reg _399498_399498 ; 
   reg __399498_399498;
   reg _399499_399499 ; 
   reg __399499_399499;
   reg _399500_399500 ; 
   reg __399500_399500;
   reg _399501_399501 ; 
   reg __399501_399501;
   reg _399502_399502 ; 
   reg __399502_399502;
   reg _399503_399503 ; 
   reg __399503_399503;
   reg _399504_399504 ; 
   reg __399504_399504;
   reg _399505_399505 ; 
   reg __399505_399505;
   reg _399506_399506 ; 
   reg __399506_399506;
   reg _399507_399507 ; 
   reg __399507_399507;
   reg _399508_399508 ; 
   reg __399508_399508;
   reg _399509_399509 ; 
   reg __399509_399509;
   reg _399510_399510 ; 
   reg __399510_399510;
   reg _399511_399511 ; 
   reg __399511_399511;
   reg _399512_399512 ; 
   reg __399512_399512;
   reg _399513_399513 ; 
   reg __399513_399513;
   reg _399514_399514 ; 
   reg __399514_399514;
   reg _399515_399515 ; 
   reg __399515_399515;
   reg _399516_399516 ; 
   reg __399516_399516;
   reg _399517_399517 ; 
   reg __399517_399517;
   reg _399518_399518 ; 
   reg __399518_399518;
   reg _399519_399519 ; 
   reg __399519_399519;
   reg _399520_399520 ; 
   reg __399520_399520;
   reg _399521_399521 ; 
   reg __399521_399521;
   reg _399522_399522 ; 
   reg __399522_399522;
   reg _399523_399523 ; 
   reg __399523_399523;
   reg _399524_399524 ; 
   reg __399524_399524;
   reg _399525_399525 ; 
   reg __399525_399525;
   reg _399526_399526 ; 
   reg __399526_399526;
   reg _399527_399527 ; 
   reg __399527_399527;
   reg _399528_399528 ; 
   reg __399528_399528;
   reg _399529_399529 ; 
   reg __399529_399529;
   reg _399530_399530 ; 
   reg __399530_399530;
   reg _399531_399531 ; 
   reg __399531_399531;
   reg _399532_399532 ; 
   reg __399532_399532;
   reg _399533_399533 ; 
   reg __399533_399533;
   reg _399534_399534 ; 
   reg __399534_399534;
   reg _399535_399535 ; 
   reg __399535_399535;
   reg _399536_399536 ; 
   reg __399536_399536;
   reg _399537_399537 ; 
   reg __399537_399537;
   reg _399538_399538 ; 
   reg __399538_399538;
   reg _399539_399539 ; 
   reg __399539_399539;
   reg _399540_399540 ; 
   reg __399540_399540;
   reg _399541_399541 ; 
   reg __399541_399541;
   reg _399542_399542 ; 
   reg __399542_399542;
   reg _399543_399543 ; 
   reg __399543_399543;
   reg _399544_399544 ; 
   reg __399544_399544;
   reg _399545_399545 ; 
   reg __399545_399545;
   reg _399546_399546 ; 
   reg __399546_399546;
   reg _399547_399547 ; 
   reg __399547_399547;
   reg _399548_399548 ; 
   reg __399548_399548;
   reg _399549_399549 ; 
   reg __399549_399549;
   reg _399550_399550 ; 
   reg __399550_399550;
   reg _399551_399551 ; 
   reg __399551_399551;
   reg _399552_399552 ; 
   reg __399552_399552;
   reg _399553_399553 ; 
   reg __399553_399553;
   reg _399554_399554 ; 
   reg __399554_399554;
   reg _399555_399555 ; 
   reg __399555_399555;
   reg _399556_399556 ; 
   reg __399556_399556;
   reg _399557_399557 ; 
   reg __399557_399557;
   reg _399558_399558 ; 
   reg __399558_399558;
   reg _399559_399559 ; 
   reg __399559_399559;
   reg _399560_399560 ; 
   reg __399560_399560;
   reg _399561_399561 ; 
   reg __399561_399561;
   reg _399562_399562 ; 
   reg __399562_399562;
   reg _399563_399563 ; 
   reg __399563_399563;
   reg _399564_399564 ; 
   reg __399564_399564;
   reg _399565_399565 ; 
   reg __399565_399565;
   reg _399566_399566 ; 
   reg __399566_399566;
   reg _399567_399567 ; 
   reg __399567_399567;
   reg _399568_399568 ; 
   reg __399568_399568;
   reg _399569_399569 ; 
   reg __399569_399569;
   reg _399570_399570 ; 
   reg __399570_399570;
   reg _399571_399571 ; 
   reg __399571_399571;
   reg _399572_399572 ; 
   reg __399572_399572;
   reg _399573_399573 ; 
   reg __399573_399573;
   reg _399574_399574 ; 
   reg __399574_399574;
   reg _399575_399575 ; 
   reg __399575_399575;
   reg _399576_399576 ; 
   reg __399576_399576;
   reg _399577_399577 ; 
   reg __399577_399577;
   reg _399578_399578 ; 
   reg __399578_399578;
   reg _399579_399579 ; 
   reg __399579_399579;
   reg _399580_399580 ; 
   reg __399580_399580;
   reg _399581_399581 ; 
   reg __399581_399581;
   reg _399582_399582 ; 
   reg __399582_399582;
   reg _399583_399583 ; 
   reg __399583_399583;
   reg _399584_399584 ; 
   reg __399584_399584;
   reg _399585_399585 ; 
   reg __399585_399585;
   reg _399586_399586 ; 
   reg __399586_399586;
   reg _399587_399587 ; 
   reg __399587_399587;
   reg _399588_399588 ; 
   reg __399588_399588;
   reg _399589_399589 ; 
   reg __399589_399589;
   reg _399590_399590 ; 
   reg __399590_399590;
   reg _399591_399591 ; 
   reg __399591_399591;
   reg _399592_399592 ; 
   reg __399592_399592;
   reg _399593_399593 ; 
   reg __399593_399593;
   reg _399594_399594 ; 
   reg __399594_399594;
   reg _399595_399595 ; 
   reg __399595_399595;
   reg _399596_399596 ; 
   reg __399596_399596;
   reg _399597_399597 ; 
   reg __399597_399597;
   reg _399598_399598 ; 
   reg __399598_399598;
   reg _399599_399599 ; 
   reg __399599_399599;
   reg _399600_399600 ; 
   reg __399600_399600;
   reg _399601_399601 ; 
   reg __399601_399601;
   reg _399602_399602 ; 
   reg __399602_399602;
   reg _399603_399603 ; 
   reg __399603_399603;
   reg _399604_399604 ; 
   reg __399604_399604;
   reg _399605_399605 ; 
   reg __399605_399605;
   reg _399606_399606 ; 
   reg __399606_399606;
   reg _399607_399607 ; 
   reg __399607_399607;
   reg _399608_399608 ; 
   reg __399608_399608;
   reg _399609_399609 ; 
   reg __399609_399609;
   reg _399610_399610 ; 
   reg __399610_399610;
   reg _399611_399611 ; 
   reg __399611_399611;
   reg _399612_399612 ; 
   reg __399612_399612;
   reg _399613_399613 ; 
   reg __399613_399613;
   reg _399614_399614 ; 
   reg __399614_399614;
   reg _399615_399615 ; 
   reg __399615_399615;
   reg _399616_399616 ; 
   reg __399616_399616;
   reg _399617_399617 ; 
   reg __399617_399617;
   reg _399618_399618 ; 
   reg __399618_399618;
   reg _399619_399619 ; 
   reg __399619_399619;
   reg _399620_399620 ; 
   reg __399620_399620;
   reg _399621_399621 ; 
   reg __399621_399621;
   reg _399622_399622 ; 
   reg __399622_399622;
   reg _399623_399623 ; 
   reg __399623_399623;
   reg _399624_399624 ; 
   reg __399624_399624;
   reg _399625_399625 ; 
   reg __399625_399625;
   reg _399626_399626 ; 
   reg __399626_399626;
   reg _399627_399627 ; 
   reg __399627_399627;
   reg _399628_399628 ; 
   reg __399628_399628;
   reg _399629_399629 ; 
   reg __399629_399629;
   reg _399630_399630 ; 
   reg __399630_399630;
   reg _399631_399631 ; 
   reg __399631_399631;
   reg _399632_399632 ; 
   reg __399632_399632;
   reg _399633_399633 ; 
   reg __399633_399633;
   reg _399634_399634 ; 
   reg __399634_399634;
   reg _399635_399635 ; 
   reg __399635_399635;
   reg _399636_399636 ; 
   reg __399636_399636;
   reg _399637_399637 ; 
   reg __399637_399637;
   reg _399638_399638 ; 
   reg __399638_399638;
   reg _399639_399639 ; 
   reg __399639_399639;
   reg _399640_399640 ; 
   reg __399640_399640;
   reg _399641_399641 ; 
   reg __399641_399641;
   reg _399642_399642 ; 
   reg __399642_399642;
   reg _399643_399643 ; 
   reg __399643_399643;
   reg _399644_399644 ; 
   reg __399644_399644;
   reg _399645_399645 ; 
   reg __399645_399645;
   reg _399646_399646 ; 
   reg __399646_399646;
   reg _399647_399647 ; 
   reg __399647_399647;
   reg _399648_399648 ; 
   reg __399648_399648;
   reg _399649_399649 ; 
   reg __399649_399649;
   reg _399650_399650 ; 
   reg __399650_399650;
   reg _399651_399651 ; 
   reg __399651_399651;
   reg _399652_399652 ; 
   reg __399652_399652;
   reg _399653_399653 ; 
   reg __399653_399653;
   reg _399654_399654 ; 
   reg __399654_399654;
   reg _399655_399655 ; 
   reg __399655_399655;
   reg _399656_399656 ; 
   reg __399656_399656;
   reg _399657_399657 ; 
   reg __399657_399657;
   reg _399658_399658 ; 
   reg __399658_399658;
   reg _399659_399659 ; 
   reg __399659_399659;
   reg _399660_399660 ; 
   reg __399660_399660;
   reg _399661_399661 ; 
   reg __399661_399661;
   reg _399662_399662 ; 
   reg __399662_399662;
   reg _399663_399663 ; 
   reg __399663_399663;
   reg _399664_399664 ; 
   reg __399664_399664;
   reg _399665_399665 ; 
   reg __399665_399665;
   reg _399666_399666 ; 
   reg __399666_399666;
   reg _399667_399667 ; 
   reg __399667_399667;
   reg _399668_399668 ; 
   reg __399668_399668;
   reg _399669_399669 ; 
   reg __399669_399669;
   reg _399670_399670 ; 
   reg __399670_399670;
   reg _399671_399671 ; 
   reg __399671_399671;
   reg _399672_399672 ; 
   reg __399672_399672;
   reg _399673_399673 ; 
   reg __399673_399673;
   reg _399674_399674 ; 
   reg __399674_399674;
   reg _399675_399675 ; 
   reg __399675_399675;
   reg _399676_399676 ; 
   reg __399676_399676;
   reg _399677_399677 ; 
   reg __399677_399677;
   reg _399678_399678 ; 
   reg __399678_399678;
   reg _399679_399679 ; 
   reg __399679_399679;
   reg _399680_399680 ; 
   reg __399680_399680;
   reg _399681_399681 ; 
   reg __399681_399681;
   reg _399682_399682 ; 
   reg __399682_399682;
   reg _399683_399683 ; 
   reg __399683_399683;
   reg _399684_399684 ; 
   reg __399684_399684;
   reg _399685_399685 ; 
   reg __399685_399685;
   reg _399686_399686 ; 
   reg __399686_399686;
   reg _399687_399687 ; 
   reg __399687_399687;
   reg _399688_399688 ; 
   reg __399688_399688;
   reg _399689_399689 ; 
   reg __399689_399689;
   reg _399690_399690 ; 
   reg __399690_399690;
   reg _399691_399691 ; 
   reg __399691_399691;
   reg _399692_399692 ; 
   reg __399692_399692;
   reg _399693_399693 ; 
   reg __399693_399693;
   reg _399694_399694 ; 
   reg __399694_399694;
   reg _399695_399695 ; 
   reg __399695_399695;
   reg _399696_399696 ; 
   reg __399696_399696;
   reg _399697_399697 ; 
   reg __399697_399697;
   reg _399698_399698 ; 
   reg __399698_399698;
   reg _399699_399699 ; 
   reg __399699_399699;
   reg _399700_399700 ; 
   reg __399700_399700;
   reg _399701_399701 ; 
   reg __399701_399701;
   reg _399702_399702 ; 
   reg __399702_399702;
   reg _399703_399703 ; 
   reg __399703_399703;
   reg _399704_399704 ; 
   reg __399704_399704;
   reg _399705_399705 ; 
   reg __399705_399705;
   reg _399706_399706 ; 
   reg __399706_399706;
   reg _399707_399707 ; 
   reg __399707_399707;
   reg _399708_399708 ; 
   reg __399708_399708;
   reg _399709_399709 ; 
   reg __399709_399709;
   reg _399710_399710 ; 
   reg __399710_399710;
   reg _399711_399711 ; 
   reg __399711_399711;
   reg _399712_399712 ; 
   reg __399712_399712;
   reg _399713_399713 ; 
   reg __399713_399713;
   reg _399714_399714 ; 
   reg __399714_399714;
   reg _399715_399715 ; 
   reg __399715_399715;
   reg _399716_399716 ; 
   reg __399716_399716;
   reg _399717_399717 ; 
   reg __399717_399717;
   reg _399718_399718 ; 
   reg __399718_399718;
   reg _399719_399719 ; 
   reg __399719_399719;
   reg _399720_399720 ; 
   reg __399720_399720;
   reg _399721_399721 ; 
   reg __399721_399721;
   reg _399722_399722 ; 
   reg __399722_399722;
   reg _399723_399723 ; 
   reg __399723_399723;
   reg _399724_399724 ; 
   reg __399724_399724;
   reg _399725_399725 ; 
   reg __399725_399725;
   reg _399726_399726 ; 
   reg __399726_399726;
   reg _399727_399727 ; 
   reg __399727_399727;
   reg _399728_399728 ; 
   reg __399728_399728;
   reg _399729_399729 ; 
   reg __399729_399729;
   reg _399730_399730 ; 
   reg __399730_399730;
   reg _399731_399731 ; 
   reg __399731_399731;
   reg _399732_399732 ; 
   reg __399732_399732;
   reg _399733_399733 ; 
   reg __399733_399733;
   reg _399734_399734 ; 
   reg __399734_399734;
   reg _399735_399735 ; 
   reg __399735_399735;
   reg _399736_399736 ; 
   reg __399736_399736;
   reg _399737_399737 ; 
   reg __399737_399737;
   reg _399738_399738 ; 
   reg __399738_399738;
   reg _399739_399739 ; 
   reg __399739_399739;
   reg _399740_399740 ; 
   reg __399740_399740;
   reg _399741_399741 ; 
   reg __399741_399741;
   reg _399742_399742 ; 
   reg __399742_399742;
   reg _399743_399743 ; 
   reg __399743_399743;
   reg _399744_399744 ; 
   reg __399744_399744;
   reg _399745_399745 ; 
   reg __399745_399745;
   reg _399746_399746 ; 
   reg __399746_399746;
   reg _399747_399747 ; 
   reg __399747_399747;
   reg _399748_399748 ; 
   reg __399748_399748;
   reg _399749_399749 ; 
   reg __399749_399749;
   reg _399750_399750 ; 
   reg __399750_399750;
   reg _399751_399751 ; 
   reg __399751_399751;
   reg _399752_399752 ; 
   reg __399752_399752;
   reg _399753_399753 ; 
   reg __399753_399753;
   reg _399754_399754 ; 
   reg __399754_399754;
   reg _399755_399755 ; 
   reg __399755_399755;
   reg _399756_399756 ; 
   reg __399756_399756;
   reg _399757_399757 ; 
   reg __399757_399757;
   reg _399758_399758 ; 
   reg __399758_399758;
   reg _399759_399759 ; 
   reg __399759_399759;
   reg _399760_399760 ; 
   reg __399760_399760;
   reg _399761_399761 ; 
   reg __399761_399761;
   reg _399762_399762 ; 
   reg __399762_399762;
   reg _399763_399763 ; 
   reg __399763_399763;
   reg _399764_399764 ; 
   reg __399764_399764;
   reg _399765_399765 ; 
   reg __399765_399765;
   reg _399766_399766 ; 
   reg __399766_399766;
   reg _399767_399767 ; 
   reg __399767_399767;
   reg _399768_399768 ; 
   reg __399768_399768;
   reg _399769_399769 ; 
   reg __399769_399769;
   reg _399770_399770 ; 
   reg __399770_399770;
   reg _399771_399771 ; 
   reg __399771_399771;
   reg _399772_399772 ; 
   reg __399772_399772;
   reg _399773_399773 ; 
   reg __399773_399773;
   reg _399774_399774 ; 
   reg __399774_399774;
   reg _399775_399775 ; 
   reg __399775_399775;
   reg _399776_399776 ; 
   reg __399776_399776;
   reg _399777_399777 ; 
   reg __399777_399777;
   reg _399778_399778 ; 
   reg __399778_399778;
   reg _399779_399779 ; 
   reg __399779_399779;
   reg _399780_399780 ; 
   reg __399780_399780;
   reg _399781_399781 ; 
   reg __399781_399781;
   reg _399782_399782 ; 
   reg __399782_399782;
   reg _399783_399783 ; 
   reg __399783_399783;
   reg _399784_399784 ; 
   reg __399784_399784;
   reg _399785_399785 ; 
   reg __399785_399785;
   reg _399786_399786 ; 
   reg __399786_399786;
   reg _399787_399787 ; 
   reg __399787_399787;
   reg _399788_399788 ; 
   reg __399788_399788;
   reg _399789_399789 ; 
   reg __399789_399789;
   reg _399790_399790 ; 
   reg __399790_399790;
   reg _399791_399791 ; 
   reg __399791_399791;
   reg _399792_399792 ; 
   reg __399792_399792;
   reg _399793_399793 ; 
   reg __399793_399793;
   reg _399794_399794 ; 
   reg __399794_399794;
   reg _399795_399795 ; 
   reg __399795_399795;
   reg _399796_399796 ; 
   reg __399796_399796;
   reg _399797_399797 ; 
   reg __399797_399797;
   reg _399798_399798 ; 
   reg __399798_399798;
   reg _399799_399799 ; 
   reg __399799_399799;
   reg _399800_399800 ; 
   reg __399800_399800;
   reg _399801_399801 ; 
   reg __399801_399801;
   reg _399802_399802 ; 
   reg __399802_399802;
   reg _399803_399803 ; 
   reg __399803_399803;
   reg _399804_399804 ; 
   reg __399804_399804;
   reg _399805_399805 ; 
   reg __399805_399805;
   reg _399806_399806 ; 
   reg __399806_399806;
   reg _399807_399807 ; 
   reg __399807_399807;
   reg _399808_399808 ; 
   reg __399808_399808;
   reg _399809_399809 ; 
   reg __399809_399809;
   reg _399810_399810 ; 
   reg __399810_399810;
   reg _399811_399811 ; 
   reg __399811_399811;
   reg _399812_399812 ; 
   reg __399812_399812;
   reg _399813_399813 ; 
   reg __399813_399813;
   reg _399814_399814 ; 
   reg __399814_399814;
   reg _399815_399815 ; 
   reg __399815_399815;
   reg _399816_399816 ; 
   reg __399816_399816;
   reg _399817_399817 ; 
   reg __399817_399817;
   reg _399818_399818 ; 
   reg __399818_399818;
   reg _399819_399819 ; 
   reg __399819_399819;
   reg _399820_399820 ; 
   reg __399820_399820;
   reg _399821_399821 ; 
   reg __399821_399821;
   reg _399822_399822 ; 
   reg __399822_399822;
   reg _399823_399823 ; 
   reg __399823_399823;
   reg _399824_399824 ; 
   reg __399824_399824;
   reg _399825_399825 ; 
   reg __399825_399825;
   reg _399826_399826 ; 
   reg __399826_399826;
   reg _399827_399827 ; 
   reg __399827_399827;
   reg _399828_399828 ; 
   reg __399828_399828;
   reg _399829_399829 ; 
   reg __399829_399829;
   reg _399830_399830 ; 
   reg __399830_399830;
   reg _399831_399831 ; 
   reg __399831_399831;
   reg _399832_399832 ; 
   reg __399832_399832;
   reg _399833_399833 ; 
   reg __399833_399833;
   reg _399834_399834 ; 
   reg __399834_399834;
   reg _399835_399835 ; 
   reg __399835_399835;
   reg _399836_399836 ; 
   reg __399836_399836;
   reg _399837_399837 ; 
   reg __399837_399837;
   reg _399838_399838 ; 
   reg __399838_399838;
   reg _399839_399839 ; 
   reg __399839_399839;
   reg _399840_399840 ; 
   reg __399840_399840;
   reg _399841_399841 ; 
   reg __399841_399841;
   reg _399842_399842 ; 
   reg __399842_399842;
   reg _399843_399843 ; 
   reg __399843_399843;
   reg _399844_399844 ; 
   reg __399844_399844;
   reg _399845_399845 ; 
   reg __399845_399845;
   reg _399846_399846 ; 
   reg __399846_399846;
   reg _399847_399847 ; 
   reg __399847_399847;
   reg _399848_399848 ; 
   reg __399848_399848;
   reg _399849_399849 ; 
   reg __399849_399849;
   reg _399850_399850 ; 
   reg __399850_399850;
   reg _399851_399851 ; 
   reg __399851_399851;
   reg _399852_399852 ; 
   reg __399852_399852;
   reg _399853_399853 ; 
   reg __399853_399853;
   reg _399854_399854 ; 
   reg __399854_399854;
   reg _399855_399855 ; 
   reg __399855_399855;
   reg _399856_399856 ; 
   reg __399856_399856;
   reg _399857_399857 ; 
   reg __399857_399857;
   reg _399858_399858 ; 
   reg __399858_399858;
   reg _399859_399859 ; 
   reg __399859_399859;
   reg _399860_399860 ; 
   reg __399860_399860;
   reg _399861_399861 ; 
   reg __399861_399861;
   reg _399862_399862 ; 
   reg __399862_399862;
   reg _399863_399863 ; 
   reg __399863_399863;
   reg _399864_399864 ; 
   reg __399864_399864;
   reg _399865_399865 ; 
   reg __399865_399865;
   reg _399866_399866 ; 
   reg __399866_399866;
   reg _399867_399867 ; 
   reg __399867_399867;
   reg _399868_399868 ; 
   reg __399868_399868;
   reg _399869_399869 ; 
   reg __399869_399869;
   reg _399870_399870 ; 
   reg __399870_399870;
   reg _399871_399871 ; 
   reg __399871_399871;
   reg _399872_399872 ; 
   reg __399872_399872;
   reg _399873_399873 ; 
   reg __399873_399873;
   reg _399874_399874 ; 
   reg __399874_399874;
   reg _399875_399875 ; 
   reg __399875_399875;
   reg _399876_399876 ; 
   reg __399876_399876;
   reg _399877_399877 ; 
   reg __399877_399877;
   reg _399878_399878 ; 
   reg __399878_399878;
   reg _399879_399879 ; 
   reg __399879_399879;
   reg _399880_399880 ; 
   reg __399880_399880;
   reg _399881_399881 ; 
   reg __399881_399881;
   reg _399882_399882 ; 
   reg __399882_399882;
   reg _399883_399883 ; 
   reg __399883_399883;
   reg _399884_399884 ; 
   reg __399884_399884;
   reg _399885_399885 ; 
   reg __399885_399885;
   reg _399886_399886 ; 
   reg __399886_399886;
   reg _399887_399887 ; 
   reg __399887_399887;
   reg _399888_399888 ; 
   reg __399888_399888;
   reg _399889_399889 ; 
   reg __399889_399889;
   reg _399890_399890 ; 
   reg __399890_399890;
   reg _399891_399891 ; 
   reg __399891_399891;
   reg _399892_399892 ; 
   reg __399892_399892;
   reg _399893_399893 ; 
   reg __399893_399893;
   reg _399894_399894 ; 
   reg __399894_399894;
   reg _399895_399895 ; 
   reg __399895_399895;
   reg _399896_399896 ; 
   reg __399896_399896;
   reg _399897_399897 ; 
   reg __399897_399897;
   reg _399898_399898 ; 
   reg __399898_399898;
   reg _399899_399899 ; 
   reg __399899_399899;
   reg _399900_399900 ; 
   reg __399900_399900;
   reg _399901_399901 ; 
   reg __399901_399901;
   reg _399902_399902 ; 
   reg __399902_399902;
   reg _399903_399903 ; 
   reg __399903_399903;
   reg _399904_399904 ; 
   reg __399904_399904;
   reg _399905_399905 ; 
   reg __399905_399905;
   reg _399906_399906 ; 
   reg __399906_399906;
   reg _399907_399907 ; 
   reg __399907_399907;
   reg _399908_399908 ; 
   reg __399908_399908;
   reg _399909_399909 ; 
   reg __399909_399909;
   reg _399910_399910 ; 
   reg __399910_399910;
   reg _399911_399911 ; 
   reg __399911_399911;
   reg _399912_399912 ; 
   reg __399912_399912;
   reg _399913_399913 ; 
   reg __399913_399913;
   reg _399914_399914 ; 
   reg __399914_399914;
   reg _399915_399915 ; 
   reg __399915_399915;
   reg _399916_399916 ; 
   reg __399916_399916;
   reg _399917_399917 ; 
   reg __399917_399917;
   reg _399918_399918 ; 
   reg __399918_399918;
   reg _399919_399919 ; 
   reg __399919_399919;
   reg _399920_399920 ; 
   reg __399920_399920;
   reg _399921_399921 ; 
   reg __399921_399921;
   reg _399922_399922 ; 
   reg __399922_399922;
   reg _399923_399923 ; 
   reg __399923_399923;
   reg _399924_399924 ; 
   reg __399924_399924;
   reg _399925_399925 ; 
   reg __399925_399925;
   reg _399926_399926 ; 
   reg __399926_399926;
   reg _399927_399927 ; 
   reg __399927_399927;
   reg _399928_399928 ; 
   reg __399928_399928;
   reg _399929_399929 ; 
   reg __399929_399929;
   reg _399930_399930 ; 
   reg __399930_399930;
   reg _399931_399931 ; 
   reg __399931_399931;
   reg _399932_399932 ; 
   reg __399932_399932;
   reg _399933_399933 ; 
   reg __399933_399933;
   reg _399934_399934 ; 
   reg __399934_399934;
   reg _399935_399935 ; 
   reg __399935_399935;
   reg _399936_399936 ; 
   reg __399936_399936;
   reg _399937_399937 ; 
   reg __399937_399937;
   reg _399938_399938 ; 
   reg __399938_399938;
   reg _399939_399939 ; 
   reg __399939_399939;
   reg _399940_399940 ; 
   reg __399940_399940;
   reg _399941_399941 ; 
   reg __399941_399941;
   reg _399942_399942 ; 
   reg __399942_399942;
   reg _399943_399943 ; 
   reg __399943_399943;
   reg _399944_399944 ; 
   reg __399944_399944;
   reg _399945_399945 ; 
   reg __399945_399945;
   reg _399946_399946 ; 
   reg __399946_399946;
   reg _399947_399947 ; 
   reg __399947_399947;
   reg _399948_399948 ; 
   reg __399948_399948;
   reg _399949_399949 ; 
   reg __399949_399949;
   reg _399950_399950 ; 
   reg __399950_399950;
   reg _399951_399951 ; 
   reg __399951_399951;
   reg _399952_399952 ; 
   reg __399952_399952;
   reg _399953_399953 ; 
   reg __399953_399953;
   reg _399954_399954 ; 
   reg __399954_399954;
   reg _399955_399955 ; 
   reg __399955_399955;
   reg _399956_399956 ; 
   reg __399956_399956;
   reg _399957_399957 ; 
   reg __399957_399957;
   reg _399958_399958 ; 
   reg __399958_399958;
   reg _399959_399959 ; 
   reg __399959_399959;
   reg _399960_399960 ; 
   reg __399960_399960;
   reg _399961_399961 ; 
   reg __399961_399961;
   reg _399962_399962 ; 
   reg __399962_399962;
   reg _399963_399963 ; 
   reg __399963_399963;
   reg _399964_399964 ; 
   reg __399964_399964;
   reg _399965_399965 ; 
   reg __399965_399965;
   reg _399966_399966 ; 
   reg __399966_399966;
   reg _399967_399967 ; 
   reg __399967_399967;
   reg _399968_399968 ; 
   reg __399968_399968;
   reg _399969_399969 ; 
   reg __399969_399969;
   reg _399970_399970 ; 
   reg __399970_399970;
   reg _399971_399971 ; 
   reg __399971_399971;
   reg _399972_399972 ; 
   reg __399972_399972;
   reg _399973_399973 ; 
   reg __399973_399973;
   reg _399974_399974 ; 
   reg __399974_399974;
   reg _399975_399975 ; 
   reg __399975_399975;
   reg _399976_399976 ; 
   reg __399976_399976;
   reg _399977_399977 ; 
   reg __399977_399977;
   reg _399978_399978 ; 
   reg __399978_399978;
   reg _399979_399979 ; 
   reg __399979_399979;
   reg _399980_399980 ; 
   reg __399980_399980;
   reg _399981_399981 ; 
   reg __399981_399981;
   reg _399982_399982 ; 
   reg __399982_399982;
   reg _399983_399983 ; 
   reg __399983_399983;
   reg _399984_399984 ; 
   reg __399984_399984;
   reg _399985_399985 ; 
   reg __399985_399985;
   reg _399986_399986 ; 
   reg __399986_399986;
   reg _399987_399987 ; 
   reg __399987_399987;
   reg _399988_399988 ; 
   reg __399988_399988;
   reg _399989_399989 ; 
   reg __399989_399989;
   reg _399990_399990 ; 
   reg __399990_399990;
   reg _399991_399991 ; 
   reg __399991_399991;
   reg _399992_399992 ; 
   reg __399992_399992;
   reg _399993_399993 ; 
   reg __399993_399993;
   reg _399994_399994 ; 
   reg __399994_399994;
   reg _399995_399995 ; 
   reg __399995_399995;
   reg _399996_399996 ; 
   reg __399996_399996;
   reg _399997_399997 ; 
   reg __399997_399997;
   reg _399998_399998 ; 
   reg __399998_399998;
   reg _399999_399999 ; 
   reg __399999_399999;
   reg _400000_400000 ; 
   reg __400000_400000;
   reg _400001_400001 ; 
   reg __400001_400001;
   reg _400002_400002 ; 
   reg __400002_400002;
   reg _400003_400003 ; 
   reg __400003_400003;
   reg _400004_400004 ; 
   reg __400004_400004;
   reg _400005_400005 ; 
   reg __400005_400005;
   reg _400006_400006 ; 
   reg __400006_400006;
   reg _400007_400007 ; 
   reg __400007_400007;
   reg _400008_400008 ; 
   reg __400008_400008;
   reg _400009_400009 ; 
   reg __400009_400009;
   reg _400010_400010 ; 
   reg __400010_400010;
   reg _400011_400011 ; 
   reg __400011_400011;
   reg _400012_400012 ; 
   reg __400012_400012;
   reg _400013_400013 ; 
   reg __400013_400013;
   reg _400014_400014 ; 
   reg __400014_400014;
   reg _400015_400015 ; 
   reg __400015_400015;
   reg _400016_400016 ; 
   reg __400016_400016;
   reg _400017_400017 ; 
   reg __400017_400017;
   reg _400018_400018 ; 
   reg __400018_400018;
   reg _400019_400019 ; 
   reg __400019_400019;
   reg _400020_400020 ; 
   reg __400020_400020;
   reg _400021_400021 ; 
   reg __400021_400021;
   reg _400022_400022 ; 
   reg __400022_400022;
   reg _400023_400023 ; 
   reg __400023_400023;
   reg _400024_400024 ; 
   reg __400024_400024;
   reg _400025_400025 ; 
   reg __400025_400025;
   reg _400026_400026 ; 
   reg __400026_400026;
   reg _400027_400027 ; 
   reg __400027_400027;
   reg _400028_400028 ; 
   reg __400028_400028;
   reg _400029_400029 ; 
   reg __400029_400029;
   reg _400030_400030 ; 
   reg __400030_400030;
   reg _400031_400031 ; 
   reg __400031_400031;
   reg _400032_400032 ; 
   reg __400032_400032;
   reg _400033_400033 ; 
   reg __400033_400033;
   reg _400034_400034 ; 
   reg __400034_400034;
   reg _400035_400035 ; 
   reg __400035_400035;
   reg _400036_400036 ; 
   reg __400036_400036;
   reg _400037_400037 ; 
   reg __400037_400037;
   reg _400038_400038 ; 
   reg __400038_400038;
   reg _400039_400039 ; 
   reg __400039_400039;
   reg _400040_400040 ; 
   reg __400040_400040;
   reg _400041_400041 ; 
   reg __400041_400041;
   reg _400042_400042 ; 
   reg __400042_400042;
   reg _400043_400043 ; 
   reg __400043_400043;
   reg _400044_400044 ; 
   reg __400044_400044;
   reg _400045_400045 ; 
   reg __400045_400045;
   reg _400046_400046 ; 
   reg __400046_400046;
   reg _400047_400047 ; 
   reg __400047_400047;
   reg _400048_400048 ; 
   reg __400048_400048;
   reg _400049_400049 ; 
   reg __400049_400049;
   reg _400050_400050 ; 
   reg __400050_400050;
   reg _400051_400051 ; 
   reg __400051_400051;
   reg _400052_400052 ; 
   reg __400052_400052;
   reg _400053_400053 ; 
   reg __400053_400053;
   reg _400054_400054 ; 
   reg __400054_400054;
   reg _400055_400055 ; 
   reg __400055_400055;
   reg _400056_400056 ; 
   reg __400056_400056;
   reg _400057_400057 ; 
   reg __400057_400057;
   reg _400058_400058 ; 
   reg __400058_400058;
   reg _400059_400059 ; 
   reg __400059_400059;
   reg _400060_400060 ; 
   reg __400060_400060;
   reg _400061_400061 ; 
   reg __400061_400061;
   reg _400062_400062 ; 
   reg __400062_400062;
   reg _400063_400063 ; 
   reg __400063_400063;
   reg _400064_400064 ; 
   reg __400064_400064;
   reg _400065_400065 ; 
   reg __400065_400065;
   reg _400066_400066 ; 
   reg __400066_400066;
   reg _400067_400067 ; 
   reg __400067_400067;
   reg _400068_400068 ; 
   reg __400068_400068;
   reg _400069_400069 ; 
   reg __400069_400069;
   reg _400070_400070 ; 
   reg __400070_400070;
   reg _400071_400071 ; 
   reg __400071_400071;
   reg _400072_400072 ; 
   reg __400072_400072;
   reg _400073_400073 ; 
   reg __400073_400073;
   reg _400074_400074 ; 
   reg __400074_400074;
   reg _400075_400075 ; 
   reg __400075_400075;
   reg _400076_400076 ; 
   reg __400076_400076;
   reg _400077_400077 ; 
   reg __400077_400077;
   reg _400078_400078 ; 
   reg __400078_400078;
   reg _400079_400079 ; 
   reg __400079_400079;
   reg _400080_400080 ; 
   reg __400080_400080;
   reg _400081_400081 ; 
   reg __400081_400081;
   reg _400082_400082 ; 
   reg __400082_400082;
   reg _400083_400083 ; 
   reg __400083_400083;
   reg _400084_400084 ; 
   reg __400084_400084;
   reg _400085_400085 ; 
   reg __400085_400085;
   reg _400086_400086 ; 
   reg __400086_400086;
   reg _400087_400087 ; 
   reg __400087_400087;
   reg _400088_400088 ; 
   reg __400088_400088;
   reg _400089_400089 ; 
   reg __400089_400089;
   reg _400090_400090 ; 
   reg __400090_400090;
   reg _400091_400091 ; 
   reg __400091_400091;
   reg _400092_400092 ; 
   reg __400092_400092;
   reg _400093_400093 ; 
   reg __400093_400093;
   reg _400094_400094 ; 
   reg __400094_400094;
   reg _400095_400095 ; 
   reg __400095_400095;
   reg _400096_400096 ; 
   reg __400096_400096;
   reg _400097_400097 ; 
   reg __400097_400097;
   reg _400098_400098 ; 
   reg __400098_400098;
   reg _400099_400099 ; 
   reg __400099_400099;
   reg _400100_400100 ; 
   reg __400100_400100;
   reg _400101_400101 ; 
   reg __400101_400101;
   reg _400102_400102 ; 
   reg __400102_400102;
   reg _400103_400103 ; 
   reg __400103_400103;
   reg _400104_400104 ; 
   reg __400104_400104;
   reg _400105_400105 ; 
   reg __400105_400105;
   reg _400106_400106 ; 
   reg __400106_400106;
   reg _400107_400107 ; 
   reg __400107_400107;
   reg _400108_400108 ; 
   reg __400108_400108;
   reg _400109_400109 ; 
   reg __400109_400109;
   reg _400110_400110 ; 
   reg __400110_400110;
   reg _400111_400111 ; 
   reg __400111_400111;
   reg _400112_400112 ; 
   reg __400112_400112;
   reg _400113_400113 ; 
   reg __400113_400113;
   reg _400114_400114 ; 
   reg __400114_400114;
   reg _400115_400115 ; 
   reg __400115_400115;
   reg _400116_400116 ; 
   reg __400116_400116;
   reg _400117_400117 ; 
   reg __400117_400117;
   reg _400118_400118 ; 
   reg __400118_400118;
   reg _400119_400119 ; 
   reg __400119_400119;
   reg _400120_400120 ; 
   reg __400120_400120;
   reg _400121_400121 ; 
   reg __400121_400121;
   reg _400122_400122 ; 
   reg __400122_400122;
   reg _400123_400123 ; 
   reg __400123_400123;
   reg _400124_400124 ; 
   reg __400124_400124;
   reg _400125_400125 ; 
   reg __400125_400125;
   reg _400126_400126 ; 
   reg __400126_400126;
   reg _400127_400127 ; 
   reg __400127_400127;
   reg _400128_400128 ; 
   reg __400128_400128;
   reg _400129_400129 ; 
   reg __400129_400129;
   reg _400130_400130 ; 
   reg __400130_400130;
   reg _400131_400131 ; 
   reg __400131_400131;
   reg _400132_400132 ; 
   reg __400132_400132;
   reg _400133_400133 ; 
   reg __400133_400133;
   reg _400134_400134 ; 
   reg __400134_400134;
   reg _400135_400135 ; 
   reg __400135_400135;
   reg _400136_400136 ; 
   reg __400136_400136;
   reg _400137_400137 ; 
   reg __400137_400137;
   reg _400138_400138 ; 
   reg __400138_400138;
   reg _400139_400139 ; 
   reg __400139_400139;
   reg _400140_400140 ; 
   reg __400140_400140;
   reg _400141_400141 ; 
   reg __400141_400141;
   reg _400142_400142 ; 
   reg __400142_400142;
   reg _400143_400143 ; 
   reg __400143_400143;
   reg _400144_400144 ; 
   reg __400144_400144;
   reg _400145_400145 ; 
   reg __400145_400145;
   reg _400146_400146 ; 
   reg __400146_400146;
   reg _400147_400147 ; 
   reg __400147_400147;
   reg _400148_400148 ; 
   reg __400148_400148;
   reg _400149_400149 ; 
   reg __400149_400149;
   reg _400150_400150 ; 
   reg __400150_400150;
   reg _400151_400151 ; 
   reg __400151_400151;
   reg _400152_400152 ; 
   reg __400152_400152;
   reg _400153_400153 ; 
   reg __400153_400153;
   reg _400154_400154 ; 
   reg __400154_400154;
   reg _400155_400155 ; 
   reg __400155_400155;
   reg _400156_400156 ; 
   reg __400156_400156;
   reg _400157_400157 ; 
   reg __400157_400157;
   reg _400158_400158 ; 
   reg __400158_400158;
   reg _400159_400159 ; 
   reg __400159_400159;
   reg _400160_400160 ; 
   reg __400160_400160;
   reg _400161_400161 ; 
   reg __400161_400161;
   reg _400162_400162 ; 
   reg __400162_400162;
   reg _400163_400163 ; 
   reg __400163_400163;
   reg _400164_400164 ; 
   reg __400164_400164;
   reg _400165_400165 ; 
   reg __400165_400165;
   reg _400166_400166 ; 
   reg __400166_400166;
   reg _400167_400167 ; 
   reg __400167_400167;
   reg _400168_400168 ; 
   reg __400168_400168;
   reg _400169_400169 ; 
   reg __400169_400169;
   reg _400170_400170 ; 
   reg __400170_400170;
   reg _400171_400171 ; 
   reg __400171_400171;
   reg _400172_400172 ; 
   reg __400172_400172;
   reg _400173_400173 ; 
   reg __400173_400173;
   reg _400174_400174 ; 
   reg __400174_400174;
   reg _400175_400175 ; 
   reg __400175_400175;
   reg _400176_400176 ; 
   reg __400176_400176;
   reg _400177_400177 ; 
   reg __400177_400177;
   reg _400178_400178 ; 
   reg __400178_400178;
   reg _400179_400179 ; 
   reg __400179_400179;
   reg _400180_400180 ; 
   reg __400180_400180;
   reg _400181_400181 ; 
   reg __400181_400181;
   reg _400182_400182 ; 
   reg __400182_400182;
   reg _400183_400183 ; 
   reg __400183_400183;
   reg _400184_400184 ; 
   reg __400184_400184;
   reg _400185_400185 ; 
   reg __400185_400185;
   reg _400186_400186 ; 
   reg __400186_400186;
   reg _400187_400187 ; 
   reg __400187_400187;
   reg _400188_400188 ; 
   reg __400188_400188;
   reg _400189_400189 ; 
   reg __400189_400189;
   reg _400190_400190 ; 
   reg __400190_400190;
   reg _400191_400191 ; 
   reg __400191_400191;
   reg _400192_400192 ; 
   reg __400192_400192;
   reg _400193_400193 ; 
   reg __400193_400193;
   reg _400194_400194 ; 
   reg __400194_400194;
   reg _400195_400195 ; 
   reg __400195_400195;
   reg _400196_400196 ; 
   reg __400196_400196;
   reg _400197_400197 ; 
   reg __400197_400197;
   reg _400198_400198 ; 
   reg __400198_400198;
   reg _400199_400199 ; 
   reg __400199_400199;
   reg _400200_400200 ; 
   reg __400200_400200;
   reg _400201_400201 ; 
   reg __400201_400201;
   reg _400202_400202 ; 
   reg __400202_400202;
   reg _400203_400203 ; 
   reg __400203_400203;
   reg _400204_400204 ; 
   reg __400204_400204;
   reg _400205_400205 ; 
   reg __400205_400205;
   reg _400206_400206 ; 
   reg __400206_400206;
   reg _400207_400207 ; 
   reg __400207_400207;
   reg _400208_400208 ; 
   reg __400208_400208;
   reg _400209_400209 ; 
   reg __400209_400209;
   reg _400210_400210 ; 
   reg __400210_400210;
   reg _400211_400211 ; 
   reg __400211_400211;
   reg _400212_400212 ; 
   reg __400212_400212;
   reg _400213_400213 ; 
   reg __400213_400213;
   reg _400214_400214 ; 
   reg __400214_400214;
   reg _400215_400215 ; 
   reg __400215_400215;
   reg _400216_400216 ; 
   reg __400216_400216;
   reg _400217_400217 ; 
   reg __400217_400217;
   reg _400218_400218 ; 
   reg __400218_400218;
   reg _400219_400219 ; 
   reg __400219_400219;
   reg _400220_400220 ; 
   reg __400220_400220;
   reg _400221_400221 ; 
   reg __400221_400221;
   reg _400222_400222 ; 
   reg __400222_400222;
   reg _400223_400223 ; 
   reg __400223_400223;
   reg _400224_400224 ; 
   reg __400224_400224;
   reg _400225_400225 ; 
   reg __400225_400225;
   reg _400226_400226 ; 
   reg __400226_400226;
   reg _400227_400227 ; 
   reg __400227_400227;
   reg _400228_400228 ; 
   reg __400228_400228;
   reg _400229_400229 ; 
   reg __400229_400229;
   reg _400230_400230 ; 
   reg __400230_400230;
   reg _400231_400231 ; 
   reg __400231_400231;
   reg _400232_400232 ; 
   reg __400232_400232;
   reg _400233_400233 ; 
   reg __400233_400233;
   reg _400234_400234 ; 
   reg __400234_400234;
   reg _400235_400235 ; 
   reg __400235_400235;
   reg _400236_400236 ; 
   reg __400236_400236;
   reg _400237_400237 ; 
   reg __400237_400237;
   reg _400238_400238 ; 
   reg __400238_400238;
   reg _400239_400239 ; 
   reg __400239_400239;
   reg _400240_400240 ; 
   reg __400240_400240;
   reg _400241_400241 ; 
   reg __400241_400241;
   reg _400242_400242 ; 
   reg __400242_400242;
   reg _400243_400243 ; 
   reg __400243_400243;
   reg _400244_400244 ; 
   reg __400244_400244;
   reg _400245_400245 ; 
   reg __400245_400245;
   reg _400246_400246 ; 
   reg __400246_400246;
   reg _400247_400247 ; 
   reg __400247_400247;
   reg _400248_400248 ; 
   reg __400248_400248;
   reg _400249_400249 ; 
   reg __400249_400249;
   reg _400250_400250 ; 
   reg __400250_400250;
   reg _400251_400251 ; 
   reg __400251_400251;
   reg _400252_400252 ; 
   reg __400252_400252;
   reg _400253_400253 ; 
   reg __400253_400253;
   reg _400254_400254 ; 
   reg __400254_400254;
   reg _400255_400255 ; 
   reg __400255_400255;
   reg _400256_400256 ; 
   reg __400256_400256;
   reg _400257_400257 ; 
   reg __400257_400257;
   reg _400258_400258 ; 
   reg __400258_400258;
   reg _400259_400259 ; 
   reg __400259_400259;
   reg _400260_400260 ; 
   reg __400260_400260;
   reg _400261_400261 ; 
   reg __400261_400261;
   reg _400262_400262 ; 
   reg __400262_400262;
   reg _400263_400263 ; 
   reg __400263_400263;
   reg _400264_400264 ; 
   reg __400264_400264;
   reg _400265_400265 ; 
   reg __400265_400265;
   reg _400266_400266 ; 
   reg __400266_400266;
   reg _400267_400267 ; 
   reg __400267_400267;
   reg _400268_400268 ; 
   reg __400268_400268;
   reg _400269_400269 ; 
   reg __400269_400269;
   reg _400270_400270 ; 
   reg __400270_400270;
   reg _400271_400271 ; 
   reg __400271_400271;
   reg _400272_400272 ; 
   reg __400272_400272;
   reg _400273_400273 ; 
   reg __400273_400273;
   reg _400274_400274 ; 
   reg __400274_400274;
   reg _400275_400275 ; 
   reg __400275_400275;
   reg _400276_400276 ; 
   reg __400276_400276;
   reg _400277_400277 ; 
   reg __400277_400277;
   reg _400278_400278 ; 
   reg __400278_400278;
   reg _400279_400279 ; 
   reg __400279_400279;
   reg _400280_400280 ; 
   reg __400280_400280;
   reg _400281_400281 ; 
   reg __400281_400281;
   reg _400282_400282 ; 
   reg __400282_400282;
   reg _400283_400283 ; 
   reg __400283_400283;
   reg _400284_400284 ; 
   reg __400284_400284;
   reg _400285_400285 ; 
   reg __400285_400285;
   reg _400286_400286 ; 
   reg __400286_400286;
   reg _400287_400287 ; 
   reg __400287_400287;
   reg _400288_400288 ; 
   reg __400288_400288;
   reg _400289_400289 ; 
   reg __400289_400289;
   reg _400290_400290 ; 
   reg __400290_400290;
   reg _400291_400291 ; 
   reg __400291_400291;
   reg _400292_400292 ; 
   reg __400292_400292;
   reg _400293_400293 ; 
   reg __400293_400293;
   reg _400294_400294 ; 
   reg __400294_400294;
   reg _400295_400295 ; 
   reg __400295_400295;
   reg _400296_400296 ; 
   reg __400296_400296;
   reg _400297_400297 ; 
   reg __400297_400297;
   reg _400298_400298 ; 
   reg __400298_400298;
   reg _400299_400299 ; 
   reg __400299_400299;
   reg _400300_400300 ; 
   reg __400300_400300;
   reg _400301_400301 ; 
   reg __400301_400301;
   reg _400302_400302 ; 
   reg __400302_400302;
   reg _400303_400303 ; 
   reg __400303_400303;
   reg _400304_400304 ; 
   reg __400304_400304;
   reg _400305_400305 ; 
   reg __400305_400305;
   reg _400306_400306 ; 
   reg __400306_400306;
   reg _400307_400307 ; 
   reg __400307_400307;
   reg _400308_400308 ; 
   reg __400308_400308;
   reg _400309_400309 ; 
   reg __400309_400309;
   reg _400310_400310 ; 
   reg __400310_400310;
   reg _400311_400311 ; 
   reg __400311_400311;
   reg _400312_400312 ; 
   reg __400312_400312;
   reg _400313_400313 ; 
   reg __400313_400313;
   reg _400314_400314 ; 
   reg __400314_400314;
   reg _400315_400315 ; 
   reg __400315_400315;
   reg _400316_400316 ; 
   reg __400316_400316;
   reg _400317_400317 ; 
   reg __400317_400317;
   reg _400318_400318 ; 
   reg __400318_400318;
   reg _400319_400319 ; 
   reg __400319_400319;
   reg _400320_400320 ; 
   reg __400320_400320;
   reg _400321_400321 ; 
   reg __400321_400321;
   reg _400322_400322 ; 
   reg __400322_400322;
   reg _400323_400323 ; 
   reg __400323_400323;
   reg _400324_400324 ; 
   reg __400324_400324;
   reg _400325_400325 ; 
   reg __400325_400325;
   reg _400326_400326 ; 
   reg __400326_400326;
   reg _400327_400327 ; 
   reg __400327_400327;
   reg _400328_400328 ; 
   reg __400328_400328;
   reg _400329_400329 ; 
   reg __400329_400329;
   reg _400330_400330 ; 
   reg __400330_400330;
   reg _400331_400331 ; 
   reg __400331_400331;
   reg _400332_400332 ; 
   reg __400332_400332;
   reg _400333_400333 ; 
   reg __400333_400333;
   reg _400334_400334 ; 
   reg __400334_400334;
   reg _400335_400335 ; 
   reg __400335_400335;
   reg _400336_400336 ; 
   reg __400336_400336;
   reg _400337_400337 ; 
   reg __400337_400337;
   reg _400338_400338 ; 
   reg __400338_400338;
   reg _400339_400339 ; 
   reg __400339_400339;
   reg _400340_400340 ; 
   reg __400340_400340;
   reg _400341_400341 ; 
   reg __400341_400341;
   reg _400342_400342 ; 
   reg __400342_400342;
   reg _400343_400343 ; 
   reg __400343_400343;
   reg _400344_400344 ; 
   reg __400344_400344;
   reg _400345_400345 ; 
   reg __400345_400345;
   reg _400346_400346 ; 
   reg __400346_400346;
   reg _400347_400347 ; 
   reg __400347_400347;
   reg _400348_400348 ; 
   reg __400348_400348;
   reg _400349_400349 ; 
   reg __400349_400349;
   reg _400350_400350 ; 
   reg __400350_400350;
   reg _400351_400351 ; 
   reg __400351_400351;
   reg _400352_400352 ; 
   reg __400352_400352;
   reg _400353_400353 ; 
   reg __400353_400353;
   reg _400354_400354 ; 
   reg __400354_400354;
   reg _400355_400355 ; 
   reg __400355_400355;
   reg _400356_400356 ; 
   reg __400356_400356;
   reg _400357_400357 ; 
   reg __400357_400357;
   reg _400358_400358 ; 
   reg __400358_400358;
   reg _400359_400359 ; 
   reg __400359_400359;
   reg _400360_400360 ; 
   reg __400360_400360;
   reg _400361_400361 ; 
   reg __400361_400361;
   reg _400362_400362 ; 
   reg __400362_400362;
   reg _400363_400363 ; 
   reg __400363_400363;
   reg _400364_400364 ; 
   reg __400364_400364;
   reg _400365_400365 ; 
   reg __400365_400365;
   reg _400366_400366 ; 
   reg __400366_400366;
   reg _400367_400367 ; 
   reg __400367_400367;
   reg _400368_400368 ; 
   reg __400368_400368;
   reg _400369_400369 ; 
   reg __400369_400369;
   reg _400370_400370 ; 
   reg __400370_400370;
   reg _400371_400371 ; 
   reg __400371_400371;
   reg _400372_400372 ; 
   reg __400372_400372;
   reg _400373_400373 ; 
   reg __400373_400373;
   reg _400374_400374 ; 
   reg __400374_400374;
   reg _400375_400375 ; 
   reg __400375_400375;
   reg _400376_400376 ; 
   reg __400376_400376;
   reg _400377_400377 ; 
   reg __400377_400377;
   reg _400378_400378 ; 
   reg __400378_400378;
   reg _400379_400379 ; 
   reg __400379_400379;
   reg _400380_400380 ; 
   reg __400380_400380;
   reg _400381_400381 ; 
   reg __400381_400381;
   reg _400382_400382 ; 
   reg __400382_400382;
   reg _400383_400383 ; 
   reg __400383_400383;
   reg _400384_400384 ; 
   reg __400384_400384;
   reg _400385_400385 ; 
   reg __400385_400385;
   reg _400386_400386 ; 
   reg __400386_400386;
   reg _400387_400387 ; 
   reg __400387_400387;
   reg _400388_400388 ; 
   reg __400388_400388;
   reg _400389_400389 ; 
   reg __400389_400389;
   reg _400390_400390 ; 
   reg __400390_400390;
   reg _400391_400391 ; 
   reg __400391_400391;
   reg _400392_400392 ; 
   reg __400392_400392;
   reg _400393_400393 ; 
   reg __400393_400393;
   reg _400394_400394 ; 
   reg __400394_400394;
   reg _400395_400395 ; 
   reg __400395_400395;
   reg _400396_400396 ; 
   reg __400396_400396;
   reg _400397_400397 ; 
   reg __400397_400397;
   reg _400398_400398 ; 
   reg __400398_400398;
   reg _400399_400399 ; 
   reg __400399_400399;
   reg _400400_400400 ; 
   reg __400400_400400;
   reg _400401_400401 ; 
   reg __400401_400401;
   reg _400402_400402 ; 
   reg __400402_400402;
   reg _400403_400403 ; 
   reg __400403_400403;
   reg _400404_400404 ; 
   reg __400404_400404;
   reg _400405_400405 ; 
   reg __400405_400405;
   reg _400406_400406 ; 
   reg __400406_400406;
   reg _400407_400407 ; 
   reg __400407_400407;
   reg _400408_400408 ; 
   reg __400408_400408;
   reg _400409_400409 ; 
   reg __400409_400409;
   reg _400410_400410 ; 
   reg __400410_400410;
   reg _400411_400411 ; 
   reg __400411_400411;
   reg _400412_400412 ; 
   reg __400412_400412;
   reg _400413_400413 ; 
   reg __400413_400413;
   reg _400414_400414 ; 
   reg __400414_400414;
   reg _400415_400415 ; 
   reg __400415_400415;
   reg _400416_400416 ; 
   reg __400416_400416;
   reg _400417_400417 ; 
   reg __400417_400417;
   reg _400418_400418 ; 
   reg __400418_400418;
   reg _400419_400419 ; 
   reg __400419_400419;
   reg _400420_400420 ; 
   reg __400420_400420;
   reg _400421_400421 ; 
   reg __400421_400421;
   reg _400422_400422 ; 
   reg __400422_400422;
   reg _400423_400423 ; 
   reg __400423_400423;
   reg _400424_400424 ; 
   reg __400424_400424;
   reg _400425_400425 ; 
   reg __400425_400425;
   reg _400426_400426 ; 
   reg __400426_400426;
   reg _400427_400427 ; 
   reg __400427_400427;
   reg _400428_400428 ; 
   reg __400428_400428;
   reg _400429_400429 ; 
   reg __400429_400429;
   reg _400430_400430 ; 
   reg __400430_400430;
   reg _400431_400431 ; 
   reg __400431_400431;
   reg _400432_400432 ; 
   reg __400432_400432;
   reg _400433_400433 ; 
   reg __400433_400433;
   reg _400434_400434 ; 
   reg __400434_400434;
   reg _400435_400435 ; 
   reg __400435_400435;
   reg _400436_400436 ; 
   reg __400436_400436;
   reg _400437_400437 ; 
   reg __400437_400437;
   reg _400438_400438 ; 
   reg __400438_400438;
   reg _400439_400439 ; 
   reg __400439_400439;
   reg _400440_400440 ; 
   reg __400440_400440;
   reg _400441_400441 ; 
   reg __400441_400441;
   reg _400442_400442 ; 
   reg __400442_400442;
   reg _400443_400443 ; 
   reg __400443_400443;
   reg _400444_400444 ; 
   reg __400444_400444;
   reg _400445_400445 ; 
   reg __400445_400445;
   reg _400446_400446 ; 
   reg __400446_400446;
   reg _400447_400447 ; 
   reg __400447_400447;
   reg _400448_400448 ; 
   reg __400448_400448;
   reg _400449_400449 ; 
   reg __400449_400449;
   reg _400450_400450 ; 
   reg __400450_400450;
   reg _400451_400451 ; 
   reg __400451_400451;
   reg _400452_400452 ; 
   reg __400452_400452;
   reg _400453_400453 ; 
   reg __400453_400453;
   reg _400454_400454 ; 
   reg __400454_400454;
   reg _400455_400455 ; 
   reg __400455_400455;
   reg _400456_400456 ; 
   reg __400456_400456;
   reg _400457_400457 ; 
   reg __400457_400457;
   reg _400458_400458 ; 
   reg __400458_400458;
   reg _400459_400459 ; 
   reg __400459_400459;
   reg _400460_400460 ; 
   reg __400460_400460;
   reg _400461_400461 ; 
   reg __400461_400461;
   reg _400462_400462 ; 
   reg __400462_400462;
   reg _400463_400463 ; 
   reg __400463_400463;
   reg _400464_400464 ; 
   reg __400464_400464;
   reg _400465_400465 ; 
   reg __400465_400465;
   reg _400466_400466 ; 
   reg __400466_400466;
   reg _400467_400467 ; 
   reg __400467_400467;
   reg _400468_400468 ; 
   reg __400468_400468;
   reg _400469_400469 ; 
   reg __400469_400469;
   reg _400470_400470 ; 
   reg __400470_400470;
   reg _400471_400471 ; 
   reg __400471_400471;
   reg _400472_400472 ; 
   reg __400472_400472;
   reg _400473_400473 ; 
   reg __400473_400473;
   reg _400474_400474 ; 
   reg __400474_400474;
   reg _400475_400475 ; 
   reg __400475_400475;
   reg _400476_400476 ; 
   reg __400476_400476;
   reg _400477_400477 ; 
   reg __400477_400477;
   reg _400478_400478 ; 
   reg __400478_400478;
   reg _400479_400479 ; 
   reg __400479_400479;
   reg _400480_400480 ; 
   reg __400480_400480;
   reg _400481_400481 ; 
   reg __400481_400481;
   reg _400482_400482 ; 
   reg __400482_400482;
   reg _400483_400483 ; 
   reg __400483_400483;
   reg _400484_400484 ; 
   reg __400484_400484;
   reg _400485_400485 ; 
   reg __400485_400485;
   reg _400486_400486 ; 
   reg __400486_400486;
   reg _400487_400487 ; 
   reg __400487_400487;
   reg _400488_400488 ; 
   reg __400488_400488;
   reg _400489_400489 ; 
   reg __400489_400489;
   reg _400490_400490 ; 
   reg __400490_400490;
   reg _400491_400491 ; 
   reg __400491_400491;
   reg _400492_400492 ; 
   reg __400492_400492;
   reg _400493_400493 ; 
   reg __400493_400493;
   reg _400494_400494 ; 
   reg __400494_400494;
   reg _400495_400495 ; 
   reg __400495_400495;
   reg _400496_400496 ; 
   reg __400496_400496;
   reg _400497_400497 ; 
   reg __400497_400497;
   reg _400498_400498 ; 
   reg __400498_400498;
   reg _400499_400499 ; 
   reg __400499_400499;
   reg _400500_400500 ; 
   reg __400500_400500;
   reg _400501_400501 ; 
   reg __400501_400501;
   reg _400502_400502 ; 
   reg __400502_400502;
   reg _400503_400503 ; 
   reg __400503_400503;
   reg _400504_400504 ; 
   reg __400504_400504;
   reg _400505_400505 ; 
   reg __400505_400505;
   reg _400506_400506 ; 
   reg __400506_400506;
   reg _400507_400507 ; 
   reg __400507_400507;
   reg _400508_400508 ; 
   reg __400508_400508;
   reg _400509_400509 ; 
   reg __400509_400509;
   reg _400510_400510 ; 
   reg __400510_400510;
   reg _400511_400511 ; 
   reg __400511_400511;
   reg _400512_400512 ; 
   reg __400512_400512;
   reg _400513_400513 ; 
   reg __400513_400513;
   reg _400514_400514 ; 
   reg __400514_400514;
   reg _400515_400515 ; 
   reg __400515_400515;
   reg _400516_400516 ; 
   reg __400516_400516;
   reg _400517_400517 ; 
   reg __400517_400517;
   reg _400518_400518 ; 
   reg __400518_400518;
   reg _400519_400519 ; 
   reg __400519_400519;
   reg _400520_400520 ; 
   reg __400520_400520;
   reg _400521_400521 ; 
   reg __400521_400521;
   reg _400522_400522 ; 
   reg __400522_400522;
   reg _400523_400523 ; 
   reg __400523_400523;
   reg _400524_400524 ; 
   reg __400524_400524;
   reg _400525_400525 ; 
   reg __400525_400525;
   reg _400526_400526 ; 
   reg __400526_400526;
   reg _400527_400527 ; 
   reg __400527_400527;
   reg _400528_400528 ; 
   reg __400528_400528;
   reg _400529_400529 ; 
   reg __400529_400529;
   reg _400530_400530 ; 
   reg __400530_400530;
   reg _400531_400531 ; 
   reg __400531_400531;
   reg _400532_400532 ; 
   reg __400532_400532;
   reg _400533_400533 ; 
   reg __400533_400533;
   reg _400534_400534 ; 
   reg __400534_400534;
   reg _400535_400535 ; 
   reg __400535_400535;
   reg _400536_400536 ; 
   reg __400536_400536;
   reg _400537_400537 ; 
   reg __400537_400537;
   reg _400538_400538 ; 
   reg __400538_400538;
   reg _400539_400539 ; 
   reg __400539_400539;
   reg _400540_400540 ; 
   reg __400540_400540;
   reg _400541_400541 ; 
   reg __400541_400541;
   reg _400542_400542 ; 
   reg __400542_400542;
   reg _400543_400543 ; 
   reg __400543_400543;
   reg _400544_400544 ; 
   reg __400544_400544;
   reg _400545_400545 ; 
   reg __400545_400545;
   reg _400546_400546 ; 
   reg __400546_400546;
   reg _400547_400547 ; 
   reg __400547_400547;
   reg _400548_400548 ; 
   reg __400548_400548;
   reg _400549_400549 ; 
   reg __400549_400549;
   reg _400550_400550 ; 
   reg __400550_400550;
   reg _400551_400551 ; 
   reg __400551_400551;
   reg _400552_400552 ; 
   reg __400552_400552;
   reg _400553_400553 ; 
   reg __400553_400553;
   reg _400554_400554 ; 
   reg __400554_400554;
   reg _400555_400555 ; 
   reg __400555_400555;
   reg _400556_400556 ; 
   reg __400556_400556;
   reg _400557_400557 ; 
   reg __400557_400557;
   reg _400558_400558 ; 
   reg __400558_400558;
   reg _400559_400559 ; 
   reg __400559_400559;
   reg _400560_400560 ; 
   reg __400560_400560;
   reg _400561_400561 ; 
   reg __400561_400561;
   reg _400562_400562 ; 
   reg __400562_400562;
   reg _400563_400563 ; 
   reg __400563_400563;
   reg _400564_400564 ; 
   reg __400564_400564;
   reg _400565_400565 ; 
   reg __400565_400565;
   reg _400566_400566 ; 
   reg __400566_400566;
   reg _400567_400567 ; 
   reg __400567_400567;
   reg _400568_400568 ; 
   reg __400568_400568;
   reg _400569_400569 ; 
   reg __400569_400569;
   reg _400570_400570 ; 
   reg __400570_400570;
   reg _400571_400571 ; 
   reg __400571_400571;
   reg _400572_400572 ; 
   reg __400572_400572;
   reg _400573_400573 ; 
   reg __400573_400573;
   reg _400574_400574 ; 
   reg __400574_400574;
   reg _400575_400575 ; 
   reg __400575_400575;
   reg _400576_400576 ; 
   reg __400576_400576;
   reg _400577_400577 ; 
   reg __400577_400577;
   reg _400578_400578 ; 
   reg __400578_400578;
   reg _400579_400579 ; 
   reg __400579_400579;
   reg _400580_400580 ; 
   reg __400580_400580;
   reg _400581_400581 ; 
   reg __400581_400581;
   reg _400582_400582 ; 
   reg __400582_400582;
   reg _400583_400583 ; 
   reg __400583_400583;
   reg _400584_400584 ; 
   reg __400584_400584;
   reg _400585_400585 ; 
   reg __400585_400585;
   reg _400586_400586 ; 
   reg __400586_400586;
   reg _400587_400587 ; 
   reg __400587_400587;
   reg _400588_400588 ; 
   reg __400588_400588;
   reg _400589_400589 ; 
   reg __400589_400589;
   reg _400590_400590 ; 
   reg __400590_400590;
   reg _400591_400591 ; 
   reg __400591_400591;
   reg _400592_400592 ; 
   reg __400592_400592;
   reg _400593_400593 ; 
   reg __400593_400593;
   reg _400594_400594 ; 
   reg __400594_400594;
   reg _400595_400595 ; 
   reg __400595_400595;
   reg _400596_400596 ; 
   reg __400596_400596;
   reg _400597_400597 ; 
   reg __400597_400597;
   reg _400598_400598 ; 
   reg __400598_400598;
   reg _400599_400599 ; 
   reg __400599_400599;
   reg _400600_400600 ; 
   reg __400600_400600;
   reg _400601_400601 ; 
   reg __400601_400601;
   reg _400602_400602 ; 
   reg __400602_400602;
   reg _400603_400603 ; 
   reg __400603_400603;
   reg _400604_400604 ; 
   reg __400604_400604;
   reg _400605_400605 ; 
   reg __400605_400605;
   reg _400606_400606 ; 
   reg __400606_400606;
   reg _400607_400607 ; 
   reg __400607_400607;
   reg _400608_400608 ; 
   reg __400608_400608;
   reg _400609_400609 ; 
   reg __400609_400609;
   reg _400610_400610 ; 
   reg __400610_400610;
   reg _400611_400611 ; 
   reg __400611_400611;
   reg _400612_400612 ; 
   reg __400612_400612;
   reg _400613_400613 ; 
   reg __400613_400613;
   reg _400614_400614 ; 
   reg __400614_400614;
   reg _400615_400615 ; 
   reg __400615_400615;
   reg _400616_400616 ; 
   reg __400616_400616;
   reg _400617_400617 ; 
   reg __400617_400617;
   reg _400618_400618 ; 
   reg __400618_400618;
   reg _400619_400619 ; 
   reg __400619_400619;
   reg _400620_400620 ; 
   reg __400620_400620;
   reg _400621_400621 ; 
   reg __400621_400621;
   reg _400622_400622 ; 
   reg __400622_400622;
   reg _400623_400623 ; 
   reg __400623_400623;
   reg _400624_400624 ; 
   reg __400624_400624;
   reg _400625_400625 ; 
   reg __400625_400625;
   reg _400626_400626 ; 
   reg __400626_400626;
   reg _400627_400627 ; 
   reg __400627_400627;
   reg _400628_400628 ; 
   reg __400628_400628;
   reg _400629_400629 ; 
   reg __400629_400629;
   reg _400630_400630 ; 
   reg __400630_400630;
   reg _400631_400631 ; 
   reg __400631_400631;
   reg _400632_400632 ; 
   reg __400632_400632;
   reg _400633_400633 ; 
   reg __400633_400633;
   reg _400634_400634 ; 
   reg __400634_400634;
   reg _400635_400635 ; 
   reg __400635_400635;
   reg _400636_400636 ; 
   reg __400636_400636;
   reg _400637_400637 ; 
   reg __400637_400637;
   reg _400638_400638 ; 
   reg __400638_400638;
   reg _400639_400639 ; 
   reg __400639_400639;
   reg _400640_400640 ; 
   reg __400640_400640;
   reg _400641_400641 ; 
   reg __400641_400641;
   reg _400642_400642 ; 
   reg __400642_400642;
   reg _400643_400643 ; 
   reg __400643_400643;
   reg _400644_400644 ; 
   reg __400644_400644;
   reg _400645_400645 ; 
   reg __400645_400645;
   reg _400646_400646 ; 
   reg __400646_400646;
   reg _400647_400647 ; 
   reg __400647_400647;
   reg _400648_400648 ; 
   reg __400648_400648;
   reg _400649_400649 ; 
   reg __400649_400649;
   reg _400650_400650 ; 
   reg __400650_400650;
   reg _400651_400651 ; 
   reg __400651_400651;
   reg _400652_400652 ; 
   reg __400652_400652;
   reg _400653_400653 ; 
   reg __400653_400653;
   reg _400654_400654 ; 
   reg __400654_400654;
   reg _400655_400655 ; 
   reg __400655_400655;
   reg _400656_400656 ; 
   reg __400656_400656;
   reg _400657_400657 ; 
   reg __400657_400657;
   reg _400658_400658 ; 
   reg __400658_400658;
   reg _400659_400659 ; 
   reg __400659_400659;
   reg _400660_400660 ; 
   reg __400660_400660;
   reg _400661_400661 ; 
   reg __400661_400661;
   reg _400662_400662 ; 
   reg __400662_400662;
   reg _400663_400663 ; 
   reg __400663_400663;
   reg _400664_400664 ; 
   reg __400664_400664;
   reg _400665_400665 ; 
   reg __400665_400665;
   reg _400666_400666 ; 
   reg __400666_400666;
   reg _400667_400667 ; 
   reg __400667_400667;
   reg _400668_400668 ; 
   reg __400668_400668;
   reg _400669_400669 ; 
   reg __400669_400669;
   reg _400670_400670 ; 
   reg __400670_400670;
   reg _400671_400671 ; 
   reg __400671_400671;
   reg _400672_400672 ; 
   reg __400672_400672;
   reg _400673_400673 ; 
   reg __400673_400673;
   reg _400674_400674 ; 
   reg __400674_400674;
   reg _400675_400675 ; 
   reg __400675_400675;
   reg _400676_400676 ; 
   reg __400676_400676;
   reg _400677_400677 ; 
   reg __400677_400677;
   reg _400678_400678 ; 
   reg __400678_400678;
   reg _400679_400679 ; 
   reg __400679_400679;
   reg _400680_400680 ; 
   reg __400680_400680;
   reg _400681_400681 ; 
   reg __400681_400681;
   reg _400682_400682 ; 
   reg __400682_400682;
   reg _400683_400683 ; 
   reg __400683_400683;
   reg _400684_400684 ; 
   reg __400684_400684;
   reg _400685_400685 ; 
   reg __400685_400685;
   reg _400686_400686 ; 
   reg __400686_400686;
   reg _400687_400687 ; 
   reg __400687_400687;
   reg _400688_400688 ; 
   reg __400688_400688;
   reg _400689_400689 ; 
   reg __400689_400689;
   reg _400690_400690 ; 
   reg __400690_400690;
   reg _400691_400691 ; 
   reg __400691_400691;
   reg _400692_400692 ; 
   reg __400692_400692;
   reg _400693_400693 ; 
   reg __400693_400693;
   reg _400694_400694 ; 
   reg __400694_400694;
   reg _400695_400695 ; 
   reg __400695_400695;
   reg _400696_400696 ; 
   reg __400696_400696;
   reg _400697_400697 ; 
   reg __400697_400697;
   reg _400698_400698 ; 
   reg __400698_400698;
   reg _400699_400699 ; 
   reg __400699_400699;
   reg _400700_400700 ; 
   reg __400700_400700;
   reg _400701_400701 ; 
   reg __400701_400701;
   reg _400702_400702 ; 
   reg __400702_400702;
   reg _400703_400703 ; 
   reg __400703_400703;
   reg _400704_400704 ; 
   reg __400704_400704;
   reg _400705_400705 ; 
   reg __400705_400705;
   reg _400706_400706 ; 
   reg __400706_400706;
   reg _400707_400707 ; 
   reg __400707_400707;
   reg _400708_400708 ; 
   reg __400708_400708;
   reg _400709_400709 ; 
   reg __400709_400709;
   reg _400710_400710 ; 
   reg __400710_400710;
   reg _400711_400711 ; 
   reg __400711_400711;
   reg _400712_400712 ; 
   reg __400712_400712;
   reg _400713_400713 ; 
   reg __400713_400713;
   reg _400714_400714 ; 
   reg __400714_400714;
   reg _400715_400715 ; 
   reg __400715_400715;
   reg _400716_400716 ; 
   reg __400716_400716;
   reg _400717_400717 ; 
   reg __400717_400717;
   reg _400718_400718 ; 
   reg __400718_400718;
   reg _400719_400719 ; 
   reg __400719_400719;
   reg _400720_400720 ; 
   reg __400720_400720;
   reg _400721_400721 ; 
   reg __400721_400721;
   reg _400722_400722 ; 
   reg __400722_400722;
   reg _400723_400723 ; 
   reg __400723_400723;
   reg _400724_400724 ; 
   reg __400724_400724;
   reg _400725_400725 ; 
   reg __400725_400725;
   reg _400726_400726 ; 
   reg __400726_400726;
   reg _400727_400727 ; 
   reg __400727_400727;
   reg _400728_400728 ; 
   reg __400728_400728;
   reg _400729_400729 ; 
   reg __400729_400729;
   reg _400730_400730 ; 
   reg __400730_400730;
   reg _400731_400731 ; 
   reg __400731_400731;
   reg _400732_400732 ; 
   reg __400732_400732;
   reg _400733_400733 ; 
   reg __400733_400733;
   reg _400734_400734 ; 
   reg __400734_400734;
   reg _400735_400735 ; 
   reg __400735_400735;
   reg _400736_400736 ; 
   reg __400736_400736;
   reg _400737_400737 ; 
   reg __400737_400737;
   reg _400738_400738 ; 
   reg __400738_400738;
   reg _400739_400739 ; 
   reg __400739_400739;
   reg _400740_400740 ; 
   reg __400740_400740;
   reg _400741_400741 ; 
   reg __400741_400741;
   reg _400742_400742 ; 
   reg __400742_400742;
   reg _400743_400743 ; 
   reg __400743_400743;
   reg _400744_400744 ; 
   reg __400744_400744;
   reg _400745_400745 ; 
   reg __400745_400745;
   reg _400746_400746 ; 
   reg __400746_400746;
   reg _400747_400747 ; 
   reg __400747_400747;
   reg _400748_400748 ; 
   reg __400748_400748;
   reg _400749_400749 ; 
   reg __400749_400749;
   reg _400750_400750 ; 
   reg __400750_400750;
   reg _400751_400751 ; 
   reg __400751_400751;
   reg _400752_400752 ; 
   reg __400752_400752;
   reg _400753_400753 ; 
   reg __400753_400753;
   reg _400754_400754 ; 
   reg __400754_400754;
   reg _400755_400755 ; 
   reg __400755_400755;
   reg _400756_400756 ; 
   reg __400756_400756;
   reg _400757_400757 ; 
   reg __400757_400757;
   reg _400758_400758 ; 
   reg __400758_400758;
   reg _400759_400759 ; 
   reg __400759_400759;
   reg _400760_400760 ; 
   reg __400760_400760;
   reg _400761_400761 ; 
   reg __400761_400761;
   reg _400762_400762 ; 
   reg __400762_400762;
   reg _400763_400763 ; 
   reg __400763_400763;
   reg _400764_400764 ; 
   reg __400764_400764;
   reg _400765_400765 ; 
   reg __400765_400765;
   reg _400766_400766 ; 
   reg __400766_400766;
   reg _400767_400767 ; 
   reg __400767_400767;
   reg _400768_400768 ; 
   reg __400768_400768;
   reg _400769_400769 ; 
   reg __400769_400769;
   reg _400770_400770 ; 
   reg __400770_400770;
   reg _400771_400771 ; 
   reg __400771_400771;
   reg _400772_400772 ; 
   reg __400772_400772;
   reg _400773_400773 ; 
   reg __400773_400773;
   reg _400774_400774 ; 
   reg __400774_400774;
   reg _400775_400775 ; 
   reg __400775_400775;
   reg _400776_400776 ; 
   reg __400776_400776;
   reg _400777_400777 ; 
   reg __400777_400777;
   reg _400778_400778 ; 
   reg __400778_400778;
   reg _400779_400779 ; 
   reg __400779_400779;
   reg _400780_400780 ; 
   reg __400780_400780;
   reg _400781_400781 ; 
   reg __400781_400781;
   reg _400782_400782 ; 
   reg __400782_400782;
   reg _400783_400783 ; 
   reg __400783_400783;
   reg _400784_400784 ; 
   reg __400784_400784;
   reg _400785_400785 ; 
   reg __400785_400785;
   reg _400786_400786 ; 
   reg __400786_400786;
   reg _400787_400787 ; 
   reg __400787_400787;
   reg _400788_400788 ; 
   reg __400788_400788;
   reg _400789_400789 ; 
   reg __400789_400789;
   reg _400790_400790 ; 
   reg __400790_400790;
   reg _400791_400791 ; 
   reg __400791_400791;
   reg _400792_400792 ; 
   reg __400792_400792;
   reg _400793_400793 ; 
   reg __400793_400793;
   reg _400794_400794 ; 
   reg __400794_400794;
   reg _400795_400795 ; 
   reg __400795_400795;
   reg _400796_400796 ; 
   reg __400796_400796;
   reg _400797_400797 ; 
   reg __400797_400797;
   reg _400798_400798 ; 
   reg __400798_400798;
   reg _400799_400799 ; 
   reg __400799_400799;
   reg _400800_400800 ; 
   reg __400800_400800;
   reg _400801_400801 ; 
   reg __400801_400801;
   reg _400802_400802 ; 
   reg __400802_400802;
   reg _400803_400803 ; 
   reg __400803_400803;
   reg _400804_400804 ; 
   reg __400804_400804;
   reg _400805_400805 ; 
   reg __400805_400805;
   reg _400806_400806 ; 
   reg __400806_400806;
   reg _400807_400807 ; 
   reg __400807_400807;
   reg _400808_400808 ; 
   reg __400808_400808;
   reg _400809_400809 ; 
   reg __400809_400809;
   reg _400810_400810 ; 
   reg __400810_400810;
   reg _400811_400811 ; 
   reg __400811_400811;
   reg _400812_400812 ; 
   reg __400812_400812;
   reg _400813_400813 ; 
   reg __400813_400813;
   reg _400814_400814 ; 
   reg __400814_400814;
   reg _400815_400815 ; 
   reg __400815_400815;
   reg _400816_400816 ; 
   reg __400816_400816;
   reg _400817_400817 ; 
   reg __400817_400817;
   reg _400818_400818 ; 
   reg __400818_400818;
   reg _400819_400819 ; 
   reg __400819_400819;
   reg _400820_400820 ; 
   reg __400820_400820;
   reg _400821_400821 ; 
   reg __400821_400821;
   reg _400822_400822 ; 
   reg __400822_400822;
   reg _400823_400823 ; 
   reg __400823_400823;
   reg _400824_400824 ; 
   reg __400824_400824;
   reg _400825_400825 ; 
   reg __400825_400825;
   reg _400826_400826 ; 
   reg __400826_400826;
   reg _400827_400827 ; 
   reg __400827_400827;
   reg _400828_400828 ; 
   reg __400828_400828;
   reg _400829_400829 ; 
   reg __400829_400829;
   reg _400830_400830 ; 
   reg __400830_400830;
   reg _400831_400831 ; 
   reg __400831_400831;
   reg _400832_400832 ; 
   reg __400832_400832;
   reg _400833_400833 ; 
   reg __400833_400833;
   reg _400834_400834 ; 
   reg __400834_400834;
   reg _400835_400835 ; 
   reg __400835_400835;
   reg _400836_400836 ; 
   reg __400836_400836;
   reg _400837_400837 ; 
   reg __400837_400837;
   reg _400838_400838 ; 
   reg __400838_400838;
   reg _400839_400839 ; 
   reg __400839_400839;
   reg _400840_400840 ; 
   reg __400840_400840;
   reg _400841_400841 ; 
   reg __400841_400841;
   reg _400842_400842 ; 
   reg __400842_400842;
   reg _400843_400843 ; 
   reg __400843_400843;
   reg _400844_400844 ; 
   reg __400844_400844;
   reg _400845_400845 ; 
   reg __400845_400845;
   reg _400846_400846 ; 
   reg __400846_400846;
   reg _400847_400847 ; 
   reg __400847_400847;
   reg _400848_400848 ; 
   reg __400848_400848;
   reg _400849_400849 ; 
   reg __400849_400849;
   reg _400850_400850 ; 
   reg __400850_400850;
   reg _400851_400851 ; 
   reg __400851_400851;
   reg _400852_400852 ; 
   reg __400852_400852;
   reg _400853_400853 ; 
   reg __400853_400853;
   reg _400854_400854 ; 
   reg __400854_400854;
   reg _400855_400855 ; 
   reg __400855_400855;
   reg _400856_400856 ; 
   reg __400856_400856;
   reg _400857_400857 ; 
   reg __400857_400857;
   reg _400858_400858 ; 
   reg __400858_400858;
   reg _400859_400859 ; 
   reg __400859_400859;
   reg _400860_400860 ; 
   reg __400860_400860;
   reg _400861_400861 ; 
   reg __400861_400861;
   reg _400862_400862 ; 
   reg __400862_400862;
   reg _400863_400863 ; 
   reg __400863_400863;
   reg _400864_400864 ; 
   reg __400864_400864;
   reg _400865_400865 ; 
   reg __400865_400865;
   reg _400866_400866 ; 
   reg __400866_400866;
   reg _400867_400867 ; 
   reg __400867_400867;
   reg _400868_400868 ; 
   reg __400868_400868;
   reg _400869_400869 ; 
   reg __400869_400869;
   reg _400870_400870 ; 
   reg __400870_400870;
   reg _400871_400871 ; 
   reg __400871_400871;
   reg _400872_400872 ; 
   reg __400872_400872;
   reg _400873_400873 ; 
   reg __400873_400873;
   reg _400874_400874 ; 
   reg __400874_400874;
   reg _400875_400875 ; 
   reg __400875_400875;
   reg _400876_400876 ; 
   reg __400876_400876;
   reg _400877_400877 ; 
   reg __400877_400877;
   reg _400878_400878 ; 
   reg __400878_400878;
   reg _400879_400879 ; 
   reg __400879_400879;
   reg _400880_400880 ; 
   reg __400880_400880;
   reg _400881_400881 ; 
   reg __400881_400881;
   reg _400882_400882 ; 
   reg __400882_400882;
   reg _400883_400883 ; 
   reg __400883_400883;
   reg _400884_400884 ; 
   reg __400884_400884;
   reg _400885_400885 ; 
   reg __400885_400885;
   reg _400886_400886 ; 
   reg __400886_400886;
   reg _400887_400887 ; 
   reg __400887_400887;
   reg _400888_400888 ; 
   reg __400888_400888;
   reg _400889_400889 ; 
   reg __400889_400889;
   reg _400890_400890 ; 
   reg __400890_400890;
   reg _400891_400891 ; 
   reg __400891_400891;
   reg _400892_400892 ; 
   reg __400892_400892;
   reg _400893_400893 ; 
   reg __400893_400893;
   reg _400894_400894 ; 
   reg __400894_400894;
   reg _400895_400895 ; 
   reg __400895_400895;
   reg _400896_400896 ; 
   reg __400896_400896;
   reg _400897_400897 ; 
   reg __400897_400897;
   reg _400898_400898 ; 
   reg __400898_400898;
   reg _400899_400899 ; 
   reg __400899_400899;
   reg _400900_400900 ; 
   reg __400900_400900;
   reg _400901_400901 ; 
   reg __400901_400901;
   reg _400902_400902 ; 
   reg __400902_400902;
   reg _400903_400903 ; 
   reg __400903_400903;
   reg _400904_400904 ; 
   reg __400904_400904;
   reg _400905_400905 ; 
   reg __400905_400905;
   reg _400906_400906 ; 
   reg __400906_400906;
   reg _400907_400907 ; 
   reg __400907_400907;
   reg _400908_400908 ; 
   reg __400908_400908;
   reg _400909_400909 ; 
   reg __400909_400909;
   reg _400910_400910 ; 
   reg __400910_400910;
   reg _400911_400911 ; 
   reg __400911_400911;
   reg _400912_400912 ; 
   reg __400912_400912;
   reg _400913_400913 ; 
   reg __400913_400913;
   reg _400914_400914 ; 
   reg __400914_400914;
   reg _400915_400915 ; 
   reg __400915_400915;
   reg _400916_400916 ; 
   reg __400916_400916;
   reg _400917_400917 ; 
   reg __400917_400917;
   reg _400918_400918 ; 
   reg __400918_400918;
   reg _400919_400919 ; 
   reg __400919_400919;
   reg _400920_400920 ; 
   reg __400920_400920;
   reg _400921_400921 ; 
   reg __400921_400921;
   reg _400922_400922 ; 
   reg __400922_400922;
   reg _400923_400923 ; 
   reg __400923_400923;
   reg _400924_400924 ; 
   reg __400924_400924;
   reg _400925_400925 ; 
   reg __400925_400925;
   reg _400926_400926 ; 
   reg __400926_400926;
   reg _400927_400927 ; 
   reg __400927_400927;
   reg _400928_400928 ; 
   reg __400928_400928;
   reg _400929_400929 ; 
   reg __400929_400929;
   reg _400930_400930 ; 
   reg __400930_400930;
   reg _400931_400931 ; 
   reg __400931_400931;
   reg _400932_400932 ; 
   reg __400932_400932;
   reg _400933_400933 ; 
   reg __400933_400933;
   reg _400934_400934 ; 
   reg __400934_400934;
   reg _400935_400935 ; 
   reg __400935_400935;
   reg _400936_400936 ; 
   reg __400936_400936;
   reg _400937_400937 ; 
   reg __400937_400937;
   reg _400938_400938 ; 
   reg __400938_400938;
   reg _400939_400939 ; 
   reg __400939_400939;
   reg _400940_400940 ; 
   reg __400940_400940;
   reg _400941_400941 ; 
   reg __400941_400941;
   reg _400942_400942 ; 
   reg __400942_400942;
   reg _400943_400943 ; 
   reg __400943_400943;
   reg _400944_400944 ; 
   reg __400944_400944;
   reg _400945_400945 ; 
   reg __400945_400945;
   reg _400946_400946 ; 
   reg __400946_400946;
   reg _400947_400947 ; 
   reg __400947_400947;
   reg _400948_400948 ; 
   reg __400948_400948;
   reg _400949_400949 ; 
   reg __400949_400949;
   reg _400950_400950 ; 
   reg __400950_400950;
   reg _400951_400951 ; 
   reg __400951_400951;
   reg _400952_400952 ; 
   reg __400952_400952;
   reg _400953_400953 ; 
   reg __400953_400953;
   reg _400954_400954 ; 
   reg __400954_400954;
   reg _400955_400955 ; 
   reg __400955_400955;
   reg _400956_400956 ; 
   reg __400956_400956;
   reg _400957_400957 ; 
   reg __400957_400957;
   reg _400958_400958 ; 
   reg __400958_400958;
   reg _400959_400959 ; 
   reg __400959_400959;
   reg _400960_400960 ; 
   reg __400960_400960;
   reg _400961_400961 ; 
   reg __400961_400961;
   reg _400962_400962 ; 
   reg __400962_400962;
   reg _400963_400963 ; 
   reg __400963_400963;
   reg _400964_400964 ; 
   reg __400964_400964;
   reg _400965_400965 ; 
   reg __400965_400965;
   reg _400966_400966 ; 
   reg __400966_400966;
   reg _400967_400967 ; 
   reg __400967_400967;
   reg _400968_400968 ; 
   reg __400968_400968;
   reg _400969_400969 ; 
   reg __400969_400969;
   reg _400970_400970 ; 
   reg __400970_400970;
   reg _400971_400971 ; 
   reg __400971_400971;
   reg _400972_400972 ; 
   reg __400972_400972;
   reg _400973_400973 ; 
   reg __400973_400973;
   reg _400974_400974 ; 
   reg __400974_400974;
   reg _400975_400975 ; 
   reg __400975_400975;
   reg _400976_400976 ; 
   reg __400976_400976;
   reg _400977_400977 ; 
   reg __400977_400977;
   reg _400978_400978 ; 
   reg __400978_400978;
   reg _400979_400979 ; 
   reg __400979_400979;
   reg _400980_400980 ; 
   reg __400980_400980;
   reg _400981_400981 ; 
   reg __400981_400981;
   reg _400982_400982 ; 
   reg __400982_400982;
   reg _400983_400983 ; 
   reg __400983_400983;
   reg _400984_400984 ; 
   reg __400984_400984;
   reg _400985_400985 ; 
   reg __400985_400985;
   reg _400986_400986 ; 
   reg __400986_400986;
   reg _400987_400987 ; 
   reg __400987_400987;
   reg _400988_400988 ; 
   reg __400988_400988;
   reg _400989_400989 ; 
   reg __400989_400989;
   reg _400990_400990 ; 
   reg __400990_400990;
   reg _400991_400991 ; 
   reg __400991_400991;
   reg _400992_400992 ; 
   reg __400992_400992;
   reg _400993_400993 ; 
   reg __400993_400993;
   reg _400994_400994 ; 
   reg __400994_400994;
   reg _400995_400995 ; 
   reg __400995_400995;
   reg _400996_400996 ; 
   reg __400996_400996;
   reg _400997_400997 ; 
   reg __400997_400997;
   reg _400998_400998 ; 
   reg __400998_400998;
   reg _400999_400999 ; 
   reg __400999_400999;
   reg _401000_401000 ; 
   reg __401000_401000;
   reg _401001_401001 ; 
   reg __401001_401001;
   reg _401002_401002 ; 
   reg __401002_401002;
   reg _401003_401003 ; 
   reg __401003_401003;
   reg _401004_401004 ; 
   reg __401004_401004;
   reg _401005_401005 ; 
   reg __401005_401005;
   reg _401006_401006 ; 
   reg __401006_401006;
   reg _401007_401007 ; 
   reg __401007_401007;
   reg _401008_401008 ; 
   reg __401008_401008;
   reg _401009_401009 ; 
   reg __401009_401009;
   reg _401010_401010 ; 
   reg __401010_401010;
   reg _401011_401011 ; 
   reg __401011_401011;
   reg _401012_401012 ; 
   reg __401012_401012;
   reg _401013_401013 ; 
   reg __401013_401013;
   reg _401014_401014 ; 
   reg __401014_401014;
   reg _401015_401015 ; 
   reg __401015_401015;
   reg _401016_401016 ; 
   reg __401016_401016;
   reg _401017_401017 ; 
   reg __401017_401017;
   reg _401018_401018 ; 
   reg __401018_401018;
   reg _401019_401019 ; 
   reg __401019_401019;
   reg _401020_401020 ; 
   reg __401020_401020;
   reg _401021_401021 ; 
   reg __401021_401021;
   reg _401022_401022 ; 
   reg __401022_401022;
   reg _401023_401023 ; 
   reg __401023_401023;
   reg _401024_401024 ; 
   reg __401024_401024;
   reg _401025_401025 ; 
   reg __401025_401025;
   reg _401026_401026 ; 
   reg __401026_401026;
   reg _401027_401027 ; 
   reg __401027_401027;
   reg _401028_401028 ; 
   reg __401028_401028;
   reg _401029_401029 ; 
   reg __401029_401029;
   reg _401030_401030 ; 
   reg __401030_401030;
   reg _401031_401031 ; 
   reg __401031_401031;
   reg _401032_401032 ; 
   reg __401032_401032;
   reg _401033_401033 ; 
   reg __401033_401033;
   reg _401034_401034 ; 
   reg __401034_401034;
   reg _401035_401035 ; 
   reg __401035_401035;
   reg _401036_401036 ; 
   reg __401036_401036;
   reg _401037_401037 ; 
   reg __401037_401037;
   reg _401038_401038 ; 
   reg __401038_401038;
   reg _401039_401039 ; 
   reg __401039_401039;
   reg _401040_401040 ; 
   reg __401040_401040;
   reg _401041_401041 ; 
   reg __401041_401041;
   reg _401042_401042 ; 
   reg __401042_401042;
   reg _401043_401043 ; 
   reg __401043_401043;
   reg _401044_401044 ; 
   reg __401044_401044;
   reg _401045_401045 ; 
   reg __401045_401045;
   reg _401046_401046 ; 
   reg __401046_401046;
   reg _401047_401047 ; 
   reg __401047_401047;
   reg _401048_401048 ; 
   reg __401048_401048;
   reg _401049_401049 ; 
   reg __401049_401049;
   reg _401050_401050 ; 
   reg __401050_401050;
   reg _401051_401051 ; 
   reg __401051_401051;
   reg _401052_401052 ; 
   reg __401052_401052;
   reg _401053_401053 ; 
   reg __401053_401053;
   reg _401054_401054 ; 
   reg __401054_401054;
   reg _401055_401055 ; 
   reg __401055_401055;
   reg _401056_401056 ; 
   reg __401056_401056;
   reg _401057_401057 ; 
   reg __401057_401057;
   reg _401058_401058 ; 
   reg __401058_401058;
   reg _401059_401059 ; 
   reg __401059_401059;
   reg _401060_401060 ; 
   reg __401060_401060;
   reg _401061_401061 ; 
   reg __401061_401061;
   reg _401062_401062 ; 
   reg __401062_401062;
   reg _401063_401063 ; 
   reg __401063_401063;
   reg _401064_401064 ; 
   reg __401064_401064;
   reg _401065_401065 ; 
   reg __401065_401065;
   reg _401066_401066 ; 
   reg __401066_401066;
   reg _401067_401067 ; 
   reg __401067_401067;
   reg _401068_401068 ; 
   reg __401068_401068;
   reg _401069_401069 ; 
   reg __401069_401069;
   reg _401070_401070 ; 
   reg __401070_401070;
   reg _401071_401071 ; 
   reg __401071_401071;
   reg _401072_401072 ; 
   reg __401072_401072;
   reg _401073_401073 ; 
   reg __401073_401073;
   reg _401074_401074 ; 
   reg __401074_401074;
   reg _401075_401075 ; 
   reg __401075_401075;
   reg _401076_401076 ; 
   reg __401076_401076;
   reg _401077_401077 ; 
   reg __401077_401077;
   reg _401078_401078 ; 
   reg __401078_401078;
   reg _401079_401079 ; 
   reg __401079_401079;
   reg _401080_401080 ; 
   reg __401080_401080;
   reg _401081_401081 ; 
   reg __401081_401081;
   reg _401082_401082 ; 
   reg __401082_401082;
   reg _401083_401083 ; 
   reg __401083_401083;
   reg _401084_401084 ; 
   reg __401084_401084;
   reg _401085_401085 ; 
   reg __401085_401085;
   reg _401086_401086 ; 
   reg __401086_401086;
   reg _401087_401087 ; 
   reg __401087_401087;
   reg _401088_401088 ; 
   reg __401088_401088;
   reg _401089_401089 ; 
   reg __401089_401089;
   reg _401090_401090 ; 
   reg __401090_401090;
   reg _401091_401091 ; 
   reg __401091_401091;
   reg _401092_401092 ; 
   reg __401092_401092;
   reg _401093_401093 ; 
   reg __401093_401093;
   reg _401094_401094 ; 
   reg __401094_401094;
   reg _401095_401095 ; 
   reg __401095_401095;
   reg _401096_401096 ; 
   reg __401096_401096;
   reg _401097_401097 ; 
   reg __401097_401097;
   reg _401098_401098 ; 
   reg __401098_401098;
   reg _401099_401099 ; 
   reg __401099_401099;
   reg _401100_401100 ; 
   reg __401100_401100;
   reg _401101_401101 ; 
   reg __401101_401101;
   reg _401102_401102 ; 
   reg __401102_401102;
   reg _401103_401103 ; 
   reg __401103_401103;
   reg _401104_401104 ; 
   reg __401104_401104;
   reg _401105_401105 ; 
   reg __401105_401105;
   reg _401106_401106 ; 
   reg __401106_401106;
   reg _401107_401107 ; 
   reg __401107_401107;
   reg _401108_401108 ; 
   reg __401108_401108;
   reg _401109_401109 ; 
   reg __401109_401109;
   reg _401110_401110 ; 
   reg __401110_401110;
   reg _401111_401111 ; 
   reg __401111_401111;
   reg _401112_401112 ; 
   reg __401112_401112;
   reg _401113_401113 ; 
   reg __401113_401113;
   reg _401114_401114 ; 
   reg __401114_401114;
   reg _401115_401115 ; 
   reg __401115_401115;
   reg _401116_401116 ; 
   reg __401116_401116;
   reg _401117_401117 ; 
   reg __401117_401117;
   reg _401118_401118 ; 
   reg __401118_401118;
   reg _401119_401119 ; 
   reg __401119_401119;
   reg _401120_401120 ; 
   reg __401120_401120;
   reg _401121_401121 ; 
   reg __401121_401121;
   reg _401122_401122 ; 
   reg __401122_401122;
   reg _401123_401123 ; 
   reg __401123_401123;
   reg _401124_401124 ; 
   reg __401124_401124;
   reg _401125_401125 ; 
   reg __401125_401125;
   reg _401126_401126 ; 
   reg __401126_401126;
   reg _401127_401127 ; 
   reg __401127_401127;
   reg _401128_401128 ; 
   reg __401128_401128;
   reg _401129_401129 ; 
   reg __401129_401129;
   reg _401130_401130 ; 
   reg __401130_401130;
   reg _401131_401131 ; 
   reg __401131_401131;
   reg _401132_401132 ; 
   reg __401132_401132;
   reg _401133_401133 ; 
   reg __401133_401133;
   reg _401134_401134 ; 
   reg __401134_401134;
   reg _401135_401135 ; 
   reg __401135_401135;
   reg _401136_401136 ; 
   reg __401136_401136;
   reg _401137_401137 ; 
   reg __401137_401137;
   reg _401138_401138 ; 
   reg __401138_401138;
   reg _401139_401139 ; 
   reg __401139_401139;
   reg _401140_401140 ; 
   reg __401140_401140;
   reg _401141_401141 ; 
   reg __401141_401141;
   reg _401142_401142 ; 
   reg __401142_401142;
   reg _401143_401143 ; 
   reg __401143_401143;
   reg _401144_401144 ; 
   reg __401144_401144;
   reg _401145_401145 ; 
   reg __401145_401145;
   reg _401146_401146 ; 
   reg __401146_401146;
   reg _401147_401147 ; 
   reg __401147_401147;
   reg _401148_401148 ; 
   reg __401148_401148;
   reg _401149_401149 ; 
   reg __401149_401149;
   reg _401150_401150 ; 
   reg __401150_401150;
   reg _401151_401151 ; 
   reg __401151_401151;
   reg _401152_401152 ; 
   reg __401152_401152;
   reg _401153_401153 ; 
   reg __401153_401153;
   reg _401154_401154 ; 
   reg __401154_401154;
   reg _401155_401155 ; 
   reg __401155_401155;
   reg _401156_401156 ; 
   reg __401156_401156;
   reg _401157_401157 ; 
   reg __401157_401157;
   reg _401158_401158 ; 
   reg __401158_401158;
   reg _401159_401159 ; 
   reg __401159_401159;
   reg _401160_401160 ; 
   reg __401160_401160;
   reg _401161_401161 ; 
   reg __401161_401161;
   reg _401162_401162 ; 
   reg __401162_401162;
   reg _401163_401163 ; 
   reg __401163_401163;
   reg _401164_401164 ; 
   reg __401164_401164;
   reg _401165_401165 ; 
   reg __401165_401165;
   reg _401166_401166 ; 
   reg __401166_401166;
   reg _401167_401167 ; 
   reg __401167_401167;
   reg _401168_401168 ; 
   reg __401168_401168;
   reg _401169_401169 ; 
   reg __401169_401169;
   reg _401170_401170 ; 
   reg __401170_401170;
   reg _401171_401171 ; 
   reg __401171_401171;
   reg _401172_401172 ; 
   reg __401172_401172;
   reg _401173_401173 ; 
   reg __401173_401173;
   reg _401174_401174 ; 
   reg __401174_401174;
   reg _401175_401175 ; 
   reg __401175_401175;
   reg _401176_401176 ; 
   reg __401176_401176;
   reg _401177_401177 ; 
   reg __401177_401177;
   reg _401178_401178 ; 
   reg __401178_401178;
   reg _401179_401179 ; 
   reg __401179_401179;
   reg _401180_401180 ; 
   reg __401180_401180;
   reg _401181_401181 ; 
   reg __401181_401181;
   reg _401182_401182 ; 
   reg __401182_401182;
   reg _401183_401183 ; 
   reg __401183_401183;
   reg _401184_401184 ; 
   reg __401184_401184;
   reg _401185_401185 ; 
   reg __401185_401185;
   reg _401186_401186 ; 
   reg __401186_401186;
   reg _401187_401187 ; 
   reg __401187_401187;
   reg _401188_401188 ; 
   reg __401188_401188;
   reg _401189_401189 ; 
   reg __401189_401189;
   reg _401190_401190 ; 
   reg __401190_401190;
   reg _401191_401191 ; 
   reg __401191_401191;
   reg _401192_401192 ; 
   reg __401192_401192;
   reg _401193_401193 ; 
   reg __401193_401193;
   reg _401194_401194 ; 
   reg __401194_401194;
   reg _401195_401195 ; 
   reg __401195_401195;
   reg _401196_401196 ; 
   reg __401196_401196;
   reg _401197_401197 ; 
   reg __401197_401197;
   reg _401198_401198 ; 
   reg __401198_401198;
   reg _401199_401199 ; 
   reg __401199_401199;
   reg _401200_401200 ; 
   reg __401200_401200;
   reg _401201_401201 ; 
   reg __401201_401201;
   reg _401202_401202 ; 
   reg __401202_401202;
   reg _401203_401203 ; 
   reg __401203_401203;
   reg _401204_401204 ; 
   reg __401204_401204;
   reg _401205_401205 ; 
   reg __401205_401205;
   reg _401206_401206 ; 
   reg __401206_401206;
   reg _401207_401207 ; 
   reg __401207_401207;
   reg _401208_401208 ; 
   reg __401208_401208;
   reg _401209_401209 ; 
   reg __401209_401209;
   reg _401210_401210 ; 
   reg __401210_401210;
   reg _401211_401211 ; 
   reg __401211_401211;
   reg _401212_401212 ; 
   reg __401212_401212;
   reg _401213_401213 ; 
   reg __401213_401213;
   reg _401214_401214 ; 
   reg __401214_401214;
   reg _401215_401215 ; 
   reg __401215_401215;
   reg _401216_401216 ; 
   reg __401216_401216;
   reg _401217_401217 ; 
   reg __401217_401217;
   reg _401218_401218 ; 
   reg __401218_401218;
   reg _401219_401219 ; 
   reg __401219_401219;
   reg _401220_401220 ; 
   reg __401220_401220;
   reg _401221_401221 ; 
   reg __401221_401221;
   reg _401222_401222 ; 
   reg __401222_401222;
   reg _401223_401223 ; 
   reg __401223_401223;
   reg _401224_401224 ; 
   reg __401224_401224;
   reg _401225_401225 ; 
   reg __401225_401225;
   reg _401226_401226 ; 
   reg __401226_401226;
   reg _401227_401227 ; 
   reg __401227_401227;
   reg _401228_401228 ; 
   reg __401228_401228;
   reg _401229_401229 ; 
   reg __401229_401229;
   reg _401230_401230 ; 
   reg __401230_401230;
   reg _401231_401231 ; 
   reg __401231_401231;
   reg _401232_401232 ; 
   reg __401232_401232;
   reg _401233_401233 ; 
   reg __401233_401233;
   reg _401234_401234 ; 
   reg __401234_401234;
   reg _401235_401235 ; 
   reg __401235_401235;
   reg _401236_401236 ; 
   reg __401236_401236;
   reg _401237_401237 ; 
   reg __401237_401237;
   reg _401238_401238 ; 
   reg __401238_401238;
   reg _401239_401239 ; 
   reg __401239_401239;
   reg _401240_401240 ; 
   reg __401240_401240;
   reg _401241_401241 ; 
   reg __401241_401241;
   reg _401242_401242 ; 
   reg __401242_401242;
   reg _401243_401243 ; 
   reg __401243_401243;
   reg _401244_401244 ; 
   reg __401244_401244;
   reg _401245_401245 ; 
   reg __401245_401245;
   reg _401246_401246 ; 
   reg __401246_401246;
   reg _401247_401247 ; 
   reg __401247_401247;
   reg _401248_401248 ; 
   reg __401248_401248;
   reg _401249_401249 ; 
   reg __401249_401249;
   reg _401250_401250 ; 
   reg __401250_401250;
   reg _401251_401251 ; 
   reg __401251_401251;
   reg _401252_401252 ; 
   reg __401252_401252;
   reg _401253_401253 ; 
   reg __401253_401253;
   reg _401254_401254 ; 
   reg __401254_401254;
   reg _401255_401255 ; 
   reg __401255_401255;
   reg _401256_401256 ; 
   reg __401256_401256;
   reg _401257_401257 ; 
   reg __401257_401257;
   reg _401258_401258 ; 
   reg __401258_401258;
   reg _401259_401259 ; 
   reg __401259_401259;
   reg _401260_401260 ; 
   reg __401260_401260;
   reg _401261_401261 ; 
   reg __401261_401261;
   reg _401262_401262 ; 
   reg __401262_401262;
   reg _401263_401263 ; 
   reg __401263_401263;
   reg _401264_401264 ; 
   reg __401264_401264;
   reg _401265_401265 ; 
   reg __401265_401265;
   reg _401266_401266 ; 
   reg __401266_401266;
   reg _401267_401267 ; 
   reg __401267_401267;
   reg _401268_401268 ; 
   reg __401268_401268;
   reg _401269_401269 ; 
   reg __401269_401269;
   reg _401270_401270 ; 
   reg __401270_401270;
   reg _401271_401271 ; 
   reg __401271_401271;
   reg _401272_401272 ; 
   reg __401272_401272;
   reg _401273_401273 ; 
   reg __401273_401273;
   reg _401274_401274 ; 
   reg __401274_401274;
   reg _401275_401275 ; 
   reg __401275_401275;
   reg _401276_401276 ; 
   reg __401276_401276;
   reg _401277_401277 ; 
   reg __401277_401277;
   reg _401278_401278 ; 
   reg __401278_401278;
   reg _401279_401279 ; 
   reg __401279_401279;
   reg _401280_401280 ; 
   reg __401280_401280;
   reg _401281_401281 ; 
   reg __401281_401281;
   reg _401282_401282 ; 
   reg __401282_401282;
   reg _401283_401283 ; 
   reg __401283_401283;
   reg _401284_401284 ; 
   reg __401284_401284;
   reg _401285_401285 ; 
   reg __401285_401285;
   reg _401286_401286 ; 
   reg __401286_401286;
   reg _401287_401287 ; 
   reg __401287_401287;
   reg _401288_401288 ; 
   reg __401288_401288;
   reg _401289_401289 ; 
   reg __401289_401289;
   reg _401290_401290 ; 
   reg __401290_401290;
   reg _401291_401291 ; 
   reg __401291_401291;
   reg _401292_401292 ; 
   reg __401292_401292;
   reg _401293_401293 ; 
   reg __401293_401293;
   reg _401294_401294 ; 
   reg __401294_401294;
   reg _401295_401295 ; 
   reg __401295_401295;
   reg _401296_401296 ; 
   reg __401296_401296;
   reg _401297_401297 ; 
   reg __401297_401297;
   reg _401298_401298 ; 
   reg __401298_401298;
   reg _401299_401299 ; 
   reg __401299_401299;
   reg _401300_401300 ; 
   reg __401300_401300;
   reg _401301_401301 ; 
   reg __401301_401301;
   reg _401302_401302 ; 
   reg __401302_401302;
   reg _401303_401303 ; 
   reg __401303_401303;
   reg _401304_401304 ; 
   reg __401304_401304;
   reg _401305_401305 ; 
   reg __401305_401305;
   reg _401306_401306 ; 
   reg __401306_401306;
   reg _401307_401307 ; 
   reg __401307_401307;
   reg _401308_401308 ; 
   reg __401308_401308;
   reg _401309_401309 ; 
   reg __401309_401309;
   reg _401310_401310 ; 
   reg __401310_401310;
   reg _401311_401311 ; 
   reg __401311_401311;
   reg _401312_401312 ; 
   reg __401312_401312;
   reg _401313_401313 ; 
   reg __401313_401313;
   reg _401314_401314 ; 
   reg __401314_401314;
   reg _401315_401315 ; 
   reg __401315_401315;
   reg _401316_401316 ; 
   reg __401316_401316;
   reg _401317_401317 ; 
   reg __401317_401317;
   reg _401318_401318 ; 
   reg __401318_401318;
   reg _401319_401319 ; 
   reg __401319_401319;
   reg _401320_401320 ; 
   reg __401320_401320;
   reg _401321_401321 ; 
   reg __401321_401321;
   reg _401322_401322 ; 
   reg __401322_401322;
   reg _401323_401323 ; 
   reg __401323_401323;
   reg _401324_401324 ; 
   reg __401324_401324;
   reg _401325_401325 ; 
   reg __401325_401325;
   reg _401326_401326 ; 
   reg __401326_401326;
   reg _401327_401327 ; 
   reg __401327_401327;
   reg _401328_401328 ; 
   reg __401328_401328;
   reg _401329_401329 ; 
   reg __401329_401329;
   reg _401330_401330 ; 
   reg __401330_401330;
   reg _401331_401331 ; 
   reg __401331_401331;
   reg _401332_401332 ; 
   reg __401332_401332;
   reg _401333_401333 ; 
   reg __401333_401333;
   reg _401334_401334 ; 
   reg __401334_401334;
   reg _401335_401335 ; 
   reg __401335_401335;
   reg _401336_401336 ; 
   reg __401336_401336;
   reg _401337_401337 ; 
   reg __401337_401337;
   reg _401338_401338 ; 
   reg __401338_401338;
   reg _401339_401339 ; 
   reg __401339_401339;
   reg _401340_401340 ; 
   reg __401340_401340;
   reg _401341_401341 ; 
   reg __401341_401341;
   reg _401342_401342 ; 
   reg __401342_401342;
   reg _401343_401343 ; 
   reg __401343_401343;
   reg _401344_401344 ; 
   reg __401344_401344;
   reg _401345_401345 ; 
   reg __401345_401345;
   reg _401346_401346 ; 
   reg __401346_401346;
   reg _401347_401347 ; 
   reg __401347_401347;
   reg _401348_401348 ; 
   reg __401348_401348;
   reg _401349_401349 ; 
   reg __401349_401349;
   reg _401350_401350 ; 
   reg __401350_401350;
   reg _401351_401351 ; 
   reg __401351_401351;
   reg _401352_401352 ; 
   reg __401352_401352;
   reg _401353_401353 ; 
   reg __401353_401353;
   reg _401354_401354 ; 
   reg __401354_401354;
   reg _401355_401355 ; 
   reg __401355_401355;
   reg _401356_401356 ; 
   reg __401356_401356;
   reg _401357_401357 ; 
   reg __401357_401357;
   reg _401358_401358 ; 
   reg __401358_401358;
   reg _401359_401359 ; 
   reg __401359_401359;
   reg _401360_401360 ; 
   reg __401360_401360;
   reg _401361_401361 ; 
   reg __401361_401361;
   reg _401362_401362 ; 
   reg __401362_401362;
   reg _401363_401363 ; 
   reg __401363_401363;
   reg _401364_401364 ; 
   reg __401364_401364;
   reg _401365_401365 ; 
   reg __401365_401365;
   reg _401366_401366 ; 
   reg __401366_401366;
   reg _401367_401367 ; 
   reg __401367_401367;
   reg _401368_401368 ; 
   reg __401368_401368;
   reg _401369_401369 ; 
   reg __401369_401369;
   reg _401370_401370 ; 
   reg __401370_401370;
   reg _401371_401371 ; 
   reg __401371_401371;
   reg _401372_401372 ; 
   reg __401372_401372;
   reg _401373_401373 ; 
   reg __401373_401373;
   reg _401374_401374 ; 
   reg __401374_401374;
   reg _401375_401375 ; 
   reg __401375_401375;
   reg _401376_401376 ; 
   reg __401376_401376;
   reg _401377_401377 ; 
   reg __401377_401377;
   reg _401378_401378 ; 
   reg __401378_401378;
   reg _401379_401379 ; 
   reg __401379_401379;
   reg _401380_401380 ; 
   reg __401380_401380;
   reg _401381_401381 ; 
   reg __401381_401381;
   reg _401382_401382 ; 
   reg __401382_401382;
   reg _401383_401383 ; 
   reg __401383_401383;
   reg _401384_401384 ; 
   reg __401384_401384;
   reg _401385_401385 ; 
   reg __401385_401385;
   reg _401386_401386 ; 
   reg __401386_401386;
   reg _401387_401387 ; 
   reg __401387_401387;
   reg _401388_401388 ; 
   reg __401388_401388;
   reg _401389_401389 ; 
   reg __401389_401389;
   reg _401390_401390 ; 
   reg __401390_401390;
   reg _401391_401391 ; 
   reg __401391_401391;
   reg _401392_401392 ; 
   reg __401392_401392;
   reg _401393_401393 ; 
   reg __401393_401393;
   reg _401394_401394 ; 
   reg __401394_401394;
   reg _401395_401395 ; 
   reg __401395_401395;
   reg _401396_401396 ; 
   reg __401396_401396;
   reg _401397_401397 ; 
   reg __401397_401397;
   reg _401398_401398 ; 
   reg __401398_401398;
   reg _401399_401399 ; 
   reg __401399_401399;
   reg _401400_401400 ; 
   reg __401400_401400;
   reg _401401_401401 ; 
   reg __401401_401401;
   reg _401402_401402 ; 
   reg __401402_401402;
   reg _401403_401403 ; 
   reg __401403_401403;
   reg _401404_401404 ; 
   reg __401404_401404;
   reg _401405_401405 ; 
   reg __401405_401405;
   reg _401406_401406 ; 
   reg __401406_401406;
   reg _401407_401407 ; 
   reg __401407_401407;
   reg _401408_401408 ; 
   reg __401408_401408;
   reg _401409_401409 ; 
   reg __401409_401409;
   reg _401410_401410 ; 
   reg __401410_401410;
   reg _401411_401411 ; 
   reg __401411_401411;
   reg _401412_401412 ; 
   reg __401412_401412;
   reg _401413_401413 ; 
   reg __401413_401413;
   reg _401414_401414 ; 
   reg __401414_401414;
   reg _401415_401415 ; 
   reg __401415_401415;
   reg _401416_401416 ; 
   reg __401416_401416;
   reg _401417_401417 ; 
   reg __401417_401417;
   reg _401418_401418 ; 
   reg __401418_401418;
   reg _401419_401419 ; 
   reg __401419_401419;
   reg _401420_401420 ; 
   reg __401420_401420;
   reg _401421_401421 ; 
   reg __401421_401421;
   reg _401422_401422 ; 
   reg __401422_401422;
   reg _401423_401423 ; 
   reg __401423_401423;
   reg _401424_401424 ; 
   reg __401424_401424;
   reg _401425_401425 ; 
   reg __401425_401425;
   reg _401426_401426 ; 
   reg __401426_401426;
   reg _401427_401427 ; 
   reg __401427_401427;
   reg _401428_401428 ; 
   reg __401428_401428;
   reg _401429_401429 ; 
   reg __401429_401429;
   reg _401430_401430 ; 
   reg __401430_401430;
   reg _401431_401431 ; 
   reg __401431_401431;
   reg _401432_401432 ; 
   reg __401432_401432;
   reg _401433_401433 ; 
   reg __401433_401433;
   reg _401434_401434 ; 
   reg __401434_401434;
   reg _401435_401435 ; 
   reg __401435_401435;
   reg _401436_401436 ; 
   reg __401436_401436;
   reg _401437_401437 ; 
   reg __401437_401437;
   reg _401438_401438 ; 
   reg __401438_401438;
   reg _401439_401439 ; 
   reg __401439_401439;
   reg _401440_401440 ; 
   reg __401440_401440;
   reg _401441_401441 ; 
   reg __401441_401441;
   reg _401442_401442 ; 
   reg __401442_401442;
   reg _401443_401443 ; 
   reg __401443_401443;
   reg _401444_401444 ; 
   reg __401444_401444;
   reg _401445_401445 ; 
   reg __401445_401445;
   reg _401446_401446 ; 
   reg __401446_401446;
   reg _401447_401447 ; 
   reg __401447_401447;
   reg _401448_401448 ; 
   reg __401448_401448;
   reg _401449_401449 ; 
   reg __401449_401449;
   reg _401450_401450 ; 
   reg __401450_401450;
   reg _401451_401451 ; 
   reg __401451_401451;
   reg _401452_401452 ; 
   reg __401452_401452;
   reg _401453_401453 ; 
   reg __401453_401453;
   reg _401454_401454 ; 
   reg __401454_401454;
   reg _401455_401455 ; 
   reg __401455_401455;
   reg _401456_401456 ; 
   reg __401456_401456;
   reg _401457_401457 ; 
   reg __401457_401457;
   reg _401458_401458 ; 
   reg __401458_401458;
   reg _401459_401459 ; 
   reg __401459_401459;
   reg _401460_401460 ; 
   reg __401460_401460;
   reg _401461_401461 ; 
   reg __401461_401461;
   reg _401462_401462 ; 
   reg __401462_401462;
   reg _401463_401463 ; 
   reg __401463_401463;
   reg _401464_401464 ; 
   reg __401464_401464;
   reg _401465_401465 ; 
   reg __401465_401465;
   reg _401466_401466 ; 
   reg __401466_401466;
   reg _401467_401467 ; 
   reg __401467_401467;
   reg _401468_401468 ; 
   reg __401468_401468;
   reg _401469_401469 ; 
   reg __401469_401469;
   reg _401470_401470 ; 
   reg __401470_401470;
   reg _401471_401471 ; 
   reg __401471_401471;
   reg _401472_401472 ; 
   reg __401472_401472;
   reg _401473_401473 ; 
   reg __401473_401473;
   reg _401474_401474 ; 
   reg __401474_401474;
   reg _401475_401475 ; 
   reg __401475_401475;
   reg _401476_401476 ; 
   reg __401476_401476;
   reg _401477_401477 ; 
   reg __401477_401477;
   reg _401478_401478 ; 
   reg __401478_401478;
   reg _401479_401479 ; 
   reg __401479_401479;
   reg _401480_401480 ; 
   reg __401480_401480;
   reg _401481_401481 ; 
   reg __401481_401481;
   reg _401482_401482 ; 
   reg __401482_401482;
   reg _401483_401483 ; 
   reg __401483_401483;
   reg _401484_401484 ; 
   reg __401484_401484;
   reg _401485_401485 ; 
   reg __401485_401485;
   reg _401486_401486 ; 
   reg __401486_401486;
   reg _401487_401487 ; 
   reg __401487_401487;
   reg _401488_401488 ; 
   reg __401488_401488;
   reg _401489_401489 ; 
   reg __401489_401489;
   reg _401490_401490 ; 
   reg __401490_401490;
   reg _401491_401491 ; 
   reg __401491_401491;
   reg _401492_401492 ; 
   reg __401492_401492;
   reg _401493_401493 ; 
   reg __401493_401493;
   reg _401494_401494 ; 
   reg __401494_401494;
   reg _401495_401495 ; 
   reg __401495_401495;
   reg _401496_401496 ; 
   reg __401496_401496;
   reg _401497_401497 ; 
   reg __401497_401497;
   reg _401498_401498 ; 
   reg __401498_401498;
   reg _401499_401499 ; 
   reg __401499_401499;
   reg _401500_401500 ; 
   reg __401500_401500;
   reg _401501_401501 ; 
   reg __401501_401501;
   reg _401502_401502 ; 
   reg __401502_401502;
   reg _401503_401503 ; 
   reg __401503_401503;
   reg _401504_401504 ; 
   reg __401504_401504;
   reg _401505_401505 ; 
   reg __401505_401505;
   reg _401506_401506 ; 
   reg __401506_401506;
   reg _401507_401507 ; 
   reg __401507_401507;
   reg _401508_401508 ; 
   reg __401508_401508;
   reg _401509_401509 ; 
   reg __401509_401509;
   reg _401510_401510 ; 
   reg __401510_401510;
   reg _401511_401511 ; 
   reg __401511_401511;
   reg _401512_401512 ; 
   reg __401512_401512;
   reg _401513_401513 ; 
   reg __401513_401513;
   reg _401514_401514 ; 
   reg __401514_401514;
   reg _401515_401515 ; 
   reg __401515_401515;
   reg _401516_401516 ; 
   reg __401516_401516;
   reg _401517_401517 ; 
   reg __401517_401517;
   reg _401518_401518 ; 
   reg __401518_401518;
   reg _401519_401519 ; 
   reg __401519_401519;
   reg _401520_401520 ; 
   reg __401520_401520;
   reg _401521_401521 ; 
   reg __401521_401521;
   reg _401522_401522 ; 
   reg __401522_401522;
   reg _401523_401523 ; 
   reg __401523_401523;
   reg _401524_401524 ; 
   reg __401524_401524;
   reg _401525_401525 ; 
   reg __401525_401525;
   reg _401526_401526 ; 
   reg __401526_401526;
   reg _401527_401527 ; 
   reg __401527_401527;
   reg _401528_401528 ; 
   reg __401528_401528;
   reg _401529_401529 ; 
   reg __401529_401529;
   reg _401530_401530 ; 
   reg __401530_401530;
   reg _401531_401531 ; 
   reg __401531_401531;
   reg _401532_401532 ; 
   reg __401532_401532;
   reg _401533_401533 ; 
   reg __401533_401533;
   reg _401534_401534 ; 
   reg __401534_401534;
   reg _401535_401535 ; 
   reg __401535_401535;
   reg _401536_401536 ; 
   reg __401536_401536;
   reg _401537_401537 ; 
   reg __401537_401537;
   reg _401538_401538 ; 
   reg __401538_401538;
   reg _401539_401539 ; 
   reg __401539_401539;
   reg _401540_401540 ; 
   reg __401540_401540;
   reg _401541_401541 ; 
   reg __401541_401541;
   reg _401542_401542 ; 
   reg __401542_401542;
   reg _401543_401543 ; 
   reg __401543_401543;
   reg _401544_401544 ; 
   reg __401544_401544;
   reg _401545_401545 ; 
   reg __401545_401545;
   reg _401546_401546 ; 
   reg __401546_401546;
   reg _401547_401547 ; 
   reg __401547_401547;
   reg _401548_401548 ; 
   reg __401548_401548;
   reg _401549_401549 ; 
   reg __401549_401549;
   reg _401550_401550 ; 
   reg __401550_401550;
   reg _401551_401551 ; 
   reg __401551_401551;
   reg _401552_401552 ; 
   reg __401552_401552;
   reg _401553_401553 ; 
   reg __401553_401553;
   reg _401554_401554 ; 
   reg __401554_401554;
   reg _401555_401555 ; 
   reg __401555_401555;
   reg _401556_401556 ; 
   reg __401556_401556;
   reg _401557_401557 ; 
   reg __401557_401557;
   reg _401558_401558 ; 
   reg __401558_401558;
   reg _401559_401559 ; 
   reg __401559_401559;
   reg _401560_401560 ; 
   reg __401560_401560;
   reg _401561_401561 ; 
   reg __401561_401561;
   reg _401562_401562 ; 
   reg __401562_401562;
   reg _401563_401563 ; 
   reg __401563_401563;
   reg _401564_401564 ; 
   reg __401564_401564;
   reg _401565_401565 ; 
   reg __401565_401565;
   reg _401566_401566 ; 
   reg __401566_401566;
   reg _401567_401567 ; 
   reg __401567_401567;
   reg _401568_401568 ; 
   reg __401568_401568;
   reg _401569_401569 ; 
   reg __401569_401569;
   reg _401570_401570 ; 
   reg __401570_401570;
   reg _401571_401571 ; 
   reg __401571_401571;
   reg _401572_401572 ; 
   reg __401572_401572;
   reg _401573_401573 ; 
   reg __401573_401573;
   reg _401574_401574 ; 
   reg __401574_401574;
   reg _401575_401575 ; 
   reg __401575_401575;
   reg _401576_401576 ; 
   reg __401576_401576;
   reg _401577_401577 ; 
   reg __401577_401577;
   reg _401578_401578 ; 
   reg __401578_401578;
   reg _401579_401579 ; 
   reg __401579_401579;
   reg _401580_401580 ; 
   reg __401580_401580;
   reg _401581_401581 ; 
   reg __401581_401581;
   reg _401582_401582 ; 
   reg __401582_401582;
   reg _401583_401583 ; 
   reg __401583_401583;
   reg _401584_401584 ; 
   reg __401584_401584;
   reg _401585_401585 ; 
   reg __401585_401585;
   reg _401586_401586 ; 
   reg __401586_401586;
   reg _401587_401587 ; 
   reg __401587_401587;
   reg _401588_401588 ; 
   reg __401588_401588;
   reg _401589_401589 ; 
   reg __401589_401589;
   reg _401590_401590 ; 
   reg __401590_401590;
   reg _401591_401591 ; 
   reg __401591_401591;
   reg _401592_401592 ; 
   reg __401592_401592;
   reg _401593_401593 ; 
   reg __401593_401593;
   reg _401594_401594 ; 
   reg __401594_401594;
   reg _401595_401595 ; 
   reg __401595_401595;
   reg _401596_401596 ; 
   reg __401596_401596;
   reg _401597_401597 ; 
   reg __401597_401597;
   reg _401598_401598 ; 
   reg __401598_401598;
   reg _401599_401599 ; 
   reg __401599_401599;
   reg _401600_401600 ; 
   reg __401600_401600;
   reg _401601_401601 ; 
   reg __401601_401601;
   reg _401602_401602 ; 
   reg __401602_401602;
   reg _401603_401603 ; 
   reg __401603_401603;
   reg _401604_401604 ; 
   reg __401604_401604;
   reg _401605_401605 ; 
   reg __401605_401605;
   reg _401606_401606 ; 
   reg __401606_401606;
   reg _401607_401607 ; 
   reg __401607_401607;
   reg _401608_401608 ; 
   reg __401608_401608;
   reg _401609_401609 ; 
   reg __401609_401609;
   reg _401610_401610 ; 
   reg __401610_401610;
   reg _401611_401611 ; 
   reg __401611_401611;
   reg _401612_401612 ; 
   reg __401612_401612;
   reg _401613_401613 ; 
   reg __401613_401613;
   reg _401614_401614 ; 
   reg __401614_401614;
   reg _401615_401615 ; 
   reg __401615_401615;
   reg _401616_401616 ; 
   reg __401616_401616;
   reg _401617_401617 ; 
   reg __401617_401617;
   reg _401618_401618 ; 
   reg __401618_401618;
   reg _401619_401619 ; 
   reg __401619_401619;
   reg _401620_401620 ; 
   reg __401620_401620;
   reg _401621_401621 ; 
   reg __401621_401621;
   reg _401622_401622 ; 
   reg __401622_401622;
   reg _401623_401623 ; 
   reg __401623_401623;
   reg _401624_401624 ; 
   reg __401624_401624;
   reg _401625_401625 ; 
   reg __401625_401625;
   reg _401626_401626 ; 
   reg __401626_401626;
   reg _401627_401627 ; 
   reg __401627_401627;
   reg _401628_401628 ; 
   reg __401628_401628;
   reg _401629_401629 ; 
   reg __401629_401629;
   reg _401630_401630 ; 
   reg __401630_401630;
   reg _401631_401631 ; 
   reg __401631_401631;
   reg _401632_401632 ; 
   reg __401632_401632;
   reg _401633_401633 ; 
   reg __401633_401633;
   reg _401634_401634 ; 
   reg __401634_401634;
   reg _401635_401635 ; 
   reg __401635_401635;
   reg _401636_401636 ; 
   reg __401636_401636;
   reg _401637_401637 ; 
   reg __401637_401637;
   reg _401638_401638 ; 
   reg __401638_401638;
   reg _401639_401639 ; 
   reg __401639_401639;
   reg _401640_401640 ; 
   reg __401640_401640;
   reg _401641_401641 ; 
   reg __401641_401641;
   reg _401642_401642 ; 
   reg __401642_401642;
   reg _401643_401643 ; 
   reg __401643_401643;
   reg _401644_401644 ; 
   reg __401644_401644;
   reg _401645_401645 ; 
   reg __401645_401645;
   reg _401646_401646 ; 
   reg __401646_401646;
   reg _401647_401647 ; 
   reg __401647_401647;
   reg _401648_401648 ; 
   reg __401648_401648;
   reg _401649_401649 ; 
   reg __401649_401649;
   reg _401650_401650 ; 
   reg __401650_401650;
   reg _401651_401651 ; 
   reg __401651_401651;
   reg _401652_401652 ; 
   reg __401652_401652;
   reg _401653_401653 ; 
   reg __401653_401653;
   reg _401654_401654 ; 
   reg __401654_401654;
   reg _401655_401655 ; 
   reg __401655_401655;
   reg _401656_401656 ; 
   reg __401656_401656;
   reg _401657_401657 ; 
   reg __401657_401657;
   reg _401658_401658 ; 
   reg __401658_401658;
   reg _401659_401659 ; 
   reg __401659_401659;
   reg _401660_401660 ; 
   reg __401660_401660;
   reg _401661_401661 ; 
   reg __401661_401661;
   reg _401662_401662 ; 
   reg __401662_401662;
   reg _401663_401663 ; 
   reg __401663_401663;
   reg _401664_401664 ; 
   reg __401664_401664;
   reg _401665_401665 ; 
   reg __401665_401665;
   reg _401666_401666 ; 
   reg __401666_401666;
   reg _401667_401667 ; 
   reg __401667_401667;
   reg _401668_401668 ; 
   reg __401668_401668;
   reg _401669_401669 ; 
   reg __401669_401669;
   reg _401670_401670 ; 
   reg __401670_401670;
   reg _401671_401671 ; 
   reg __401671_401671;
   reg _401672_401672 ; 
   reg __401672_401672;
   reg _401673_401673 ; 
   reg __401673_401673;
   reg _401674_401674 ; 
   reg __401674_401674;
   reg _401675_401675 ; 
   reg __401675_401675;
   reg _401676_401676 ; 
   reg __401676_401676;
   reg _401677_401677 ; 
   reg __401677_401677;
   reg _401678_401678 ; 
   reg __401678_401678;
   reg _401679_401679 ; 
   reg __401679_401679;
   reg _401680_401680 ; 
   reg __401680_401680;
   reg _401681_401681 ; 
   reg __401681_401681;
   reg _401682_401682 ; 
   reg __401682_401682;
   reg _401683_401683 ; 
   reg __401683_401683;
   reg _401684_401684 ; 
   reg __401684_401684;
   reg _401685_401685 ; 
   reg __401685_401685;
   reg _401686_401686 ; 
   reg __401686_401686;
   reg _401687_401687 ; 
   reg __401687_401687;
   reg _401688_401688 ; 
   reg __401688_401688;
   reg _401689_401689 ; 
   reg __401689_401689;
   reg _401690_401690 ; 
   reg __401690_401690;
   reg _401691_401691 ; 
   reg __401691_401691;
   reg _401692_401692 ; 
   reg __401692_401692;
   reg _401693_401693 ; 
   reg __401693_401693;
   reg _401694_401694 ; 
   reg __401694_401694;
   reg _401695_401695 ; 
   reg __401695_401695;
   reg _401696_401696 ; 
   reg __401696_401696;
   reg _401697_401697 ; 
   reg __401697_401697;
   reg _401698_401698 ; 
   reg __401698_401698;
   reg _401699_401699 ; 
   reg __401699_401699;
   reg _401700_401700 ; 
   reg __401700_401700;
   reg _401701_401701 ; 
   reg __401701_401701;
   reg _401702_401702 ; 
   reg __401702_401702;
   reg _401703_401703 ; 
   reg __401703_401703;
   reg _401704_401704 ; 
   reg __401704_401704;
   reg _401705_401705 ; 
   reg __401705_401705;
   reg _401706_401706 ; 
   reg __401706_401706;
   reg _401707_401707 ; 
   reg __401707_401707;
   reg _401708_401708 ; 
   reg __401708_401708;
   reg _401709_401709 ; 
   reg __401709_401709;
   reg _401710_401710 ; 
   reg __401710_401710;
   reg _401711_401711 ; 
   reg __401711_401711;
   reg _401712_401712 ; 
   reg __401712_401712;
   reg _401713_401713 ; 
   reg __401713_401713;
   reg _401714_401714 ; 
   reg __401714_401714;
   reg _401715_401715 ; 
   reg __401715_401715;
   reg _401716_401716 ; 
   reg __401716_401716;
   reg _401717_401717 ; 
   reg __401717_401717;
   reg _401718_401718 ; 
   reg __401718_401718;
   reg _401719_401719 ; 
   reg __401719_401719;
   reg _401720_401720 ; 
   reg __401720_401720;
   reg _401721_401721 ; 
   reg __401721_401721;
   reg _401722_401722 ; 
   reg __401722_401722;
   reg _401723_401723 ; 
   reg __401723_401723;
   reg _401724_401724 ; 
   reg __401724_401724;
   reg _401725_401725 ; 
   reg __401725_401725;
   reg _401726_401726 ; 
   reg __401726_401726;
   reg _401727_401727 ; 
   reg __401727_401727;
   reg _401728_401728 ; 
   reg __401728_401728;
   reg _401729_401729 ; 
   reg __401729_401729;
   reg _401730_401730 ; 
   reg __401730_401730;
   reg _401731_401731 ; 
   reg __401731_401731;
   reg _401732_401732 ; 
   reg __401732_401732;
   reg _401733_401733 ; 
   reg __401733_401733;
   reg _401734_401734 ; 
   reg __401734_401734;
   reg _401735_401735 ; 
   reg __401735_401735;
   reg _401736_401736 ; 
   reg __401736_401736;
   reg _401737_401737 ; 
   reg __401737_401737;
   reg _401738_401738 ; 
   reg __401738_401738;
   reg _401739_401739 ; 
   reg __401739_401739;
   reg _401740_401740 ; 
   reg __401740_401740;
   reg _401741_401741 ; 
   reg __401741_401741;
   reg _401742_401742 ; 
   reg __401742_401742;
   reg _401743_401743 ; 
   reg __401743_401743;
   reg _401744_401744 ; 
   reg __401744_401744;
   reg _401745_401745 ; 
   reg __401745_401745;
   reg _401746_401746 ; 
   reg __401746_401746;
   reg _401747_401747 ; 
   reg __401747_401747;
   reg _401748_401748 ; 
   reg __401748_401748;
   reg _401749_401749 ; 
   reg __401749_401749;
   reg _401750_401750 ; 
   reg __401750_401750;
   reg _401751_401751 ; 
   reg __401751_401751;
   reg _401752_401752 ; 
   reg __401752_401752;
   reg _401753_401753 ; 
   reg __401753_401753;
   reg _401754_401754 ; 
   reg __401754_401754;
   reg _401755_401755 ; 
   reg __401755_401755;
   reg _401756_401756 ; 
   reg __401756_401756;
   reg _401757_401757 ; 
   reg __401757_401757;
   reg _401758_401758 ; 
   reg __401758_401758;
   reg _401759_401759 ; 
   reg __401759_401759;
   reg _401760_401760 ; 
   reg __401760_401760;
   reg _401761_401761 ; 
   reg __401761_401761;
   reg _401762_401762 ; 
   reg __401762_401762;
   reg _401763_401763 ; 
   reg __401763_401763;
   reg _401764_401764 ; 
   reg __401764_401764;
   reg _401765_401765 ; 
   reg __401765_401765;
   reg _401766_401766 ; 
   reg __401766_401766;
   reg _401767_401767 ; 
   reg __401767_401767;
   reg _401768_401768 ; 
   reg __401768_401768;
   reg _401769_401769 ; 
   reg __401769_401769;
   reg _401770_401770 ; 
   reg __401770_401770;
   reg _401771_401771 ; 
   reg __401771_401771;
   reg _401772_401772 ; 
   reg __401772_401772;
   reg _401773_401773 ; 
   reg __401773_401773;
   reg _401774_401774 ; 
   reg __401774_401774;
   reg _401775_401775 ; 
   reg __401775_401775;
   reg _401776_401776 ; 
   reg __401776_401776;
   reg _401777_401777 ; 
   reg __401777_401777;
   reg _401778_401778 ; 
   reg __401778_401778;
   reg _401779_401779 ; 
   reg __401779_401779;
   reg _401780_401780 ; 
   reg __401780_401780;
   reg _401781_401781 ; 
   reg __401781_401781;
   reg _401782_401782 ; 
   reg __401782_401782;
   reg _401783_401783 ; 
   reg __401783_401783;
   reg _401784_401784 ; 
   reg __401784_401784;
   reg _401785_401785 ; 
   reg __401785_401785;
   reg _401786_401786 ; 
   reg __401786_401786;
   reg _401787_401787 ; 
   reg __401787_401787;
   reg _401788_401788 ; 
   reg __401788_401788;
   reg _401789_401789 ; 
   reg __401789_401789;
   reg _401790_401790 ; 
   reg __401790_401790;
   reg _401791_401791 ; 
   reg __401791_401791;
   reg _401792_401792 ; 
   reg __401792_401792;
   reg _401793_401793 ; 
   reg __401793_401793;
   reg _401794_401794 ; 
   reg __401794_401794;
   reg _401795_401795 ; 
   reg __401795_401795;
   reg _401796_401796 ; 
   reg __401796_401796;
   reg _401797_401797 ; 
   reg __401797_401797;
   reg _401798_401798 ; 
   reg __401798_401798;
   reg _401799_401799 ; 
   reg __401799_401799;
   reg _401800_401800 ; 
   reg __401800_401800;
   reg _401801_401801 ; 
   reg __401801_401801;
   reg _401802_401802 ; 
   reg __401802_401802;
   reg _401803_401803 ; 
   reg __401803_401803;
   reg _401804_401804 ; 
   reg __401804_401804;
   reg _401805_401805 ; 
   reg __401805_401805;
   reg _401806_401806 ; 
   reg __401806_401806;
   reg _401807_401807 ; 
   reg __401807_401807;
   reg _401808_401808 ; 
   reg __401808_401808;
   reg _401809_401809 ; 
   reg __401809_401809;
   reg _401810_401810 ; 
   reg __401810_401810;
   reg _401811_401811 ; 
   reg __401811_401811;
   reg _401812_401812 ; 
   reg __401812_401812;
   reg _401813_401813 ; 
   reg __401813_401813;
   reg _401814_401814 ; 
   reg __401814_401814;
   reg _401815_401815 ; 
   reg __401815_401815;
   reg _401816_401816 ; 
   reg __401816_401816;
   reg _401817_401817 ; 
   reg __401817_401817;
   reg _401818_401818 ; 
   reg __401818_401818;
   reg _401819_401819 ; 
   reg __401819_401819;
   reg _401820_401820 ; 
   reg __401820_401820;
   reg _401821_401821 ; 
   reg __401821_401821;
   reg _401822_401822 ; 
   reg __401822_401822;
   reg _401823_401823 ; 
   reg __401823_401823;
   reg _401824_401824 ; 
   reg __401824_401824;
   reg _401825_401825 ; 
   reg __401825_401825;
   reg _401826_401826 ; 
   reg __401826_401826;
   reg _401827_401827 ; 
   reg __401827_401827;
   reg _401828_401828 ; 
   reg __401828_401828;
   reg _401829_401829 ; 
   reg __401829_401829;
   reg _401830_401830 ; 
   reg __401830_401830;
   reg _401831_401831 ; 
   reg __401831_401831;
   reg _401832_401832 ; 
   reg __401832_401832;
   reg _401833_401833 ; 
   reg __401833_401833;
   reg _401834_401834 ; 
   reg __401834_401834;
   reg _401835_401835 ; 
   reg __401835_401835;
   reg _401836_401836 ; 
   reg __401836_401836;
   reg _401837_401837 ; 
   reg __401837_401837;
   reg _401838_401838 ; 
   reg __401838_401838;
   reg _401839_401839 ; 
   reg __401839_401839;
   reg _401840_401840 ; 
   reg __401840_401840;
   reg _401841_401841 ; 
   reg __401841_401841;
   reg _401842_401842 ; 
   reg __401842_401842;
   reg _401843_401843 ; 
   reg __401843_401843;
   reg _401844_401844 ; 
   reg __401844_401844;
   reg _401845_401845 ; 
   reg __401845_401845;
   reg _401846_401846 ; 
   reg __401846_401846;
   reg _401847_401847 ; 
   reg __401847_401847;
   reg _401848_401848 ; 
   reg __401848_401848;
   reg _401849_401849 ; 
   reg __401849_401849;
   reg _401850_401850 ; 
   reg __401850_401850;
   reg _401851_401851 ; 
   reg __401851_401851;
   reg _401852_401852 ; 
   reg __401852_401852;
   reg _401853_401853 ; 
   reg __401853_401853;
   reg _401854_401854 ; 
   reg __401854_401854;
   reg _401855_401855 ; 
   reg __401855_401855;
   reg _401856_401856 ; 
   reg __401856_401856;
   reg _401857_401857 ; 
   reg __401857_401857;
   reg _401858_401858 ; 
   reg __401858_401858;
   reg _401859_401859 ; 
   reg __401859_401859;
   reg _401860_401860 ; 
   reg __401860_401860;
   reg _401861_401861 ; 
   reg __401861_401861;
   reg _401862_401862 ; 
   reg __401862_401862;
   reg _401863_401863 ; 
   reg __401863_401863;
   reg _401864_401864 ; 
   reg __401864_401864;
   reg _401865_401865 ; 
   reg __401865_401865;
   reg _401866_401866 ; 
   reg __401866_401866;
   reg _401867_401867 ; 
   reg __401867_401867;
   reg _401868_401868 ; 
   reg __401868_401868;
   reg _401869_401869 ; 
   reg __401869_401869;
   reg _401870_401870 ; 
   reg __401870_401870;
   reg _401871_401871 ; 
   reg __401871_401871;
   reg _401872_401872 ; 
   reg __401872_401872;
   reg _401873_401873 ; 
   reg __401873_401873;
   reg _401874_401874 ; 
   reg __401874_401874;
   reg _401875_401875 ; 
   reg __401875_401875;
   reg _401876_401876 ; 
   reg __401876_401876;
   reg _401877_401877 ; 
   reg __401877_401877;
   reg _401878_401878 ; 
   reg __401878_401878;
   reg _401879_401879 ; 
   reg __401879_401879;
   reg _401880_401880 ; 
   reg __401880_401880;
   reg _401881_401881 ; 
   reg __401881_401881;
   reg _401882_401882 ; 
   reg __401882_401882;
   reg _401883_401883 ; 
   reg __401883_401883;
   reg _401884_401884 ; 
   reg __401884_401884;
   reg _401885_401885 ; 
   reg __401885_401885;
   reg _401886_401886 ; 
   reg __401886_401886;
   reg _401887_401887 ; 
   reg __401887_401887;
   reg _401888_401888 ; 
   reg __401888_401888;
   reg _401889_401889 ; 
   reg __401889_401889;
   reg _401890_401890 ; 
   reg __401890_401890;
   reg _401891_401891 ; 
   reg __401891_401891;
   reg _401892_401892 ; 
   reg __401892_401892;
   reg _401893_401893 ; 
   reg __401893_401893;
   reg _401894_401894 ; 
   reg __401894_401894;
   reg _401895_401895 ; 
   reg __401895_401895;
   reg _401896_401896 ; 
   reg __401896_401896;
   reg _401897_401897 ; 
   reg __401897_401897;
   reg _401898_401898 ; 
   reg __401898_401898;
   reg _401899_401899 ; 
   reg __401899_401899;
   reg _401900_401900 ; 
   reg __401900_401900;
   reg _401901_401901 ; 
   reg __401901_401901;
   reg _401902_401902 ; 
   reg __401902_401902;
   reg _401903_401903 ; 
   reg __401903_401903;
   reg _401904_401904 ; 
   reg __401904_401904;
   reg _401905_401905 ; 
   reg __401905_401905;
   reg _401906_401906 ; 
   reg __401906_401906;
   reg _401907_401907 ; 
   reg __401907_401907;
   reg _401908_401908 ; 
   reg __401908_401908;
   reg _401909_401909 ; 
   reg __401909_401909;
   reg _401910_401910 ; 
   reg __401910_401910;
   reg _401911_401911 ; 
   reg __401911_401911;
   reg _401912_401912 ; 
   reg __401912_401912;
   reg _401913_401913 ; 
   reg __401913_401913;
   reg _401914_401914 ; 
   reg __401914_401914;
   reg _401915_401915 ; 
   reg __401915_401915;
   reg _401916_401916 ; 
   reg __401916_401916;
   reg _401917_401917 ; 
   reg __401917_401917;
   reg _401918_401918 ; 
   reg __401918_401918;
   reg _401919_401919 ; 
   reg __401919_401919;
   reg _401920_401920 ; 
   reg __401920_401920;
   reg _401921_401921 ; 
   reg __401921_401921;
   reg _401922_401922 ; 
   reg __401922_401922;
   reg _401923_401923 ; 
   reg __401923_401923;
   reg _401924_401924 ; 
   reg __401924_401924;
   reg _401925_401925 ; 
   reg __401925_401925;
   reg _401926_401926 ; 
   reg __401926_401926;
   reg _401927_401927 ; 
   reg __401927_401927;
   reg _401928_401928 ; 
   reg __401928_401928;
   reg _401929_401929 ; 
   reg __401929_401929;
   reg _401930_401930 ; 
   reg __401930_401930;
   reg _401931_401931 ; 
   reg __401931_401931;
   reg _401932_401932 ; 
   reg __401932_401932;
   reg _401933_401933 ; 
   reg __401933_401933;
   reg _401934_401934 ; 
   reg __401934_401934;
   reg _401935_401935 ; 
   reg __401935_401935;
   reg _401936_401936 ; 
   reg __401936_401936;
   reg _401937_401937 ; 
   reg __401937_401937;
   reg _401938_401938 ; 
   reg __401938_401938;
   reg _401939_401939 ; 
   reg __401939_401939;
   reg _401940_401940 ; 
   reg __401940_401940;
   reg _401941_401941 ; 
   reg __401941_401941;
   reg _401942_401942 ; 
   reg __401942_401942;
   reg _401943_401943 ; 
   reg __401943_401943;
   reg _401944_401944 ; 
   reg __401944_401944;
   reg _401945_401945 ; 
   reg __401945_401945;
   reg _401946_401946 ; 
   reg __401946_401946;
   reg _401947_401947 ; 
   reg __401947_401947;
   reg _401948_401948 ; 
   reg __401948_401948;
   reg _401949_401949 ; 
   reg __401949_401949;
   reg _401950_401950 ; 
   reg __401950_401950;
   reg _401951_401951 ; 
   reg __401951_401951;
   reg _401952_401952 ; 
   reg __401952_401952;
   reg _401953_401953 ; 
   reg __401953_401953;
   reg _401954_401954 ; 
   reg __401954_401954;
   reg _401955_401955 ; 
   reg __401955_401955;
   reg _401956_401956 ; 
   reg __401956_401956;
   reg _401957_401957 ; 
   reg __401957_401957;
   reg _401958_401958 ; 
   reg __401958_401958;
   reg _401959_401959 ; 
   reg __401959_401959;
   reg _401960_401960 ; 
   reg __401960_401960;
   reg _401961_401961 ; 
   reg __401961_401961;
   reg _401962_401962 ; 
   reg __401962_401962;
   reg _401963_401963 ; 
   reg __401963_401963;
   reg _401964_401964 ; 
   reg __401964_401964;
   reg _401965_401965 ; 
   reg __401965_401965;
   reg _401966_401966 ; 
   reg __401966_401966;
   reg _401967_401967 ; 
   reg __401967_401967;
   reg _401968_401968 ; 
   reg __401968_401968;
   reg _401969_401969 ; 
   reg __401969_401969;
   reg _401970_401970 ; 
   reg __401970_401970;
   reg _401971_401971 ; 
   reg __401971_401971;
   reg _401972_401972 ; 
   reg __401972_401972;
   reg _401973_401973 ; 
   reg __401973_401973;
   reg _401974_401974 ; 
   reg __401974_401974;
   reg _401975_401975 ; 
   reg __401975_401975;
   reg _401976_401976 ; 
   reg __401976_401976;
   reg _401977_401977 ; 
   reg __401977_401977;
   reg _401978_401978 ; 
   reg __401978_401978;
   reg _401979_401979 ; 
   reg __401979_401979;
   reg _401980_401980 ; 
   reg __401980_401980;
   reg _401981_401981 ; 
   reg __401981_401981;
   reg _401982_401982 ; 
   reg __401982_401982;
   reg _401983_401983 ; 
   reg __401983_401983;
   reg _401984_401984 ; 
   reg __401984_401984;
   reg _401985_401985 ; 
   reg __401985_401985;
   reg _401986_401986 ; 
   reg __401986_401986;
   reg _401987_401987 ; 
   reg __401987_401987;
   reg _401988_401988 ; 
   reg __401988_401988;
   reg _401989_401989 ; 
   reg __401989_401989;
   reg _401990_401990 ; 
   reg __401990_401990;
   reg _401991_401991 ; 
   reg __401991_401991;
   reg _401992_401992 ; 
   reg __401992_401992;
   reg _401993_401993 ; 
   reg __401993_401993;
   reg _401994_401994 ; 
   reg __401994_401994;
   reg _401995_401995 ; 
   reg __401995_401995;
   reg _401996_401996 ; 
   reg __401996_401996;
   reg _401997_401997 ; 
   reg __401997_401997;
   reg _401998_401998 ; 
   reg __401998_401998;
   reg _401999_401999 ; 
   reg __401999_401999;
   reg _402000_402000 ; 
   reg __402000_402000;
   reg _402001_402001 ; 
   reg __402001_402001;
   reg _402002_402002 ; 
   reg __402002_402002;
   reg _402003_402003 ; 
   reg __402003_402003;
   reg _402004_402004 ; 
   reg __402004_402004;
   reg _402005_402005 ; 
   reg __402005_402005;
   reg _402006_402006 ; 
   reg __402006_402006;
   reg _402007_402007 ; 
   reg __402007_402007;
   reg _402008_402008 ; 
   reg __402008_402008;
   reg _402009_402009 ; 
   reg __402009_402009;
   reg _402010_402010 ; 
   reg __402010_402010;
   reg _402011_402011 ; 
   reg __402011_402011;
   reg _402012_402012 ; 
   reg __402012_402012;
   reg _402013_402013 ; 
   reg __402013_402013;
   reg _402014_402014 ; 
   reg __402014_402014;
   reg _402015_402015 ; 
   reg __402015_402015;
   reg _402016_402016 ; 
   reg __402016_402016;
   reg _402017_402017 ; 
   reg __402017_402017;
   reg _402018_402018 ; 
   reg __402018_402018;
   reg _402019_402019 ; 
   reg __402019_402019;
   reg _402020_402020 ; 
   reg __402020_402020;
   reg _402021_402021 ; 
   reg __402021_402021;
   reg _402022_402022 ; 
   reg __402022_402022;
   reg _402023_402023 ; 
   reg __402023_402023;
   reg _402024_402024 ; 
   reg __402024_402024;
   reg _402025_402025 ; 
   reg __402025_402025;
   reg _402026_402026 ; 
   reg __402026_402026;
   reg _402027_402027 ; 
   reg __402027_402027;
   reg _402028_402028 ; 
   reg __402028_402028;
   reg _402029_402029 ; 
   reg __402029_402029;
   reg _402030_402030 ; 
   reg __402030_402030;
   reg _402031_402031 ; 
   reg __402031_402031;
   reg _402032_402032 ; 
   reg __402032_402032;
   reg _402033_402033 ; 
   reg __402033_402033;
   reg _402034_402034 ; 
   reg __402034_402034;
   reg _402035_402035 ; 
   reg __402035_402035;
   reg _402036_402036 ; 
   reg __402036_402036;
   reg _402037_402037 ; 
   reg __402037_402037;
   reg _402038_402038 ; 
   reg __402038_402038;
   reg _402039_402039 ; 
   reg __402039_402039;
   reg _402040_402040 ; 
   reg __402040_402040;
   reg _402041_402041 ; 
   reg __402041_402041;
   reg _402042_402042 ; 
   reg __402042_402042;
   reg _402043_402043 ; 
   reg __402043_402043;
   reg _402044_402044 ; 
   reg __402044_402044;
   reg _402045_402045 ; 
   reg __402045_402045;
   reg _402046_402046 ; 
   reg __402046_402046;
   reg _402047_402047 ; 
   reg __402047_402047;
   reg _402048_402048 ; 
   reg __402048_402048;
   reg _402049_402049 ; 
   reg __402049_402049;
   reg _402050_402050 ; 
   reg __402050_402050;
   reg _402051_402051 ; 
   reg __402051_402051;
   reg _402052_402052 ; 
   reg __402052_402052;
   reg _402053_402053 ; 
   reg __402053_402053;
   reg _402054_402054 ; 
   reg __402054_402054;
   reg _402055_402055 ; 
   reg __402055_402055;
   reg _402056_402056 ; 
   reg __402056_402056;
   reg _402057_402057 ; 
   reg __402057_402057;
   reg _402058_402058 ; 
   reg __402058_402058;
   reg _402059_402059 ; 
   reg __402059_402059;
   reg _402060_402060 ; 
   reg __402060_402060;
   reg _402061_402061 ; 
   reg __402061_402061;
   reg _402062_402062 ; 
   reg __402062_402062;
   reg _402063_402063 ; 
   reg __402063_402063;
   reg _402064_402064 ; 
   reg __402064_402064;
   reg _402065_402065 ; 
   reg __402065_402065;
   reg _402066_402066 ; 
   reg __402066_402066;
   reg _402067_402067 ; 
   reg __402067_402067;
   reg _402068_402068 ; 
   reg __402068_402068;
   reg _402069_402069 ; 
   reg __402069_402069;
   reg _402070_402070 ; 
   reg __402070_402070;
   reg _402071_402071 ; 
   reg __402071_402071;
   reg _402072_402072 ; 
   reg __402072_402072;
   reg _402073_402073 ; 
   reg __402073_402073;
   reg _402074_402074 ; 
   reg __402074_402074;
   reg _402075_402075 ; 
   reg __402075_402075;
   reg _402076_402076 ; 
   reg __402076_402076;
   reg _402077_402077 ; 
   reg __402077_402077;
   reg _402078_402078 ; 
   reg __402078_402078;
   reg _402079_402079 ; 
   reg __402079_402079;
   reg _402080_402080 ; 
   reg __402080_402080;
   reg _402081_402081 ; 
   reg __402081_402081;
   reg _402082_402082 ; 
   reg __402082_402082;
   reg _402083_402083 ; 
   reg __402083_402083;
   reg _402084_402084 ; 
   reg __402084_402084;
   reg _402085_402085 ; 
   reg __402085_402085;
   reg _402086_402086 ; 
   reg __402086_402086;
   reg _402087_402087 ; 
   reg __402087_402087;
   reg _402088_402088 ; 
   reg __402088_402088;
   reg _402089_402089 ; 
   reg __402089_402089;
   reg _402090_402090 ; 
   reg __402090_402090;
   reg _402091_402091 ; 
   reg __402091_402091;
   reg _402092_402092 ; 
   reg __402092_402092;
   reg _402093_402093 ; 
   reg __402093_402093;
   reg _402094_402094 ; 
   reg __402094_402094;
   reg _402095_402095 ; 
   reg __402095_402095;
   reg _402096_402096 ; 
   reg __402096_402096;
   reg _402097_402097 ; 
   reg __402097_402097;
   reg _402098_402098 ; 
   reg __402098_402098;
   reg _402099_402099 ; 
   reg __402099_402099;
   reg _402100_402100 ; 
   reg __402100_402100;
   reg _402101_402101 ; 
   reg __402101_402101;
   reg _402102_402102 ; 
   reg __402102_402102;
   reg _402103_402103 ; 
   reg __402103_402103;
   reg _402104_402104 ; 
   reg __402104_402104;
   reg _402105_402105 ; 
   reg __402105_402105;
   reg _402106_402106 ; 
   reg __402106_402106;
   reg _402107_402107 ; 
   reg __402107_402107;
   reg _402108_402108 ; 
   reg __402108_402108;
   reg _402109_402109 ; 
   reg __402109_402109;
   reg _402110_402110 ; 
   reg __402110_402110;
   reg _402111_402111 ; 
   reg __402111_402111;
   reg _402112_402112 ; 
   reg __402112_402112;
   reg _402113_402113 ; 
   reg __402113_402113;
   reg _402114_402114 ; 
   reg __402114_402114;
   reg _402115_402115 ; 
   reg __402115_402115;
   reg _402116_402116 ; 
   reg __402116_402116;
   reg _402117_402117 ; 
   reg __402117_402117;
   reg _402118_402118 ; 
   reg __402118_402118;
   reg _402119_402119 ; 
   reg __402119_402119;
   reg _402120_402120 ; 
   reg __402120_402120;
   reg _402121_402121 ; 
   reg __402121_402121;
   reg _402122_402122 ; 
   reg __402122_402122;
   reg _402123_402123 ; 
   reg __402123_402123;
   reg _402124_402124 ; 
   reg __402124_402124;
   reg _402125_402125 ; 
   reg __402125_402125;
   reg _402126_402126 ; 
   reg __402126_402126;
   reg _402127_402127 ; 
   reg __402127_402127;
   reg _402128_402128 ; 
   reg __402128_402128;
   reg _402129_402129 ; 
   reg __402129_402129;
   reg _402130_402130 ; 
   reg __402130_402130;
   reg _402131_402131 ; 
   reg __402131_402131;
   reg _402132_402132 ; 
   reg __402132_402132;
   reg _402133_402133 ; 
   reg __402133_402133;
   reg _402134_402134 ; 
   reg __402134_402134;
   reg _402135_402135 ; 
   reg __402135_402135;
   reg _402136_402136 ; 
   reg __402136_402136;
   reg _402137_402137 ; 
   reg __402137_402137;
   reg _402138_402138 ; 
   reg __402138_402138;
   reg _402139_402139 ; 
   reg __402139_402139;
   reg _402140_402140 ; 
   reg __402140_402140;
   reg _402141_402141 ; 
   reg __402141_402141;
   reg _402142_402142 ; 
   reg __402142_402142;
   reg _402143_402143 ; 
   reg __402143_402143;
   reg _402144_402144 ; 
   reg __402144_402144;
   reg _402145_402145 ; 
   reg __402145_402145;
   reg _402146_402146 ; 
   reg __402146_402146;
   reg _402147_402147 ; 
   reg __402147_402147;
   reg _402148_402148 ; 
   reg __402148_402148;
   reg _402149_402149 ; 
   reg __402149_402149;
   reg _402150_402150 ; 
   reg __402150_402150;
   reg _402151_402151 ; 
   reg __402151_402151;
   reg _402152_402152 ; 
   reg __402152_402152;
   reg _402153_402153 ; 
   reg __402153_402153;
   reg _402154_402154 ; 
   reg __402154_402154;
   reg _402155_402155 ; 
   reg __402155_402155;
   reg _402156_402156 ; 
   reg __402156_402156;
   reg _402157_402157 ; 
   reg __402157_402157;
   reg _402158_402158 ; 
   reg __402158_402158;
   reg _402159_402159 ; 
   reg __402159_402159;
   reg _402160_402160 ; 
   reg __402160_402160;
   reg _402161_402161 ; 
   reg __402161_402161;
   reg _402162_402162 ; 
   reg __402162_402162;
   reg _402163_402163 ; 
   reg __402163_402163;
   reg _402164_402164 ; 
   reg __402164_402164;
   reg _402165_402165 ; 
   reg __402165_402165;
   reg _402166_402166 ; 
   reg __402166_402166;
   reg _402167_402167 ; 
   reg __402167_402167;
   reg _402168_402168 ; 
   reg __402168_402168;
   reg _402169_402169 ; 
   reg __402169_402169;
   reg _402170_402170 ; 
   reg __402170_402170;
   reg _402171_402171 ; 
   reg __402171_402171;
   reg _402172_402172 ; 
   reg __402172_402172;
   reg _402173_402173 ; 
   reg __402173_402173;
   reg _402174_402174 ; 
   reg __402174_402174;
   reg _402175_402175 ; 
   reg __402175_402175;
   reg _402176_402176 ; 
   reg __402176_402176;
   reg _402177_402177 ; 
   reg __402177_402177;
   reg _402178_402178 ; 
   reg __402178_402178;
   reg _402179_402179 ; 
   reg __402179_402179;
   reg _402180_402180 ; 
   reg __402180_402180;
   reg _402181_402181 ; 
   reg __402181_402181;
   reg _402182_402182 ; 
   reg __402182_402182;
   reg _402183_402183 ; 
   reg __402183_402183;
   reg _402184_402184 ; 
   reg __402184_402184;
   reg _402185_402185 ; 
   reg __402185_402185;
   reg _402186_402186 ; 
   reg __402186_402186;
   reg _402187_402187 ; 
   reg __402187_402187;
   reg _402188_402188 ; 
   reg __402188_402188;
   reg _402189_402189 ; 
   reg __402189_402189;
   reg _402190_402190 ; 
   reg __402190_402190;
   reg _402191_402191 ; 
   reg __402191_402191;
   reg _402192_402192 ; 
   reg __402192_402192;
   reg _402193_402193 ; 
   reg __402193_402193;
   reg _402194_402194 ; 
   reg __402194_402194;
   reg _402195_402195 ; 
   reg __402195_402195;
   reg _402196_402196 ; 
   reg __402196_402196;
   reg _402197_402197 ; 
   reg __402197_402197;
   reg _402198_402198 ; 
   reg __402198_402198;
   reg _402199_402199 ; 
   reg __402199_402199;
   reg _402200_402200 ; 
   reg __402200_402200;
   reg _402201_402201 ; 
   reg __402201_402201;
   reg _402202_402202 ; 
   reg __402202_402202;
   reg _402203_402203 ; 
   reg __402203_402203;
   reg _402204_402204 ; 
   reg __402204_402204;
   reg _402205_402205 ; 
   reg __402205_402205;
   reg _402206_402206 ; 
   reg __402206_402206;
   reg _402207_402207 ; 
   reg __402207_402207;
   reg _402208_402208 ; 
   reg __402208_402208;
   reg _402209_402209 ; 
   reg __402209_402209;
   reg _402210_402210 ; 
   reg __402210_402210;
   reg _402211_402211 ; 
   reg __402211_402211;
   reg _402212_402212 ; 
   reg __402212_402212;
   reg _402213_402213 ; 
   reg __402213_402213;
   reg _402214_402214 ; 
   reg __402214_402214;
   reg _402215_402215 ; 
   reg __402215_402215;
   reg _402216_402216 ; 
   reg __402216_402216;
   reg _402217_402217 ; 
   reg __402217_402217;
   reg _402218_402218 ; 
   reg __402218_402218;
   reg _402219_402219 ; 
   reg __402219_402219;
   reg _402220_402220 ; 
   reg __402220_402220;
   reg _402221_402221 ; 
   reg __402221_402221;
   reg _402222_402222 ; 
   reg __402222_402222;
   reg _402223_402223 ; 
   reg __402223_402223;
   reg _402224_402224 ; 
   reg __402224_402224;
   reg _402225_402225 ; 
   reg __402225_402225;
   reg _402226_402226 ; 
   reg __402226_402226;
   reg _402227_402227 ; 
   reg __402227_402227;
   reg _402228_402228 ; 
   reg __402228_402228;
   reg _402229_402229 ; 
   reg __402229_402229;
   reg _402230_402230 ; 
   reg __402230_402230;
   reg _402231_402231 ; 
   reg __402231_402231;
   reg _402232_402232 ; 
   reg __402232_402232;
   reg _402233_402233 ; 
   reg __402233_402233;
   reg _402234_402234 ; 
   reg __402234_402234;
   reg _402235_402235 ; 
   reg __402235_402235;
   reg _402236_402236 ; 
   reg __402236_402236;
   reg _402237_402237 ; 
   reg __402237_402237;
   reg _402238_402238 ; 
   reg __402238_402238;
   reg _402239_402239 ; 
   reg __402239_402239;
   reg _402240_402240 ; 
   reg __402240_402240;
   reg _402241_402241 ; 
   reg __402241_402241;
   reg _402242_402242 ; 
   reg __402242_402242;
   reg _402243_402243 ; 
   reg __402243_402243;
   reg _402244_402244 ; 
   reg __402244_402244;
   reg _402245_402245 ; 
   reg __402245_402245;
   reg _402246_402246 ; 
   reg __402246_402246;
   reg _402247_402247 ; 
   reg __402247_402247;
   reg _402248_402248 ; 
   reg __402248_402248;
   reg _402249_402249 ; 
   reg __402249_402249;
   reg _402250_402250 ; 
   reg __402250_402250;
   reg _402251_402251 ; 
   reg __402251_402251;
   reg _402252_402252 ; 
   reg __402252_402252;
   reg _402253_402253 ; 
   reg __402253_402253;
   reg _402254_402254 ; 
   reg __402254_402254;
   reg _402255_402255 ; 
   reg __402255_402255;
   reg _402256_402256 ; 
   reg __402256_402256;
   reg _402257_402257 ; 
   reg __402257_402257;
   reg _402258_402258 ; 
   reg __402258_402258;
   reg _402259_402259 ; 
   reg __402259_402259;
   reg _402260_402260 ; 
   reg __402260_402260;
   reg _402261_402261 ; 
   reg __402261_402261;
   reg _402262_402262 ; 
   reg __402262_402262;
   reg _402263_402263 ; 
   reg __402263_402263;
   reg _402264_402264 ; 
   reg __402264_402264;
   reg _402265_402265 ; 
   reg __402265_402265;
   reg _402266_402266 ; 
   reg __402266_402266;
   reg _402267_402267 ; 
   reg __402267_402267;
   reg _402268_402268 ; 
   reg __402268_402268;
   reg _402269_402269 ; 
   reg __402269_402269;
   reg _402270_402270 ; 
   reg __402270_402270;
   reg _402271_402271 ; 
   reg __402271_402271;
   reg _402272_402272 ; 
   reg __402272_402272;
   reg _402273_402273 ; 
   reg __402273_402273;
   reg _402274_402274 ; 
   reg __402274_402274;
   reg _402275_402275 ; 
   reg __402275_402275;
   reg _402276_402276 ; 
   reg __402276_402276;
   reg _402277_402277 ; 
   reg __402277_402277;
   reg _402278_402278 ; 
   reg __402278_402278;
   reg _402279_402279 ; 
   reg __402279_402279;
   reg _402280_402280 ; 
   reg __402280_402280;
   reg _402281_402281 ; 
   reg __402281_402281;
   reg _402282_402282 ; 
   reg __402282_402282;
   reg _402283_402283 ; 
   reg __402283_402283;
   reg _402284_402284 ; 
   reg __402284_402284;
   reg _402285_402285 ; 
   reg __402285_402285;
   reg _402286_402286 ; 
   reg __402286_402286;
   reg _402287_402287 ; 
   reg __402287_402287;
   reg _402288_402288 ; 
   reg __402288_402288;
   reg _402289_402289 ; 
   reg __402289_402289;
   reg _402290_402290 ; 
   reg __402290_402290;
   reg _402291_402291 ; 
   reg __402291_402291;
   reg _402292_402292 ; 
   reg __402292_402292;
   reg _402293_402293 ; 
   reg __402293_402293;
   reg _402294_402294 ; 
   reg __402294_402294;
   reg _402295_402295 ; 
   reg __402295_402295;
   reg _402296_402296 ; 
   reg __402296_402296;
   reg _402297_402297 ; 
   reg __402297_402297;
   reg _402298_402298 ; 
   reg __402298_402298;
   reg _402299_402299 ; 
   reg __402299_402299;
   reg _402300_402300 ; 
   reg __402300_402300;
   reg _402301_402301 ; 
   reg __402301_402301;
   reg _402302_402302 ; 
   reg __402302_402302;
   reg _402303_402303 ; 
   reg __402303_402303;
   reg _402304_402304 ; 
   reg __402304_402304;
   reg _402305_402305 ; 
   reg __402305_402305;
   reg _402306_402306 ; 
   reg __402306_402306;
   reg _402307_402307 ; 
   reg __402307_402307;
   reg _402308_402308 ; 
   reg __402308_402308;
   reg _402309_402309 ; 
   reg __402309_402309;
   reg _402310_402310 ; 
   reg __402310_402310;
   reg _402311_402311 ; 
   reg __402311_402311;
   reg _402312_402312 ; 
   reg __402312_402312;
   reg _402313_402313 ; 
   reg __402313_402313;
   reg _402314_402314 ; 
   reg __402314_402314;
   reg _402315_402315 ; 
   reg __402315_402315;
   reg _402316_402316 ; 
   reg __402316_402316;
   reg _402317_402317 ; 
   reg __402317_402317;
   reg _402318_402318 ; 
   reg __402318_402318;
   reg _402319_402319 ; 
   reg __402319_402319;
   reg _402320_402320 ; 
   reg __402320_402320;
   reg _402321_402321 ; 
   reg __402321_402321;
   reg _402322_402322 ; 
   reg __402322_402322;
   reg _402323_402323 ; 
   reg __402323_402323;
   reg _402324_402324 ; 
   reg __402324_402324;
   reg _402325_402325 ; 
   reg __402325_402325;
   reg _402326_402326 ; 
   reg __402326_402326;
   reg _402327_402327 ; 
   reg __402327_402327;
   reg _402328_402328 ; 
   reg __402328_402328;
   reg _402329_402329 ; 
   reg __402329_402329;
   reg _402330_402330 ; 
   reg __402330_402330;
   reg _402331_402331 ; 
   reg __402331_402331;
   reg _402332_402332 ; 
   reg __402332_402332;
   reg _402333_402333 ; 
   reg __402333_402333;
   reg _402334_402334 ; 
   reg __402334_402334;
   reg _402335_402335 ; 
   reg __402335_402335;
   reg _402336_402336 ; 
   reg __402336_402336;
   reg _402337_402337 ; 
   reg __402337_402337;
   reg _402338_402338 ; 
   reg __402338_402338;
   reg _402339_402339 ; 
   reg __402339_402339;
   reg _402340_402340 ; 
   reg __402340_402340;
   reg _402341_402341 ; 
   reg __402341_402341;
   reg _402342_402342 ; 
   reg __402342_402342;
   reg _402343_402343 ; 
   reg __402343_402343;
   reg _402344_402344 ; 
   reg __402344_402344;
   reg _402345_402345 ; 
   reg __402345_402345;
   reg _402346_402346 ; 
   reg __402346_402346;
   reg _402347_402347 ; 
   reg __402347_402347;
   reg _402348_402348 ; 
   reg __402348_402348;
   reg _402349_402349 ; 
   reg __402349_402349;
   reg _402350_402350 ; 
   reg __402350_402350;
   reg _402351_402351 ; 
   reg __402351_402351;
   reg _402352_402352 ; 
   reg __402352_402352;
   reg _402353_402353 ; 
   reg __402353_402353;
   reg _402354_402354 ; 
   reg __402354_402354;
   reg _402355_402355 ; 
   reg __402355_402355;
   reg _402356_402356 ; 
   reg __402356_402356;
   reg _402357_402357 ; 
   reg __402357_402357;
   reg _402358_402358 ; 
   reg __402358_402358;
   reg _402359_402359 ; 
   reg __402359_402359;
   reg _402360_402360 ; 
   reg __402360_402360;
   reg _402361_402361 ; 
   reg __402361_402361;
   reg _402362_402362 ; 
   reg __402362_402362;
   reg _402363_402363 ; 
   reg __402363_402363;
   reg _402364_402364 ; 
   reg __402364_402364;
   reg _402365_402365 ; 
   reg __402365_402365;
   reg _402366_402366 ; 
   reg __402366_402366;
   reg _402367_402367 ; 
   reg __402367_402367;
   reg _402368_402368 ; 
   reg __402368_402368;
   reg _402369_402369 ; 
   reg __402369_402369;
   reg _402370_402370 ; 
   reg __402370_402370;
   reg _402371_402371 ; 
   reg __402371_402371;
   reg _402372_402372 ; 
   reg __402372_402372;
   reg _402373_402373 ; 
   reg __402373_402373;
   reg _402374_402374 ; 
   reg __402374_402374;
   reg _402375_402375 ; 
   reg __402375_402375;
   reg _402376_402376 ; 
   reg __402376_402376;
   reg _402377_402377 ; 
   reg __402377_402377;
   reg _402378_402378 ; 
   reg __402378_402378;
   reg _402379_402379 ; 
   reg __402379_402379;
   reg _402380_402380 ; 
   reg __402380_402380;
   reg _402381_402381 ; 
   reg __402381_402381;
   reg _402382_402382 ; 
   reg __402382_402382;
   reg _402383_402383 ; 
   reg __402383_402383;
   reg _402384_402384 ; 
   reg __402384_402384;
   reg _402385_402385 ; 
   reg __402385_402385;
   reg _402386_402386 ; 
   reg __402386_402386;
   reg _402387_402387 ; 
   reg __402387_402387;
   reg _402388_402388 ; 
   reg __402388_402388;
   reg _402389_402389 ; 
   reg __402389_402389;
   reg _402390_402390 ; 
   reg __402390_402390;
   reg _402391_402391 ; 
   reg __402391_402391;
   reg _402392_402392 ; 
   reg __402392_402392;
   reg _402393_402393 ; 
   reg __402393_402393;
   reg _402394_402394 ; 
   reg __402394_402394;
   reg _402395_402395 ; 
   reg __402395_402395;
   reg _402396_402396 ; 
   reg __402396_402396;
   reg _402397_402397 ; 
   reg __402397_402397;
   reg _402398_402398 ; 
   reg __402398_402398;
   reg _402399_402399 ; 
   reg __402399_402399;
   reg _402400_402400 ; 
   reg __402400_402400;
   reg _402401_402401 ; 
   reg __402401_402401;
   reg _402402_402402 ; 
   reg __402402_402402;
   reg _402403_402403 ; 
   reg __402403_402403;
   reg _402404_402404 ; 
   reg __402404_402404;
   reg _402405_402405 ; 
   reg __402405_402405;
   reg _402406_402406 ; 
   reg __402406_402406;
   reg _402407_402407 ; 
   reg __402407_402407;
   reg _402408_402408 ; 
   reg __402408_402408;
   reg _402409_402409 ; 
   reg __402409_402409;
   reg _402410_402410 ; 
   reg __402410_402410;
   reg _402411_402411 ; 
   reg __402411_402411;
   reg _402412_402412 ; 
   reg __402412_402412;
   reg _402413_402413 ; 
   reg __402413_402413;
   reg _402414_402414 ; 
   reg __402414_402414;
   reg _402415_402415 ; 
   reg __402415_402415;
   reg _402416_402416 ; 
   reg __402416_402416;
   reg _402417_402417 ; 
   reg __402417_402417;
   reg _402418_402418 ; 
   reg __402418_402418;
   reg _402419_402419 ; 
   reg __402419_402419;
   reg _402420_402420 ; 
   reg __402420_402420;
   reg _402421_402421 ; 
   reg __402421_402421;
   reg _402422_402422 ; 
   reg __402422_402422;
   reg _402423_402423 ; 
   reg __402423_402423;
   reg _402424_402424 ; 
   reg __402424_402424;
   reg _402425_402425 ; 
   reg __402425_402425;
   reg _402426_402426 ; 
   reg __402426_402426;
   reg _402427_402427 ; 
   reg __402427_402427;
   reg _402428_402428 ; 
   reg __402428_402428;
   reg _402429_402429 ; 
   reg __402429_402429;
   reg _402430_402430 ; 
   reg __402430_402430;
   reg _402431_402431 ; 
   reg __402431_402431;
   reg _402432_402432 ; 
   reg __402432_402432;
   reg _402433_402433 ; 
   reg __402433_402433;
   reg _402434_402434 ; 
   reg __402434_402434;
   reg _402435_402435 ; 
   reg __402435_402435;
   reg _402436_402436 ; 
   reg __402436_402436;
   reg _402437_402437 ; 
   reg __402437_402437;
   reg _402438_402438 ; 
   reg __402438_402438;
   reg _402439_402439 ; 
   reg __402439_402439;
   reg _402440_402440 ; 
   reg __402440_402440;
   reg _402441_402441 ; 
   reg __402441_402441;
   reg _402442_402442 ; 
   reg __402442_402442;
   reg _402443_402443 ; 
   reg __402443_402443;
   reg _402444_402444 ; 
   reg __402444_402444;
   reg _402445_402445 ; 
   reg __402445_402445;
   reg _402446_402446 ; 
   reg __402446_402446;
   reg _402447_402447 ; 
   reg __402447_402447;
   reg _402448_402448 ; 
   reg __402448_402448;
   reg _402449_402449 ; 
   reg __402449_402449;
   reg _402450_402450 ; 
   reg __402450_402450;
   reg _402451_402451 ; 
   reg __402451_402451;
   reg _402452_402452 ; 
   reg __402452_402452;
   reg _402453_402453 ; 
   reg __402453_402453;
   reg _402454_402454 ; 
   reg __402454_402454;
   reg _402455_402455 ; 
   reg __402455_402455;
   reg _402456_402456 ; 
   reg __402456_402456;
   reg _402457_402457 ; 
   reg __402457_402457;
   reg _402458_402458 ; 
   reg __402458_402458;
   reg _402459_402459 ; 
   reg __402459_402459;
   reg _402460_402460 ; 
   reg __402460_402460;
   reg _402461_402461 ; 
   reg __402461_402461;
   reg _402462_402462 ; 
   reg __402462_402462;
   reg _402463_402463 ; 
   reg __402463_402463;
   reg _402464_402464 ; 
   reg __402464_402464;
   reg _402465_402465 ; 
   reg __402465_402465;
   reg _402466_402466 ; 
   reg __402466_402466;
   reg _402467_402467 ; 
   reg __402467_402467;
   reg _402468_402468 ; 
   reg __402468_402468;
   reg _402469_402469 ; 
   reg __402469_402469;
   reg _402470_402470 ; 
   reg __402470_402470;
   reg _402471_402471 ; 
   reg __402471_402471;
   reg _402472_402472 ; 
   reg __402472_402472;
   reg _402473_402473 ; 
   reg __402473_402473;
   reg _402474_402474 ; 
   reg __402474_402474;
   reg _402475_402475 ; 
   reg __402475_402475;
   reg _402476_402476 ; 
   reg __402476_402476;
   reg _402477_402477 ; 
   reg __402477_402477;
   reg _402478_402478 ; 
   reg __402478_402478;
   reg _402479_402479 ; 
   reg __402479_402479;
   reg _402480_402480 ; 
   reg __402480_402480;
   reg _402481_402481 ; 
   reg __402481_402481;
   reg _402482_402482 ; 
   reg __402482_402482;
   reg _402483_402483 ; 
   reg __402483_402483;
   reg _402484_402484 ; 
   reg __402484_402484;
   reg _402485_402485 ; 
   reg __402485_402485;
   reg _402486_402486 ; 
   reg __402486_402486;
   reg _402487_402487 ; 
   reg __402487_402487;
   reg _402488_402488 ; 
   reg __402488_402488;
   reg _402489_402489 ; 
   reg __402489_402489;
   reg _402490_402490 ; 
   reg __402490_402490;
   reg _402491_402491 ; 
   reg __402491_402491;
   reg _402492_402492 ; 
   reg __402492_402492;
   reg _402493_402493 ; 
   reg __402493_402493;
   reg _402494_402494 ; 
   reg __402494_402494;
   reg _402495_402495 ; 
   reg __402495_402495;
   reg _402496_402496 ; 
   reg __402496_402496;
   reg _402497_402497 ; 
   reg __402497_402497;
   reg _402498_402498 ; 
   reg __402498_402498;
   reg _402499_402499 ; 
   reg __402499_402499;
   reg _402500_402500 ; 
   reg __402500_402500;
   reg _402501_402501 ; 
   reg __402501_402501;
   reg _402502_402502 ; 
   reg __402502_402502;
   reg _402503_402503 ; 
   reg __402503_402503;
   reg _402504_402504 ; 
   reg __402504_402504;
   reg _402505_402505 ; 
   reg __402505_402505;
   reg _402506_402506 ; 
   reg __402506_402506;
   reg _402507_402507 ; 
   reg __402507_402507;
   reg _402508_402508 ; 
   reg __402508_402508;
   reg _402509_402509 ; 
   reg __402509_402509;
   reg _402510_402510 ; 
   reg __402510_402510;
   reg _402511_402511 ; 
   reg __402511_402511;
   reg _402512_402512 ; 
   reg __402512_402512;
   reg _402513_402513 ; 
   reg __402513_402513;
   reg _402514_402514 ; 
   reg __402514_402514;
   reg _402515_402515 ; 
   reg __402515_402515;
   reg _402516_402516 ; 
   reg __402516_402516;
   reg _402517_402517 ; 
   reg __402517_402517;
   reg _402518_402518 ; 
   reg __402518_402518;
   reg _402519_402519 ; 
   reg __402519_402519;
   reg _402520_402520 ; 
   reg __402520_402520;
   reg _402521_402521 ; 
   reg __402521_402521;
   reg _402522_402522 ; 
   reg __402522_402522;
   reg _402523_402523 ; 
   reg __402523_402523;
   reg _402524_402524 ; 
   reg __402524_402524;
   reg _402525_402525 ; 
   reg __402525_402525;
   reg _402526_402526 ; 
   reg __402526_402526;
   reg _402527_402527 ; 
   reg __402527_402527;
   reg _402528_402528 ; 
   reg __402528_402528;
   reg _402529_402529 ; 
   reg __402529_402529;
   reg _402530_402530 ; 
   reg __402530_402530;
   reg _402531_402531 ; 
   reg __402531_402531;
   reg _402532_402532 ; 
   reg __402532_402532;
   reg _402533_402533 ; 
   reg __402533_402533;
   reg _402534_402534 ; 
   reg __402534_402534;
   reg _402535_402535 ; 
   reg __402535_402535;
   reg _402536_402536 ; 
   reg __402536_402536;
   reg _402537_402537 ; 
   reg __402537_402537;
   reg _402538_402538 ; 
   reg __402538_402538;
   reg _402539_402539 ; 
   reg __402539_402539;
   reg _402540_402540 ; 
   reg __402540_402540;
   reg _402541_402541 ; 
   reg __402541_402541;
   reg _402542_402542 ; 
   reg __402542_402542;
   reg _402543_402543 ; 
   reg __402543_402543;
   reg _402544_402544 ; 
   reg __402544_402544;
   reg _402545_402545 ; 
   reg __402545_402545;
   reg _402546_402546 ; 
   reg __402546_402546;
   reg _402547_402547 ; 
   reg __402547_402547;
   reg _402548_402548 ; 
   reg __402548_402548;
   reg _402549_402549 ; 
   reg __402549_402549;
   reg _402550_402550 ; 
   reg __402550_402550;
   reg _402551_402551 ; 
   reg __402551_402551;
   reg _402552_402552 ; 
   reg __402552_402552;
   reg _402553_402553 ; 
   reg __402553_402553;
   reg _402554_402554 ; 
   reg __402554_402554;
   reg _402555_402555 ; 
   reg __402555_402555;
   reg _402556_402556 ; 
   reg __402556_402556;
   reg _402557_402557 ; 
   reg __402557_402557;
   reg _402558_402558 ; 
   reg __402558_402558;
   reg _402559_402559 ; 
   reg __402559_402559;
   reg _402560_402560 ; 
   reg __402560_402560;
   reg _402561_402561 ; 
   reg __402561_402561;
   reg _402562_402562 ; 
   reg __402562_402562;
   reg _402563_402563 ; 
   reg __402563_402563;
   reg _402564_402564 ; 
   reg __402564_402564;
   reg _402565_402565 ; 
   reg __402565_402565;
   reg _402566_402566 ; 
   reg __402566_402566;
   reg _402567_402567 ; 
   reg __402567_402567;
   reg _402568_402568 ; 
   reg __402568_402568;
   reg _402569_402569 ; 
   reg __402569_402569;
   reg _402570_402570 ; 
   reg __402570_402570;
   reg _402571_402571 ; 
   reg __402571_402571;
   reg _402572_402572 ; 
   reg __402572_402572;
   reg _402573_402573 ; 
   reg __402573_402573;
   reg _402574_402574 ; 
   reg __402574_402574;
   reg _402575_402575 ; 
   reg __402575_402575;
   reg _402576_402576 ; 
   reg __402576_402576;
   reg _402577_402577 ; 
   reg __402577_402577;
   reg _402578_402578 ; 
   reg __402578_402578;
   reg _402579_402579 ; 
   reg __402579_402579;
   reg _402580_402580 ; 
   reg __402580_402580;
   reg _402581_402581 ; 
   reg __402581_402581;
   reg _402582_402582 ; 
   reg __402582_402582;
   reg _402583_402583 ; 
   reg __402583_402583;
   reg _402584_402584 ; 
   reg __402584_402584;
   reg _402585_402585 ; 
   reg __402585_402585;
   reg _402586_402586 ; 
   reg __402586_402586;
   reg _402587_402587 ; 
   reg __402587_402587;
   reg _402588_402588 ; 
   reg __402588_402588;
   reg _402589_402589 ; 
   reg __402589_402589;
   reg _402590_402590 ; 
   reg __402590_402590;
   reg _402591_402591 ; 
   reg __402591_402591;
   reg _402592_402592 ; 
   reg __402592_402592;
   reg _402593_402593 ; 
   reg __402593_402593;
   reg _402594_402594 ; 
   reg __402594_402594;
   reg _402595_402595 ; 
   reg __402595_402595;
   reg _402596_402596 ; 
   reg __402596_402596;
   reg _402597_402597 ; 
   reg __402597_402597;
   reg _402598_402598 ; 
   reg __402598_402598;
   reg _402599_402599 ; 
   reg __402599_402599;
   reg _402600_402600 ; 
   reg __402600_402600;
   reg _402601_402601 ; 
   reg __402601_402601;
   reg _402602_402602 ; 
   reg __402602_402602;
   reg _402603_402603 ; 
   reg __402603_402603;
   reg _402604_402604 ; 
   reg __402604_402604;
   reg _402605_402605 ; 
   reg __402605_402605;
   reg _402606_402606 ; 
   reg __402606_402606;
   reg _402607_402607 ; 
   reg __402607_402607;
   reg _402608_402608 ; 
   reg __402608_402608;
   reg _402609_402609 ; 
   reg __402609_402609;
   reg _402610_402610 ; 
   reg __402610_402610;
   reg _402611_402611 ; 
   reg __402611_402611;
   reg _402612_402612 ; 
   reg __402612_402612;
   reg _402613_402613 ; 
   reg __402613_402613;
   reg _402614_402614 ; 
   reg __402614_402614;
   reg _402615_402615 ; 
   reg __402615_402615;
   reg _402616_402616 ; 
   reg __402616_402616;
   reg _402617_402617 ; 
   reg __402617_402617;
   reg _402618_402618 ; 
   reg __402618_402618;
   reg _402619_402619 ; 
   reg __402619_402619;
   reg _402620_402620 ; 
   reg __402620_402620;
   reg _402621_402621 ; 
   reg __402621_402621;
   reg _402622_402622 ; 
   reg __402622_402622;
   reg _402623_402623 ; 
   reg __402623_402623;
   reg _402624_402624 ; 
   reg __402624_402624;
   reg _402625_402625 ; 
   reg __402625_402625;
   reg _402626_402626 ; 
   reg __402626_402626;
   reg _402627_402627 ; 
   reg __402627_402627;
   reg _402628_402628 ; 
   reg __402628_402628;
   reg _402629_402629 ; 
   reg __402629_402629;
   reg _402630_402630 ; 
   reg __402630_402630;
   reg _402631_402631 ; 
   reg __402631_402631;
   reg _402632_402632 ; 
   reg __402632_402632;
   reg _402633_402633 ; 
   reg __402633_402633;
   reg _402634_402634 ; 
   reg __402634_402634;
   reg _402635_402635 ; 
   reg __402635_402635;
   reg _402636_402636 ; 
   reg __402636_402636;
   reg _402637_402637 ; 
   reg __402637_402637;
   reg _402638_402638 ; 
   reg __402638_402638;
   reg _402639_402639 ; 
   reg __402639_402639;
   reg _402640_402640 ; 
   reg __402640_402640;
   reg _402641_402641 ; 
   reg __402641_402641;
   reg _402642_402642 ; 
   reg __402642_402642;
   reg _402643_402643 ; 
   reg __402643_402643;
   reg _402644_402644 ; 
   reg __402644_402644;
   reg _402645_402645 ; 
   reg __402645_402645;
   reg _402646_402646 ; 
   reg __402646_402646;
   reg _402647_402647 ; 
   reg __402647_402647;
   reg _402648_402648 ; 
   reg __402648_402648;
   reg _402649_402649 ; 
   reg __402649_402649;
   reg _402650_402650 ; 
   reg __402650_402650;
   reg _402651_402651 ; 
   reg __402651_402651;
   reg _402652_402652 ; 
   reg __402652_402652;
   reg _402653_402653 ; 
   reg __402653_402653;
   reg _402654_402654 ; 
   reg __402654_402654;
   reg _402655_402655 ; 
   reg __402655_402655;
   reg _402656_402656 ; 
   reg __402656_402656;
   reg _402657_402657 ; 
   reg __402657_402657;
   reg _402658_402658 ; 
   reg __402658_402658;
   reg _402659_402659 ; 
   reg __402659_402659;
   reg _402660_402660 ; 
   reg __402660_402660;
   reg _402661_402661 ; 
   reg __402661_402661;
   reg _402662_402662 ; 
   reg __402662_402662;
   reg _402663_402663 ; 
   reg __402663_402663;
   reg _402664_402664 ; 
   reg __402664_402664;
   reg _402665_402665 ; 
   reg __402665_402665;
   reg _402666_402666 ; 
   reg __402666_402666;
   reg _402667_402667 ; 
   reg __402667_402667;
   reg _402668_402668 ; 
   reg __402668_402668;
   reg _402669_402669 ; 
   reg __402669_402669;
   reg _402670_402670 ; 
   reg __402670_402670;
   reg _402671_402671 ; 
   reg __402671_402671;
   reg _402672_402672 ; 
   reg __402672_402672;
   reg _402673_402673 ; 
   reg __402673_402673;
   reg _402674_402674 ; 
   reg __402674_402674;
   reg _402675_402675 ; 
   reg __402675_402675;
   reg _402676_402676 ; 
   reg __402676_402676;
   reg _402677_402677 ; 
   reg __402677_402677;
   reg _402678_402678 ; 
   reg __402678_402678;
   reg _402679_402679 ; 
   reg __402679_402679;
   reg _402680_402680 ; 
   reg __402680_402680;
   reg _402681_402681 ; 
   reg __402681_402681;
   reg _402682_402682 ; 
   reg __402682_402682;
   reg _402683_402683 ; 
   reg __402683_402683;
   reg _402684_402684 ; 
   reg __402684_402684;
   reg _402685_402685 ; 
   reg __402685_402685;
   reg _402686_402686 ; 
   reg __402686_402686;
   reg _402687_402687 ; 
   reg __402687_402687;
   reg _402688_402688 ; 
   reg __402688_402688;
   reg _402689_402689 ; 
   reg __402689_402689;
   reg _402690_402690 ; 
   reg __402690_402690;
   reg _402691_402691 ; 
   reg __402691_402691;
   reg _402692_402692 ; 
   reg __402692_402692;
   reg _402693_402693 ; 
   reg __402693_402693;
   reg _402694_402694 ; 
   reg __402694_402694;
   reg _402695_402695 ; 
   reg __402695_402695;
   reg _402696_402696 ; 
   reg __402696_402696;
   reg _402697_402697 ; 
   reg __402697_402697;
   reg _402698_402698 ; 
   reg __402698_402698;
   reg _402699_402699 ; 
   reg __402699_402699;
   reg _402700_402700 ; 
   reg __402700_402700;
   reg _402701_402701 ; 
   reg __402701_402701;
   reg _402702_402702 ; 
   reg __402702_402702;
   reg _402703_402703 ; 
   reg __402703_402703;
   reg _402704_402704 ; 
   reg __402704_402704;
   reg _402705_402705 ; 
   reg __402705_402705;
   reg _402706_402706 ; 
   reg __402706_402706;
   reg _402707_402707 ; 
   reg __402707_402707;
   reg _402708_402708 ; 
   reg __402708_402708;
   reg _402709_402709 ; 
   reg __402709_402709;
   reg _402710_402710 ; 
   reg __402710_402710;
   reg _402711_402711 ; 
   reg __402711_402711;
   reg _402712_402712 ; 
   reg __402712_402712;
   reg _402713_402713 ; 
   reg __402713_402713;
   reg _402714_402714 ; 
   reg __402714_402714;
   reg _402715_402715 ; 
   reg __402715_402715;
   reg _402716_402716 ; 
   reg __402716_402716;
   reg _402717_402717 ; 
   reg __402717_402717;
   reg _402718_402718 ; 
   reg __402718_402718;
   reg _402719_402719 ; 
   reg __402719_402719;
   reg _402720_402720 ; 
   reg __402720_402720;
   reg _402721_402721 ; 
   reg __402721_402721;
   reg _402722_402722 ; 
   reg __402722_402722;
   reg _402723_402723 ; 
   reg __402723_402723;
   reg _402724_402724 ; 
   reg __402724_402724;
   reg _402725_402725 ; 
   reg __402725_402725;
   reg _402726_402726 ; 
   reg __402726_402726;
   reg _402727_402727 ; 
   reg __402727_402727;
   reg _402728_402728 ; 
   reg __402728_402728;
   reg _402729_402729 ; 
   reg __402729_402729;
   reg _402730_402730 ; 
   reg __402730_402730;
   reg _402731_402731 ; 
   reg __402731_402731;
   reg _402732_402732 ; 
   reg __402732_402732;
   reg _402733_402733 ; 
   reg __402733_402733;
   reg _402734_402734 ; 
   reg __402734_402734;
   reg _402735_402735 ; 
   reg __402735_402735;
   reg _402736_402736 ; 
   reg __402736_402736;
   reg _402737_402737 ; 
   reg __402737_402737;
   reg _402738_402738 ; 
   reg __402738_402738;
   reg _402739_402739 ; 
   reg __402739_402739;
   reg _402740_402740 ; 
   reg __402740_402740;
   reg _402741_402741 ; 
   reg __402741_402741;
   reg _402742_402742 ; 
   reg __402742_402742;
   reg _402743_402743 ; 
   reg __402743_402743;
   reg _402744_402744 ; 
   reg __402744_402744;
   reg _402745_402745 ; 
   reg __402745_402745;
   reg _402746_402746 ; 
   reg __402746_402746;
   reg _402747_402747 ; 
   reg __402747_402747;
   reg _402748_402748 ; 
   reg __402748_402748;
   reg _402749_402749 ; 
   reg __402749_402749;
   reg _402750_402750 ; 
   reg __402750_402750;
   reg _402751_402751 ; 
   reg __402751_402751;
   reg _402752_402752 ; 
   reg __402752_402752;
   reg _402753_402753 ; 
   reg __402753_402753;
   reg _402754_402754 ; 
   reg __402754_402754;
   reg _402755_402755 ; 
   reg __402755_402755;
   reg _402756_402756 ; 
   reg __402756_402756;
   reg _402757_402757 ; 
   reg __402757_402757;
   reg _402758_402758 ; 
   reg __402758_402758;
   reg _402759_402759 ; 
   reg __402759_402759;
   reg _402760_402760 ; 
   reg __402760_402760;
   reg _402761_402761 ; 
   reg __402761_402761;
   reg _402762_402762 ; 
   reg __402762_402762;
   reg _402763_402763 ; 
   reg __402763_402763;
   reg _402764_402764 ; 
   reg __402764_402764;
   reg _402765_402765 ; 
   reg __402765_402765;
   reg _402766_402766 ; 
   reg __402766_402766;
   reg _402767_402767 ; 
   reg __402767_402767;
   reg _402768_402768 ; 
   reg __402768_402768;
   reg _402769_402769 ; 
   reg __402769_402769;
   reg _402770_402770 ; 
   reg __402770_402770;
   reg _402771_402771 ; 
   reg __402771_402771;
   reg _402772_402772 ; 
   reg __402772_402772;
   reg _402773_402773 ; 
   reg __402773_402773;
   reg _402774_402774 ; 
   reg __402774_402774;
   reg _402775_402775 ; 
   reg __402775_402775;
   reg _402776_402776 ; 
   reg __402776_402776;
   reg _402777_402777 ; 
   reg __402777_402777;
   reg _402778_402778 ; 
   reg __402778_402778;
   reg _402779_402779 ; 
   reg __402779_402779;
   reg _402780_402780 ; 
   reg __402780_402780;
   reg _402781_402781 ; 
   reg __402781_402781;
   reg _402782_402782 ; 
   reg __402782_402782;
   reg _402783_402783 ; 
   reg __402783_402783;
   reg _402784_402784 ; 
   reg __402784_402784;
   reg _402785_402785 ; 
   reg __402785_402785;
   reg _402786_402786 ; 
   reg __402786_402786;
   reg _402787_402787 ; 
   reg __402787_402787;
   reg _402788_402788 ; 
   reg __402788_402788;
   reg _402789_402789 ; 
   reg __402789_402789;
   reg _402790_402790 ; 
   reg __402790_402790;
   reg _402791_402791 ; 
   reg __402791_402791;
   reg _402792_402792 ; 
   reg __402792_402792;
   reg _402793_402793 ; 
   reg __402793_402793;
   reg _402794_402794 ; 
   reg __402794_402794;
   reg _402795_402795 ; 
   reg __402795_402795;
   reg _402796_402796 ; 
   reg __402796_402796;
   reg _402797_402797 ; 
   reg __402797_402797;
   reg _402798_402798 ; 
   reg __402798_402798;
   reg _402799_402799 ; 
   reg __402799_402799;
   reg _402800_402800 ; 
   reg __402800_402800;
   reg _402801_402801 ; 
   reg __402801_402801;
   reg _402802_402802 ; 
   reg __402802_402802;
   reg _402803_402803 ; 
   reg __402803_402803;
   reg _402804_402804 ; 
   reg __402804_402804;
   reg _402805_402805 ; 
   reg __402805_402805;
   reg _402806_402806 ; 
   reg __402806_402806;
   reg _402807_402807 ; 
   reg __402807_402807;
   reg _402808_402808 ; 
   reg __402808_402808;
   reg _402809_402809 ; 
   reg __402809_402809;
   reg _402810_402810 ; 
   reg __402810_402810;
   reg _402811_402811 ; 
   reg __402811_402811;
   reg _402812_402812 ; 
   reg __402812_402812;
   reg _402813_402813 ; 
   reg __402813_402813;
   reg _402814_402814 ; 
   reg __402814_402814;
   reg _402815_402815 ; 
   reg __402815_402815;
   reg _402816_402816 ; 
   reg __402816_402816;
   reg _402817_402817 ; 
   reg __402817_402817;
   reg _402818_402818 ; 
   reg __402818_402818;
   reg _402819_402819 ; 
   reg __402819_402819;
   reg _402820_402820 ; 
   reg __402820_402820;
   reg _402821_402821 ; 
   reg __402821_402821;
   reg _402822_402822 ; 
   reg __402822_402822;
   reg _402823_402823 ; 
   reg __402823_402823;
   reg _402824_402824 ; 
   reg __402824_402824;
   reg _402825_402825 ; 
   reg __402825_402825;
   reg _402826_402826 ; 
   reg __402826_402826;
   reg _402827_402827 ; 
   reg __402827_402827;
   reg _402828_402828 ; 
   reg __402828_402828;
   reg _402829_402829 ; 
   reg __402829_402829;
   reg _402830_402830 ; 
   reg __402830_402830;
   reg _402831_402831 ; 
   reg __402831_402831;
   reg _402832_402832 ; 
   reg __402832_402832;
   reg _402833_402833 ; 
   reg __402833_402833;
   reg _402834_402834 ; 
   reg __402834_402834;
   reg _402835_402835 ; 
   reg __402835_402835;
   reg _402836_402836 ; 
   reg __402836_402836;
   reg _402837_402837 ; 
   reg __402837_402837;
   reg _402838_402838 ; 
   reg __402838_402838;
   reg _402839_402839 ; 
   reg __402839_402839;
   reg _402840_402840 ; 
   reg __402840_402840;
   reg _402841_402841 ; 
   reg __402841_402841;
   reg _402842_402842 ; 
   reg __402842_402842;
   reg _402843_402843 ; 
   reg __402843_402843;
   reg _402844_402844 ; 
   reg __402844_402844;
   reg _402845_402845 ; 
   reg __402845_402845;
   reg _402846_402846 ; 
   reg __402846_402846;
   reg _402847_402847 ; 
   reg __402847_402847;
   reg _402848_402848 ; 
   reg __402848_402848;
   reg _402849_402849 ; 
   reg __402849_402849;
   reg _402850_402850 ; 
   reg __402850_402850;
   reg _402851_402851 ; 
   reg __402851_402851;
   reg _402852_402852 ; 
   reg __402852_402852;
   reg _402853_402853 ; 
   reg __402853_402853;
   reg _402854_402854 ; 
   reg __402854_402854;
   reg _402855_402855 ; 
   reg __402855_402855;
   reg _402856_402856 ; 
   reg __402856_402856;
   reg _402857_402857 ; 
   reg __402857_402857;
   reg _402858_402858 ; 
   reg __402858_402858;
   reg _402859_402859 ; 
   reg __402859_402859;
   reg _402860_402860 ; 
   reg __402860_402860;
   reg _402861_402861 ; 
   reg __402861_402861;
   reg _402862_402862 ; 
   reg __402862_402862;
   reg _402863_402863 ; 
   reg __402863_402863;
   reg _402864_402864 ; 
   reg __402864_402864;
   reg _402865_402865 ; 
   reg __402865_402865;
   reg _402866_402866 ; 
   reg __402866_402866;
   reg _402867_402867 ; 
   reg __402867_402867;
   reg _402868_402868 ; 
   reg __402868_402868;
   reg _402869_402869 ; 
   reg __402869_402869;
   reg _402870_402870 ; 
   reg __402870_402870;
   reg _402871_402871 ; 
   reg __402871_402871;
   reg _402872_402872 ; 
   reg __402872_402872;
   reg _402873_402873 ; 
   reg __402873_402873;
   reg _402874_402874 ; 
   reg __402874_402874;
   reg _402875_402875 ; 
   reg __402875_402875;
   reg _402876_402876 ; 
   reg __402876_402876;
   reg _402877_402877 ; 
   reg __402877_402877;
   reg _402878_402878 ; 
   reg __402878_402878;
   reg _402879_402879 ; 
   reg __402879_402879;
   reg _402880_402880 ; 
   reg __402880_402880;
   reg _402881_402881 ; 
   reg __402881_402881;
   reg _402882_402882 ; 
   reg __402882_402882;
   reg _402883_402883 ; 
   reg __402883_402883;
   reg _402884_402884 ; 
   reg __402884_402884;
   reg _402885_402885 ; 
   reg __402885_402885;
   reg _402886_402886 ; 
   reg __402886_402886;
   reg _402887_402887 ; 
   reg __402887_402887;
   reg _402888_402888 ; 
   reg __402888_402888;
   reg _402889_402889 ; 
   reg __402889_402889;
   reg _402890_402890 ; 
   reg __402890_402890;
   reg _402891_402891 ; 
   reg __402891_402891;
   reg _402892_402892 ; 
   reg __402892_402892;
   reg _402893_402893 ; 
   reg __402893_402893;
   reg _402894_402894 ; 
   reg __402894_402894;
   reg _402895_402895 ; 
   reg __402895_402895;
   reg _402896_402896 ; 
   reg __402896_402896;
   reg _402897_402897 ; 
   reg __402897_402897;
   reg _402898_402898 ; 
   reg __402898_402898;
   reg _402899_402899 ; 
   reg __402899_402899;
   reg _402900_402900 ; 
   reg __402900_402900;
   reg _402901_402901 ; 
   reg __402901_402901;
   reg _402902_402902 ; 
   reg __402902_402902;
   reg _402903_402903 ; 
   reg __402903_402903;
   reg _402904_402904 ; 
   reg __402904_402904;
   reg _402905_402905 ; 
   reg __402905_402905;
   reg _402906_402906 ; 
   reg __402906_402906;
   reg _402907_402907 ; 
   reg __402907_402907;
   reg _402908_402908 ; 
   reg __402908_402908;
   reg _402909_402909 ; 
   reg __402909_402909;
   reg _402910_402910 ; 
   reg __402910_402910;
   reg _402911_402911 ; 
   reg __402911_402911;
   reg _402912_402912 ; 
   reg __402912_402912;
   reg _402913_402913 ; 
   reg __402913_402913;
   reg _402914_402914 ; 
   reg __402914_402914;
   reg _402915_402915 ; 
   reg __402915_402915;
   reg _402916_402916 ; 
   reg __402916_402916;
   reg _402917_402917 ; 
   reg __402917_402917;
   reg _402918_402918 ; 
   reg __402918_402918;
   reg _402919_402919 ; 
   reg __402919_402919;
   reg _402920_402920 ; 
   reg __402920_402920;
   reg _402921_402921 ; 
   reg __402921_402921;
   reg _402922_402922 ; 
   reg __402922_402922;
   reg _402923_402923 ; 
   reg __402923_402923;
   reg _402924_402924 ; 
   reg __402924_402924;
   reg _402925_402925 ; 
   reg __402925_402925;
   reg _402926_402926 ; 
   reg __402926_402926;
   reg _402927_402927 ; 
   reg __402927_402927;
   reg _402928_402928 ; 
   reg __402928_402928;
   reg _402929_402929 ; 
   reg __402929_402929;
   reg _402930_402930 ; 
   reg __402930_402930;
   reg _402931_402931 ; 
   reg __402931_402931;
   reg _402932_402932 ; 
   reg __402932_402932;
   reg _402933_402933 ; 
   reg __402933_402933;
   reg _402934_402934 ; 
   reg __402934_402934;
   reg _402935_402935 ; 
   reg __402935_402935;
   reg _402936_402936 ; 
   reg __402936_402936;
   reg _402937_402937 ; 
   reg __402937_402937;
   reg _402938_402938 ; 
   reg __402938_402938;
   reg _402939_402939 ; 
   reg __402939_402939;
   reg _402940_402940 ; 
   reg __402940_402940;
   reg _402941_402941 ; 
   reg __402941_402941;
   reg _402942_402942 ; 
   reg __402942_402942;
   reg _402943_402943 ; 
   reg __402943_402943;
   reg _402944_402944 ; 
   reg __402944_402944;
   reg _402945_402945 ; 
   reg __402945_402945;
   reg _402946_402946 ; 
   reg __402946_402946;
   reg _402947_402947 ; 
   reg __402947_402947;
   reg _402948_402948 ; 
   reg __402948_402948;
   reg _402949_402949 ; 
   reg __402949_402949;
   reg _402950_402950 ; 
   reg __402950_402950;
   reg _402951_402951 ; 
   reg __402951_402951;
   reg _402952_402952 ; 
   reg __402952_402952;
   reg _402953_402953 ; 
   reg __402953_402953;
   reg _402954_402954 ; 
   reg __402954_402954;
   reg _402955_402955 ; 
   reg __402955_402955;
   reg _402956_402956 ; 
   reg __402956_402956;
   reg _402957_402957 ; 
   reg __402957_402957;
   reg _402958_402958 ; 
   reg __402958_402958;
   reg _402959_402959 ; 
   reg __402959_402959;
   reg _402960_402960 ; 
   reg __402960_402960;
   reg _402961_402961 ; 
   reg __402961_402961;
   reg _402962_402962 ; 
   reg __402962_402962;
   reg _402963_402963 ; 
   reg __402963_402963;
   reg _402964_402964 ; 
   reg __402964_402964;
   reg _402965_402965 ; 
   reg __402965_402965;
   reg _402966_402966 ; 
   reg __402966_402966;
   reg _402967_402967 ; 
   reg __402967_402967;
   reg _402968_402968 ; 
   reg __402968_402968;
   reg _402969_402969 ; 
   reg __402969_402969;
   reg _402970_402970 ; 
   reg __402970_402970;
   reg _402971_402971 ; 
   reg __402971_402971;
   reg _402972_402972 ; 
   reg __402972_402972;
   reg _402973_402973 ; 
   reg __402973_402973;
   reg _402974_402974 ; 
   reg __402974_402974;
   reg _402975_402975 ; 
   reg __402975_402975;
   reg _402976_402976 ; 
   reg __402976_402976;
   reg _402977_402977 ; 
   reg __402977_402977;
   reg _402978_402978 ; 
   reg __402978_402978;
   reg _402979_402979 ; 
   reg __402979_402979;
   reg _402980_402980 ; 
   reg __402980_402980;
   reg _402981_402981 ; 
   reg __402981_402981;
   reg _402982_402982 ; 
   reg __402982_402982;
   reg _402983_402983 ; 
   reg __402983_402983;
   reg _402984_402984 ; 
   reg __402984_402984;
   reg _402985_402985 ; 
   reg __402985_402985;
   reg _402986_402986 ; 
   reg __402986_402986;
   reg _402987_402987 ; 
   reg __402987_402987;
   reg _402988_402988 ; 
   reg __402988_402988;
   reg _402989_402989 ; 
   reg __402989_402989;
   reg _402990_402990 ; 
   reg __402990_402990;
   reg _402991_402991 ; 
   reg __402991_402991;
   reg _402992_402992 ; 
   reg __402992_402992;
   reg _402993_402993 ; 
   reg __402993_402993;
   reg _402994_402994 ; 
   reg __402994_402994;
   reg _402995_402995 ; 
   reg __402995_402995;
   reg _402996_402996 ; 
   reg __402996_402996;
   reg _402997_402997 ; 
   reg __402997_402997;
   reg _402998_402998 ; 
   reg __402998_402998;
   reg _402999_402999 ; 
   reg __402999_402999;
   reg _403000_403000 ; 
   reg __403000_403000;
   reg _403001_403001 ; 
   reg __403001_403001;
   reg _403002_403002 ; 
   reg __403002_403002;
   reg _403003_403003 ; 
   reg __403003_403003;
   reg _403004_403004 ; 
   reg __403004_403004;
   reg _403005_403005 ; 
   reg __403005_403005;
   reg _403006_403006 ; 
   reg __403006_403006;
   reg _403007_403007 ; 
   reg __403007_403007;
   reg _403008_403008 ; 
   reg __403008_403008;
   reg _403009_403009 ; 
   reg __403009_403009;
   reg _403010_403010 ; 
   reg __403010_403010;
   reg _403011_403011 ; 
   reg __403011_403011;
   reg _403012_403012 ; 
   reg __403012_403012;
   reg _403013_403013 ; 
   reg __403013_403013;
   reg _403014_403014 ; 
   reg __403014_403014;
   reg _403015_403015 ; 
   reg __403015_403015;
   reg _403016_403016 ; 
   reg __403016_403016;
   reg _403017_403017 ; 
   reg __403017_403017;
   reg _403018_403018 ; 
   reg __403018_403018;
   reg _403019_403019 ; 
   reg __403019_403019;
   reg _403020_403020 ; 
   reg __403020_403020;
   reg _403021_403021 ; 
   reg __403021_403021;
   reg _403022_403022 ; 
   reg __403022_403022;
   reg _403023_403023 ; 
   reg __403023_403023;
   reg _403024_403024 ; 
   reg __403024_403024;
   reg _403025_403025 ; 
   reg __403025_403025;
   reg _403026_403026 ; 
   reg __403026_403026;
   reg _403027_403027 ; 
   reg __403027_403027;
   reg _403028_403028 ; 
   reg __403028_403028;
   reg _403029_403029 ; 
   reg __403029_403029;
   reg _403030_403030 ; 
   reg __403030_403030;
   reg _403031_403031 ; 
   reg __403031_403031;
   reg _403032_403032 ; 
   reg __403032_403032;
   reg _403033_403033 ; 
   reg __403033_403033;
   reg _403034_403034 ; 
   reg __403034_403034;
   reg _403035_403035 ; 
   reg __403035_403035;
   reg _403036_403036 ; 
   reg __403036_403036;
   reg _403037_403037 ; 
   reg __403037_403037;
   reg _403038_403038 ; 
   reg __403038_403038;
   reg _403039_403039 ; 
   reg __403039_403039;
   reg _403040_403040 ; 
   reg __403040_403040;
   reg _403041_403041 ; 
   reg __403041_403041;
   reg _403042_403042 ; 
   reg __403042_403042;
   reg _403043_403043 ; 
   reg __403043_403043;
   reg _403044_403044 ; 
   reg __403044_403044;
   reg _403045_403045 ; 
   reg __403045_403045;
   reg _403046_403046 ; 
   reg __403046_403046;
   reg _403047_403047 ; 
   reg __403047_403047;
   reg _403048_403048 ; 
   reg __403048_403048;
   reg _403049_403049 ; 
   reg __403049_403049;
   reg _403050_403050 ; 
   reg __403050_403050;
   reg _403051_403051 ; 
   reg __403051_403051;
   reg _403052_403052 ; 
   reg __403052_403052;
   reg _403053_403053 ; 
   reg __403053_403053;
   reg _403054_403054 ; 
   reg __403054_403054;
   reg _403055_403055 ; 
   reg __403055_403055;
   reg _403056_403056 ; 
   reg __403056_403056;
   reg _403057_403057 ; 
   reg __403057_403057;
   reg _403058_403058 ; 
   reg __403058_403058;
   reg _403059_403059 ; 
   reg __403059_403059;
   reg _403060_403060 ; 
   reg __403060_403060;
   reg _403061_403061 ; 
   reg __403061_403061;
   reg _403062_403062 ; 
   reg __403062_403062;
   reg _403063_403063 ; 
   reg __403063_403063;
   reg _403064_403064 ; 
   reg __403064_403064;
   reg _403065_403065 ; 
   reg __403065_403065;
   reg _403066_403066 ; 
   reg __403066_403066;
   reg _403067_403067 ; 
   reg __403067_403067;
   reg _403068_403068 ; 
   reg __403068_403068;
   reg _403069_403069 ; 
   reg __403069_403069;
   reg _403070_403070 ; 
   reg __403070_403070;
   reg _403071_403071 ; 
   reg __403071_403071;
   reg _403072_403072 ; 
   reg __403072_403072;
   reg _403073_403073 ; 
   reg __403073_403073;
   reg _403074_403074 ; 
   reg __403074_403074;
   reg _403075_403075 ; 
   reg __403075_403075;
   reg _403076_403076 ; 
   reg __403076_403076;
   reg _403077_403077 ; 
   reg __403077_403077;
   reg _403078_403078 ; 
   reg __403078_403078;
   reg _403079_403079 ; 
   reg __403079_403079;
   reg _403080_403080 ; 
   reg __403080_403080;
   reg _403081_403081 ; 
   reg __403081_403081;
   reg _403082_403082 ; 
   reg __403082_403082;
   reg _403083_403083 ; 
   reg __403083_403083;
   reg _403084_403084 ; 
   reg __403084_403084;
   reg _403085_403085 ; 
   reg __403085_403085;
   reg _403086_403086 ; 
   reg __403086_403086;
   reg _403087_403087 ; 
   reg __403087_403087;
   reg _403088_403088 ; 
   reg __403088_403088;
   reg _403089_403089 ; 
   reg __403089_403089;
   reg _403090_403090 ; 
   reg __403090_403090;
   reg _403091_403091 ; 
   reg __403091_403091;
   reg _403092_403092 ; 
   reg __403092_403092;
   reg _403093_403093 ; 
   reg __403093_403093;
   reg _403094_403094 ; 
   reg __403094_403094;
   reg _403095_403095 ; 
   reg __403095_403095;
   reg _403096_403096 ; 
   reg __403096_403096;
   reg _403097_403097 ; 
   reg __403097_403097;
   reg _403098_403098 ; 
   reg __403098_403098;
   reg _403099_403099 ; 
   reg __403099_403099;
   reg _403100_403100 ; 
   reg __403100_403100;
   reg _403101_403101 ; 
   reg __403101_403101;
   reg _403102_403102 ; 
   reg __403102_403102;
   reg _403103_403103 ; 
   reg __403103_403103;
   reg _403104_403104 ; 
   reg __403104_403104;
   reg _403105_403105 ; 
   reg __403105_403105;
   reg _403106_403106 ; 
   reg __403106_403106;
   reg _403107_403107 ; 
   reg __403107_403107;
   reg _403108_403108 ; 
   reg __403108_403108;
   reg _403109_403109 ; 
   reg __403109_403109;
   reg _403110_403110 ; 
   reg __403110_403110;
   reg _403111_403111 ; 
   reg __403111_403111;
   reg _403112_403112 ; 
   reg __403112_403112;
   reg _403113_403113 ; 
   reg __403113_403113;
   reg _403114_403114 ; 
   reg __403114_403114;
   reg _403115_403115 ; 
   reg __403115_403115;
   reg _403116_403116 ; 
   reg __403116_403116;
   reg _403117_403117 ; 
   reg __403117_403117;
   reg _403118_403118 ; 
   reg __403118_403118;
   reg _403119_403119 ; 
   reg __403119_403119;
   reg _403120_403120 ; 
   reg __403120_403120;
   reg _403121_403121 ; 
   reg __403121_403121;
   reg _403122_403122 ; 
   reg __403122_403122;
   reg _403123_403123 ; 
   reg __403123_403123;
   reg _403124_403124 ; 
   reg __403124_403124;
   reg _403125_403125 ; 
   reg __403125_403125;
   reg _403126_403126 ; 
   reg __403126_403126;
   reg _403127_403127 ; 
   reg __403127_403127;
   reg _403128_403128 ; 
   reg __403128_403128;
   reg _403129_403129 ; 
   reg __403129_403129;
   reg _403130_403130 ; 
   reg __403130_403130;
   reg _403131_403131 ; 
   reg __403131_403131;
   reg _403132_403132 ; 
   reg __403132_403132;
   reg _403133_403133 ; 
   reg __403133_403133;
   reg _403134_403134 ; 
   reg __403134_403134;
   reg _403135_403135 ; 
   reg __403135_403135;
   reg _403136_403136 ; 
   reg __403136_403136;
   reg _403137_403137 ; 
   reg __403137_403137;
   reg _403138_403138 ; 
   reg __403138_403138;
   reg _403139_403139 ; 
   reg __403139_403139;
   reg _403140_403140 ; 
   reg __403140_403140;
   reg _403141_403141 ; 
   reg __403141_403141;
   reg _403142_403142 ; 
   reg __403142_403142;
   reg _403143_403143 ; 
   reg __403143_403143;
   reg _403144_403144 ; 
   reg __403144_403144;
   reg _403145_403145 ; 
   reg __403145_403145;
   reg _403146_403146 ; 
   reg __403146_403146;
   reg _403147_403147 ; 
   reg __403147_403147;
   reg _403148_403148 ; 
   reg __403148_403148;
   reg _403149_403149 ; 
   reg __403149_403149;
   reg _403150_403150 ; 
   reg __403150_403150;
   reg _403151_403151 ; 
   reg __403151_403151;
   reg _403152_403152 ; 
   reg __403152_403152;
   reg _403153_403153 ; 
   reg __403153_403153;
   reg _403154_403154 ; 
   reg __403154_403154;
   reg _403155_403155 ; 
   reg __403155_403155;
   reg _403156_403156 ; 
   reg __403156_403156;
   reg _403157_403157 ; 
   reg __403157_403157;
   reg _403158_403158 ; 
   reg __403158_403158;
   reg _403159_403159 ; 
   reg __403159_403159;
   reg _403160_403160 ; 
   reg __403160_403160;
   reg _403161_403161 ; 
   reg __403161_403161;
   reg _403162_403162 ; 
   reg __403162_403162;
   reg _403163_403163 ; 
   reg __403163_403163;
   reg _403164_403164 ; 
   reg __403164_403164;
   reg _403165_403165 ; 
   reg __403165_403165;
   reg _403166_403166 ; 
   reg __403166_403166;
   reg _403167_403167 ; 
   reg __403167_403167;
   reg _403168_403168 ; 
   reg __403168_403168;
   reg _403169_403169 ; 
   reg __403169_403169;
   reg _403170_403170 ; 
   reg __403170_403170;
   reg _403171_403171 ; 
   reg __403171_403171;
   reg _403172_403172 ; 
   reg __403172_403172;
   reg _403173_403173 ; 
   reg __403173_403173;
   reg _403174_403174 ; 
   reg __403174_403174;
   reg _403175_403175 ; 
   reg __403175_403175;
   reg _403176_403176 ; 
   reg __403176_403176;
   reg _403177_403177 ; 
   reg __403177_403177;
   reg _403178_403178 ; 
   reg __403178_403178;
   reg _403179_403179 ; 
   reg __403179_403179;
   reg _403180_403180 ; 
   reg __403180_403180;
   reg _403181_403181 ; 
   reg __403181_403181;
   reg _403182_403182 ; 
   reg __403182_403182;
   reg _403183_403183 ; 
   reg __403183_403183;
   reg _403184_403184 ; 
   reg __403184_403184;
   reg _403185_403185 ; 
   reg __403185_403185;
   reg _403186_403186 ; 
   reg __403186_403186;
   reg _403187_403187 ; 
   reg __403187_403187;
   reg _403188_403188 ; 
   reg __403188_403188;
   reg _403189_403189 ; 
   reg __403189_403189;
   reg _403190_403190 ; 
   reg __403190_403190;
   reg _403191_403191 ; 
   reg __403191_403191;
   reg _403192_403192 ; 
   reg __403192_403192;
   reg _403193_403193 ; 
   reg __403193_403193;
   reg _403194_403194 ; 
   reg __403194_403194;
   reg _403195_403195 ; 
   reg __403195_403195;
   reg _403196_403196 ; 
   reg __403196_403196;
   reg _403197_403197 ; 
   reg __403197_403197;
   reg _403198_403198 ; 
   reg __403198_403198;
   reg _403199_403199 ; 
   reg __403199_403199;
   reg _403200_403200 ; 
   reg __403200_403200;
   reg _403201_403201 ; 
   reg __403201_403201;
   reg _403202_403202 ; 
   reg __403202_403202;
   reg _403203_403203 ; 
   reg __403203_403203;
   reg _403204_403204 ; 
   reg __403204_403204;
   reg _403205_403205 ; 
   reg __403205_403205;
   reg _403206_403206 ; 
   reg __403206_403206;
   reg _403207_403207 ; 
   reg __403207_403207;
   reg _403208_403208 ; 
   reg __403208_403208;
   reg _403209_403209 ; 
   reg __403209_403209;
   reg _403210_403210 ; 
   reg __403210_403210;
   reg _403211_403211 ; 
   reg __403211_403211;
   reg _403212_403212 ; 
   reg __403212_403212;
   reg _403213_403213 ; 
   reg __403213_403213;
   reg _403214_403214 ; 
   reg __403214_403214;
   reg _403215_403215 ; 
   reg __403215_403215;
   reg _403216_403216 ; 
   reg __403216_403216;
   reg _403217_403217 ; 
   reg __403217_403217;
   reg _403218_403218 ; 
   reg __403218_403218;
   reg _403219_403219 ; 
   reg __403219_403219;
   reg _403220_403220 ; 
   reg __403220_403220;
   reg _403221_403221 ; 
   reg __403221_403221;
   reg _403222_403222 ; 
   reg __403222_403222;
   reg _403223_403223 ; 
   reg __403223_403223;
   reg _403224_403224 ; 
   reg __403224_403224;
   reg _403225_403225 ; 
   reg __403225_403225;
   reg _403226_403226 ; 
   reg __403226_403226;
   reg _403227_403227 ; 
   reg __403227_403227;
   reg _403228_403228 ; 
   reg __403228_403228;
   reg _403229_403229 ; 
   reg __403229_403229;
   reg _403230_403230 ; 
   reg __403230_403230;
   reg _403231_403231 ; 
   reg __403231_403231;
   reg _403232_403232 ; 
   reg __403232_403232;
   reg _403233_403233 ; 
   reg __403233_403233;
   reg _403234_403234 ; 
   reg __403234_403234;
   reg _403235_403235 ; 
   reg __403235_403235;
   reg _403236_403236 ; 
   reg __403236_403236;
   reg _403237_403237 ; 
   reg __403237_403237;
   reg _403238_403238 ; 
   reg __403238_403238;
   reg _403239_403239 ; 
   reg __403239_403239;
   reg _403240_403240 ; 
   reg __403240_403240;
   reg _403241_403241 ; 
   reg __403241_403241;
   reg _403242_403242 ; 
   reg __403242_403242;
   reg _403243_403243 ; 
   reg __403243_403243;
   reg _403244_403244 ; 
   reg __403244_403244;
   reg _403245_403245 ; 
   reg __403245_403245;
   reg _403246_403246 ; 
   reg __403246_403246;
   reg _403247_403247 ; 
   reg __403247_403247;
   reg _403248_403248 ; 
   reg __403248_403248;
   reg _403249_403249 ; 
   reg __403249_403249;
   reg _403250_403250 ; 
   reg __403250_403250;
   reg _403251_403251 ; 
   reg __403251_403251;
   reg _403252_403252 ; 
   reg __403252_403252;
   reg _403253_403253 ; 
   reg __403253_403253;
   reg _403254_403254 ; 
   reg __403254_403254;
   reg _403255_403255 ; 
   reg __403255_403255;
   reg _403256_403256 ; 
   reg __403256_403256;
   reg _403257_403257 ; 
   reg __403257_403257;
   reg _403258_403258 ; 
   reg __403258_403258;
   reg _403259_403259 ; 
   reg __403259_403259;
   reg _403260_403260 ; 
   reg __403260_403260;
   reg _403261_403261 ; 
   reg __403261_403261;
   reg _403262_403262 ; 
   reg __403262_403262;
   reg _403263_403263 ; 
   reg __403263_403263;
   reg _403264_403264 ; 
   reg __403264_403264;
   reg _403265_403265 ; 
   reg __403265_403265;
   reg _403266_403266 ; 
   reg __403266_403266;
   reg _403267_403267 ; 
   reg __403267_403267;
   reg _403268_403268 ; 
   reg __403268_403268;
   reg _403269_403269 ; 
   reg __403269_403269;
   reg _403270_403270 ; 
   reg __403270_403270;
   reg _403271_403271 ; 
   reg __403271_403271;
   reg _403272_403272 ; 
   reg __403272_403272;
   reg _403273_403273 ; 
   reg __403273_403273;
   reg _403274_403274 ; 
   reg __403274_403274;
   reg _403275_403275 ; 
   reg __403275_403275;
   reg _403276_403276 ; 
   reg __403276_403276;
   reg _403277_403277 ; 
   reg __403277_403277;
   reg _403278_403278 ; 
   reg __403278_403278;
   reg _403279_403279 ; 
   reg __403279_403279;
   reg _403280_403280 ; 
   reg __403280_403280;
   reg _403281_403281 ; 
   reg __403281_403281;
   reg _403282_403282 ; 
   reg __403282_403282;
   reg _403283_403283 ; 
   reg __403283_403283;
   reg _403284_403284 ; 
   reg __403284_403284;
   reg _403285_403285 ; 
   reg __403285_403285;
   reg _403286_403286 ; 
   reg __403286_403286;
   reg _403287_403287 ; 
   reg __403287_403287;
   reg _403288_403288 ; 
   reg __403288_403288;
   reg _403289_403289 ; 
   reg __403289_403289;
   reg _403290_403290 ; 
   reg __403290_403290;
   reg _403291_403291 ; 
   reg __403291_403291;
   reg _403292_403292 ; 
   reg __403292_403292;
   reg _403293_403293 ; 
   reg __403293_403293;
   reg _403294_403294 ; 
   reg __403294_403294;
   reg _403295_403295 ; 
   reg __403295_403295;
   reg _403296_403296 ; 
   reg __403296_403296;
   reg _403297_403297 ; 
   reg __403297_403297;
   reg _403298_403298 ; 
   reg __403298_403298;
   reg _403299_403299 ; 
   reg __403299_403299;
   reg _403300_403300 ; 
   reg __403300_403300;
   reg _403301_403301 ; 
   reg __403301_403301;
   reg _403302_403302 ; 
   reg __403302_403302;
   reg _403303_403303 ; 
   reg __403303_403303;
   reg _403304_403304 ; 
   reg __403304_403304;
   reg _403305_403305 ; 
   reg __403305_403305;
   reg _403306_403306 ; 
   reg __403306_403306;
   reg _403307_403307 ; 
   reg __403307_403307;
   reg _403308_403308 ; 
   reg __403308_403308;
   reg _403309_403309 ; 
   reg __403309_403309;
   reg _403310_403310 ; 
   reg __403310_403310;
   reg _403311_403311 ; 
   reg __403311_403311;
   reg _403312_403312 ; 
   reg __403312_403312;
   reg _403313_403313 ; 
   reg __403313_403313;
   reg _403314_403314 ; 
   reg __403314_403314;
   reg _403315_403315 ; 
   reg __403315_403315;
   reg _403316_403316 ; 
   reg __403316_403316;
   reg _403317_403317 ; 
   reg __403317_403317;
   reg _403318_403318 ; 
   reg __403318_403318;
   reg _403319_403319 ; 
   reg __403319_403319;
   reg _403320_403320 ; 
   reg __403320_403320;
   reg _403321_403321 ; 
   reg __403321_403321;
   reg _403322_403322 ; 
   reg __403322_403322;
   reg _403323_403323 ; 
   reg __403323_403323;
   reg _403324_403324 ; 
   reg __403324_403324;
   reg _403325_403325 ; 
   reg __403325_403325;
   reg _403326_403326 ; 
   reg __403326_403326;
   reg _403327_403327 ; 
   reg __403327_403327;
   reg _403328_403328 ; 
   reg __403328_403328;
   reg _403329_403329 ; 
   reg __403329_403329;
   reg _403330_403330 ; 
   reg __403330_403330;
   reg _403331_403331 ; 
   reg __403331_403331;
   reg _403332_403332 ; 
   reg __403332_403332;
   reg _403333_403333 ; 
   reg __403333_403333;
   reg _403334_403334 ; 
   reg __403334_403334;
   reg _403335_403335 ; 
   reg __403335_403335;
   reg _403336_403336 ; 
   reg __403336_403336;
   reg _403337_403337 ; 
   reg __403337_403337;
   reg _403338_403338 ; 
   reg __403338_403338;
   reg _403339_403339 ; 
   reg __403339_403339;
   reg _403340_403340 ; 
   reg __403340_403340;
   reg _403341_403341 ; 
   reg __403341_403341;
   reg _403342_403342 ; 
   reg __403342_403342;
   reg _403343_403343 ; 
   reg __403343_403343;
   reg _403344_403344 ; 
   reg __403344_403344;
   reg _403345_403345 ; 
   reg __403345_403345;
   reg _403346_403346 ; 
   reg __403346_403346;
   reg _403347_403347 ; 
   reg __403347_403347;
   reg _403348_403348 ; 
   reg __403348_403348;
   reg _403349_403349 ; 
   reg __403349_403349;
   reg _403350_403350 ; 
   reg __403350_403350;
   reg _403351_403351 ; 
   reg __403351_403351;
   reg _403352_403352 ; 
   reg __403352_403352;
   reg _403353_403353 ; 
   reg __403353_403353;
   reg _403354_403354 ; 
   reg __403354_403354;
   reg _403355_403355 ; 
   reg __403355_403355;
   reg _403356_403356 ; 
   reg __403356_403356;
   reg _403357_403357 ; 
   reg __403357_403357;
   reg _403358_403358 ; 
   reg __403358_403358;
   reg _403359_403359 ; 
   reg __403359_403359;
   reg _403360_403360 ; 
   reg __403360_403360;
   reg _403361_403361 ; 
   reg __403361_403361;
   reg _403362_403362 ; 
   reg __403362_403362;
   reg _403363_403363 ; 
   reg __403363_403363;
   reg _403364_403364 ; 
   reg __403364_403364;
   reg _403365_403365 ; 
   reg __403365_403365;
   reg _403366_403366 ; 
   reg __403366_403366;
   reg _403367_403367 ; 
   reg __403367_403367;
   reg _403368_403368 ; 
   reg __403368_403368;
   reg _403369_403369 ; 
   reg __403369_403369;
   reg _403370_403370 ; 
   reg __403370_403370;
   reg _403371_403371 ; 
   reg __403371_403371;
   reg _403372_403372 ; 
   reg __403372_403372;
   reg _403373_403373 ; 
   reg __403373_403373;
   reg _403374_403374 ; 
   reg __403374_403374;
   reg _403375_403375 ; 
   reg __403375_403375;
   reg _403376_403376 ; 
   reg __403376_403376;
   reg _403377_403377 ; 
   reg __403377_403377;
   reg _403378_403378 ; 
   reg __403378_403378;
   reg _403379_403379 ; 
   reg __403379_403379;
   reg _403380_403380 ; 
   reg __403380_403380;
   reg _403381_403381 ; 
   reg __403381_403381;
   reg _403382_403382 ; 
   reg __403382_403382;
   reg _403383_403383 ; 
   reg __403383_403383;
   reg _403384_403384 ; 
   reg __403384_403384;
   reg _403385_403385 ; 
   reg __403385_403385;
   reg _403386_403386 ; 
   reg __403386_403386;
   reg _403387_403387 ; 
   reg __403387_403387;
   reg _403388_403388 ; 
   reg __403388_403388;
   reg _403389_403389 ; 
   reg __403389_403389;
   reg _403390_403390 ; 
   reg __403390_403390;
   reg _403391_403391 ; 
   reg __403391_403391;
   reg _403392_403392 ; 
   reg __403392_403392;
   reg _403393_403393 ; 
   reg __403393_403393;
   reg _403394_403394 ; 
   reg __403394_403394;
   reg _403395_403395 ; 
   reg __403395_403395;
   reg _403396_403396 ; 
   reg __403396_403396;
   reg _403397_403397 ; 
   reg __403397_403397;
   reg _403398_403398 ; 
   reg __403398_403398;
   reg _403399_403399 ; 
   reg __403399_403399;
   reg _403400_403400 ; 
   reg __403400_403400;
   reg _403401_403401 ; 
   reg __403401_403401;
   reg _403402_403402 ; 
   reg __403402_403402;
   reg _403403_403403 ; 
   reg __403403_403403;
   reg _403404_403404 ; 
   reg __403404_403404;
   reg _403405_403405 ; 
   reg __403405_403405;
   reg _403406_403406 ; 
   reg __403406_403406;
   reg _403407_403407 ; 
   reg __403407_403407;
   reg _403408_403408 ; 
   reg __403408_403408;
   reg _403409_403409 ; 
   reg __403409_403409;
   reg _403410_403410 ; 
   reg __403410_403410;
   reg _403411_403411 ; 
   reg __403411_403411;
   reg _403412_403412 ; 
   reg __403412_403412;
   reg _403413_403413 ; 
   reg __403413_403413;
   reg _403414_403414 ; 
   reg __403414_403414;
   reg _403415_403415 ; 
   reg __403415_403415;
   reg _403416_403416 ; 
   reg __403416_403416;
   reg _403417_403417 ; 
   reg __403417_403417;
   reg _403418_403418 ; 
   reg __403418_403418;
   reg _403419_403419 ; 
   reg __403419_403419;
   reg _403420_403420 ; 
   reg __403420_403420;
   reg _403421_403421 ; 
   reg __403421_403421;
   reg _403422_403422 ; 
   reg __403422_403422;
   reg _403423_403423 ; 
   reg __403423_403423;
   reg _403424_403424 ; 
   reg __403424_403424;
   reg _403425_403425 ; 
   reg __403425_403425;
   reg _403426_403426 ; 
   reg __403426_403426;
   reg _403427_403427 ; 
   reg __403427_403427;
   reg _403428_403428 ; 
   reg __403428_403428;
   reg _403429_403429 ; 
   reg __403429_403429;
   reg _403430_403430 ; 
   reg __403430_403430;
   reg _403431_403431 ; 
   reg __403431_403431;
   reg _403432_403432 ; 
   reg __403432_403432;
   reg _403433_403433 ; 
   reg __403433_403433;
   reg _403434_403434 ; 
   reg __403434_403434;
   reg _403435_403435 ; 
   reg __403435_403435;
   reg _403436_403436 ; 
   reg __403436_403436;
   reg _403437_403437 ; 
   reg __403437_403437;
   reg _403438_403438 ; 
   reg __403438_403438;
   reg _403439_403439 ; 
   reg __403439_403439;
   reg _403440_403440 ; 
   reg __403440_403440;
   reg _403441_403441 ; 
   reg __403441_403441;
   reg _403442_403442 ; 
   reg __403442_403442;
   reg _403443_403443 ; 
   reg __403443_403443;
   reg _403444_403444 ; 
   reg __403444_403444;
   reg _403445_403445 ; 
   reg __403445_403445;
   reg _403446_403446 ; 
   reg __403446_403446;
   reg _403447_403447 ; 
   reg __403447_403447;
   reg _403448_403448 ; 
   reg __403448_403448;
   reg _403449_403449 ; 
   reg __403449_403449;
   reg _403450_403450 ; 
   reg __403450_403450;
   reg _403451_403451 ; 
   reg __403451_403451;
   reg _403452_403452 ; 
   reg __403452_403452;
   reg _403453_403453 ; 
   reg __403453_403453;
   reg _403454_403454 ; 
   reg __403454_403454;
   reg _403455_403455 ; 
   reg __403455_403455;
   reg _403456_403456 ; 
   reg __403456_403456;
   reg _403457_403457 ; 
   reg __403457_403457;
   reg _403458_403458 ; 
   reg __403458_403458;
   reg _403459_403459 ; 
   reg __403459_403459;
   reg _403460_403460 ; 
   reg __403460_403460;
   reg _403461_403461 ; 
   reg __403461_403461;
   reg _403462_403462 ; 
   reg __403462_403462;
   reg _403463_403463 ; 
   reg __403463_403463;
   reg _403464_403464 ; 
   reg __403464_403464;
   reg _403465_403465 ; 
   reg __403465_403465;
   reg _403466_403466 ; 
   reg __403466_403466;
   reg _403467_403467 ; 
   reg __403467_403467;
   reg _403468_403468 ; 
   reg __403468_403468;
   reg _403469_403469 ; 
   reg __403469_403469;
   reg _403470_403470 ; 
   reg __403470_403470;
   reg _403471_403471 ; 
   reg __403471_403471;
   reg _403472_403472 ; 
   reg __403472_403472;
   reg _403473_403473 ; 
   reg __403473_403473;
   reg _403474_403474 ; 
   reg __403474_403474;
   reg _403475_403475 ; 
   reg __403475_403475;
   reg _403476_403476 ; 
   reg __403476_403476;
   reg _403477_403477 ; 
   reg __403477_403477;
   reg _403478_403478 ; 
   reg __403478_403478;
   reg _403479_403479 ; 
   reg __403479_403479;
   reg _403480_403480 ; 
   reg __403480_403480;
   reg _403481_403481 ; 
   reg __403481_403481;
   reg _403482_403482 ; 
   reg __403482_403482;
   reg _403483_403483 ; 
   reg __403483_403483;
   reg _403484_403484 ; 
   reg __403484_403484;
   reg _403485_403485 ; 
   reg __403485_403485;
   reg _403486_403486 ; 
   reg __403486_403486;
   reg _403487_403487 ; 
   reg __403487_403487;
   reg _403488_403488 ; 
   reg __403488_403488;
   reg _403489_403489 ; 
   reg __403489_403489;
   reg _403490_403490 ; 
   reg __403490_403490;
   reg _403491_403491 ; 
   reg __403491_403491;
   reg _403492_403492 ; 
   reg __403492_403492;
   reg _403493_403493 ; 
   reg __403493_403493;
   reg _403494_403494 ; 
   reg __403494_403494;
   reg _403495_403495 ; 
   reg __403495_403495;
   reg _403496_403496 ; 
   reg __403496_403496;
   reg _403497_403497 ; 
   reg __403497_403497;
   reg _403498_403498 ; 
   reg __403498_403498;
   reg _403499_403499 ; 
   reg __403499_403499;
   reg _403500_403500 ; 
   reg __403500_403500;
   reg _403501_403501 ; 
   reg __403501_403501;
   reg _403502_403502 ; 
   reg __403502_403502;
   reg _403503_403503 ; 
   reg __403503_403503;
   reg _403504_403504 ; 
   reg __403504_403504;
   reg _403505_403505 ; 
   reg __403505_403505;
   reg _403506_403506 ; 
   reg __403506_403506;
   reg _403507_403507 ; 
   reg __403507_403507;
   reg _403508_403508 ; 
   reg __403508_403508;
   reg _403509_403509 ; 
   reg __403509_403509;
   reg _403510_403510 ; 
   reg __403510_403510;
   reg _403511_403511 ; 
   reg __403511_403511;
   reg _403512_403512 ; 
   reg __403512_403512;
   reg _403513_403513 ; 
   reg __403513_403513;
   reg _403514_403514 ; 
   reg __403514_403514;
   reg _403515_403515 ; 
   reg __403515_403515;
   reg _403516_403516 ; 
   reg __403516_403516;
   reg _403517_403517 ; 
   reg __403517_403517;
   reg _403518_403518 ; 
   reg __403518_403518;
   reg _403519_403519 ; 
   reg __403519_403519;
   reg _403520_403520 ; 
   reg __403520_403520;
   reg _403521_403521 ; 
   reg __403521_403521;
   reg _403522_403522 ; 
   reg __403522_403522;
   reg _403523_403523 ; 
   reg __403523_403523;
   reg _403524_403524 ; 
   reg __403524_403524;
   reg _403525_403525 ; 
   reg __403525_403525;
   reg _403526_403526 ; 
   reg __403526_403526;
   reg _403527_403527 ; 
   reg __403527_403527;
   reg _403528_403528 ; 
   reg __403528_403528;
   reg _403529_403529 ; 
   reg __403529_403529;
   reg _403530_403530 ; 
   reg __403530_403530;
   reg _403531_403531 ; 
   reg __403531_403531;
   reg _403532_403532 ; 
   reg __403532_403532;
   reg _403533_403533 ; 
   reg __403533_403533;
   reg _403534_403534 ; 
   reg __403534_403534;
   reg _403535_403535 ; 
   reg __403535_403535;
   reg _403536_403536 ; 
   reg __403536_403536;
   reg _403537_403537 ; 
   reg __403537_403537;
   reg _403538_403538 ; 
   reg __403538_403538;
   reg _403539_403539 ; 
   reg __403539_403539;
   reg _403540_403540 ; 
   reg __403540_403540;
   reg _403541_403541 ; 
   reg __403541_403541;
   reg _403542_403542 ; 
   reg __403542_403542;
   reg _403543_403543 ; 
   reg __403543_403543;
   reg _403544_403544 ; 
   reg __403544_403544;
   reg _403545_403545 ; 
   reg __403545_403545;
   reg _403546_403546 ; 
   reg __403546_403546;
   reg _403547_403547 ; 
   reg __403547_403547;
   reg _403548_403548 ; 
   reg __403548_403548;
   reg _403549_403549 ; 
   reg __403549_403549;
   reg _403550_403550 ; 
   reg __403550_403550;
   reg _403551_403551 ; 
   reg __403551_403551;
   reg _403552_403552 ; 
   reg __403552_403552;
   reg _403553_403553 ; 
   reg __403553_403553;
   reg _403554_403554 ; 
   reg __403554_403554;
   reg _403555_403555 ; 
   reg __403555_403555;
   reg _403556_403556 ; 
   reg __403556_403556;
   reg _403557_403557 ; 
   reg __403557_403557;
   reg _403558_403558 ; 
   reg __403558_403558;
   reg _403559_403559 ; 
   reg __403559_403559;
   reg _403560_403560 ; 
   reg __403560_403560;
   reg _403561_403561 ; 
   reg __403561_403561;
   reg _403562_403562 ; 
   reg __403562_403562;
   reg _403563_403563 ; 
   reg __403563_403563;
   reg _403564_403564 ; 
   reg __403564_403564;
   reg _403565_403565 ; 
   reg __403565_403565;
   reg _403566_403566 ; 
   reg __403566_403566;
   reg _403567_403567 ; 
   reg __403567_403567;
   reg _403568_403568 ; 
   reg __403568_403568;
   reg _403569_403569 ; 
   reg __403569_403569;
   reg _403570_403570 ; 
   reg __403570_403570;
   reg _403571_403571 ; 
   reg __403571_403571;
   reg _403572_403572 ; 
   reg __403572_403572;
   reg _403573_403573 ; 
   reg __403573_403573;
   reg _403574_403574 ; 
   reg __403574_403574;
   reg _403575_403575 ; 
   reg __403575_403575;
   reg _403576_403576 ; 
   reg __403576_403576;
   reg _403577_403577 ; 
   reg __403577_403577;
   reg _403578_403578 ; 
   reg __403578_403578;
   reg _403579_403579 ; 
   reg __403579_403579;
   reg _403580_403580 ; 
   reg __403580_403580;
   reg _403581_403581 ; 
   reg __403581_403581;
   reg _403582_403582 ; 
   reg __403582_403582;
   reg _403583_403583 ; 
   reg __403583_403583;
   reg _403584_403584 ; 
   reg __403584_403584;
   reg _403585_403585 ; 
   reg __403585_403585;
   reg _403586_403586 ; 
   reg __403586_403586;
   reg _403587_403587 ; 
   reg __403587_403587;
   reg _403588_403588 ; 
   reg __403588_403588;
   reg _403589_403589 ; 
   reg __403589_403589;
   reg _403590_403590 ; 
   reg __403590_403590;
   reg _403591_403591 ; 
   reg __403591_403591;
   reg _403592_403592 ; 
   reg __403592_403592;
   reg _403593_403593 ; 
   reg __403593_403593;
   reg _403594_403594 ; 
   reg __403594_403594;
   reg _403595_403595 ; 
   reg __403595_403595;
   reg _403596_403596 ; 
   reg __403596_403596;
   reg _403597_403597 ; 
   reg __403597_403597;
   reg _403598_403598 ; 
   reg __403598_403598;
   reg _403599_403599 ; 
   reg __403599_403599;
   reg _403600_403600 ; 
   reg __403600_403600;
   reg _403601_403601 ; 
   reg __403601_403601;
   reg _403602_403602 ; 
   reg __403602_403602;
   reg _403603_403603 ; 
   reg __403603_403603;
   reg _403604_403604 ; 
   reg __403604_403604;
   reg _403605_403605 ; 
   reg __403605_403605;
   reg _403606_403606 ; 
   reg __403606_403606;
   reg _403607_403607 ; 
   reg __403607_403607;
   reg _403608_403608 ; 
   reg __403608_403608;
   reg _403609_403609 ; 
   reg __403609_403609;
   reg _403610_403610 ; 
   reg __403610_403610;
   reg _403611_403611 ; 
   reg __403611_403611;
   reg _403612_403612 ; 
   reg __403612_403612;
   reg _403613_403613 ; 
   reg __403613_403613;
   reg _403614_403614 ; 
   reg __403614_403614;
   reg _403615_403615 ; 
   reg __403615_403615;
   reg _403616_403616 ; 
   reg __403616_403616;
   reg _403617_403617 ; 
   reg __403617_403617;
   reg _403618_403618 ; 
   reg __403618_403618;
   reg _403619_403619 ; 
   reg __403619_403619;
   reg _403620_403620 ; 
   reg __403620_403620;
   reg _403621_403621 ; 
   reg __403621_403621;
   reg _403622_403622 ; 
   reg __403622_403622;
   reg _403623_403623 ; 
   reg __403623_403623;
   reg _403624_403624 ; 
   reg __403624_403624;
   reg _403625_403625 ; 
   reg __403625_403625;
   reg _403626_403626 ; 
   reg __403626_403626;
   reg _403627_403627 ; 
   reg __403627_403627;
   reg _403628_403628 ; 
   reg __403628_403628;
   reg _403629_403629 ; 
   reg __403629_403629;
   reg _403630_403630 ; 
   reg __403630_403630;
   reg _403631_403631 ; 
   reg __403631_403631;
   reg _403632_403632 ; 
   reg __403632_403632;
   reg _403633_403633 ; 
   reg __403633_403633;
   reg _403634_403634 ; 
   reg __403634_403634;
   reg _403635_403635 ; 
   reg __403635_403635;
   reg _403636_403636 ; 
   reg __403636_403636;
   reg _403637_403637 ; 
   reg __403637_403637;
   reg _403638_403638 ; 
   reg __403638_403638;
   reg _403639_403639 ; 
   reg __403639_403639;
   reg _403640_403640 ; 
   reg __403640_403640;
   reg _403641_403641 ; 
   reg __403641_403641;
   reg _403642_403642 ; 
   reg __403642_403642;
   reg _403643_403643 ; 
   reg __403643_403643;
   reg _403644_403644 ; 
   reg __403644_403644;
   reg _403645_403645 ; 
   reg __403645_403645;
   reg _403646_403646 ; 
   reg __403646_403646;
   reg _403647_403647 ; 
   reg __403647_403647;
   reg _403648_403648 ; 
   reg __403648_403648;
   reg _403649_403649 ; 
   reg __403649_403649;
   reg _403650_403650 ; 
   reg __403650_403650;
   reg _403651_403651 ; 
   reg __403651_403651;
   reg _403652_403652 ; 
   reg __403652_403652;
   reg _403653_403653 ; 
   reg __403653_403653;
   reg _403654_403654 ; 
   reg __403654_403654;
   reg _403655_403655 ; 
   reg __403655_403655;
   reg _403656_403656 ; 
   reg __403656_403656;
   reg _403657_403657 ; 
   reg __403657_403657;
   reg _403658_403658 ; 
   reg __403658_403658;
   reg _403659_403659 ; 
   reg __403659_403659;
   reg _403660_403660 ; 
   reg __403660_403660;
   reg _403661_403661 ; 
   reg __403661_403661;
   reg _403662_403662 ; 
   reg __403662_403662;
   reg _403663_403663 ; 
   reg __403663_403663;
   reg _403664_403664 ; 
   reg __403664_403664;
   reg _403665_403665 ; 
   reg __403665_403665;
   reg _403666_403666 ; 
   reg __403666_403666;
   reg _403667_403667 ; 
   reg __403667_403667;
   reg _403668_403668 ; 
   reg __403668_403668;
   reg _403669_403669 ; 
   reg __403669_403669;
   reg _403670_403670 ; 
   reg __403670_403670;
   reg _403671_403671 ; 
   reg __403671_403671;
   reg _403672_403672 ; 
   reg __403672_403672;
   reg _403673_403673 ; 
   reg __403673_403673;
   reg _403674_403674 ; 
   reg __403674_403674;
   reg _403675_403675 ; 
   reg __403675_403675;
   reg _403676_403676 ; 
   reg __403676_403676;
   reg _403677_403677 ; 
   reg __403677_403677;
   reg _403678_403678 ; 
   reg __403678_403678;
   reg _403679_403679 ; 
   reg __403679_403679;
   reg _403680_403680 ; 
   reg __403680_403680;
   reg _403681_403681 ; 
   reg __403681_403681;
   reg _403682_403682 ; 
   reg __403682_403682;
   reg _403683_403683 ; 
   reg __403683_403683;
   reg _403684_403684 ; 
   reg __403684_403684;
   reg _403685_403685 ; 
   reg __403685_403685;
   reg _403686_403686 ; 
   reg __403686_403686;
   reg _403687_403687 ; 
   reg __403687_403687;
   reg _403688_403688 ; 
   reg __403688_403688;
   reg _403689_403689 ; 
   reg __403689_403689;
   reg _403690_403690 ; 
   reg __403690_403690;
   reg _403691_403691 ; 
   reg __403691_403691;
   reg _403692_403692 ; 
   reg __403692_403692;
   reg _403693_403693 ; 
   reg __403693_403693;
   reg _403694_403694 ; 
   reg __403694_403694;
   reg _403695_403695 ; 
   reg __403695_403695;
   reg _403696_403696 ; 
   reg __403696_403696;
   reg _403697_403697 ; 
   reg __403697_403697;
   reg _403698_403698 ; 
   reg __403698_403698;
   reg _403699_403699 ; 
   reg __403699_403699;
   reg _403700_403700 ; 
   reg __403700_403700;
   reg _403701_403701 ; 
   reg __403701_403701;
   reg _403702_403702 ; 
   reg __403702_403702;
   reg _403703_403703 ; 
   reg __403703_403703;
   reg _403704_403704 ; 
   reg __403704_403704;
   reg _403705_403705 ; 
   reg __403705_403705;
   reg _403706_403706 ; 
   reg __403706_403706;
   reg _403707_403707 ; 
   reg __403707_403707;
   reg _403708_403708 ; 
   reg __403708_403708;
   reg _403709_403709 ; 
   reg __403709_403709;
   reg _403710_403710 ; 
   reg __403710_403710;
   reg _403711_403711 ; 
   reg __403711_403711;
   reg _403712_403712 ; 
   reg __403712_403712;
   reg _403713_403713 ; 
   reg __403713_403713;
   reg _403714_403714 ; 
   reg __403714_403714;
   reg _403715_403715 ; 
   reg __403715_403715;
   reg _403716_403716 ; 
   reg __403716_403716;
   reg _403717_403717 ; 
   reg __403717_403717;
   reg _403718_403718 ; 
   reg __403718_403718;
   reg _403719_403719 ; 
   reg __403719_403719;
   reg _403720_403720 ; 
   reg __403720_403720;
   reg _403721_403721 ; 
   reg __403721_403721;
   reg _403722_403722 ; 
   reg __403722_403722;
   reg _403723_403723 ; 
   reg __403723_403723;
   reg _403724_403724 ; 
   reg __403724_403724;
   reg _403725_403725 ; 
   reg __403725_403725;
   reg _403726_403726 ; 
   reg __403726_403726;
   reg _403727_403727 ; 
   reg __403727_403727;
   reg _403728_403728 ; 
   reg __403728_403728;
   reg _403729_403729 ; 
   reg __403729_403729;
   reg _403730_403730 ; 
   reg __403730_403730;
   reg _403731_403731 ; 
   reg __403731_403731;
   reg _403732_403732 ; 
   reg __403732_403732;
   reg _403733_403733 ; 
   reg __403733_403733;
   reg _403734_403734 ; 
   reg __403734_403734;
   reg _403735_403735 ; 
   reg __403735_403735;
   reg _403736_403736 ; 
   reg __403736_403736;
   reg _403737_403737 ; 
   reg __403737_403737;
   reg _403738_403738 ; 
   reg __403738_403738;
   reg _403739_403739 ; 
   reg __403739_403739;
   reg _403740_403740 ; 
   reg __403740_403740;
   reg _403741_403741 ; 
   reg __403741_403741;
   reg _403742_403742 ; 
   reg __403742_403742;
   reg _403743_403743 ; 
   reg __403743_403743;
   reg _403744_403744 ; 
   reg __403744_403744;
   reg _403745_403745 ; 
   reg __403745_403745;
   reg _403746_403746 ; 
   reg __403746_403746;
   reg _403747_403747 ; 
   reg __403747_403747;
   reg _403748_403748 ; 
   reg __403748_403748;
   reg _403749_403749 ; 
   reg __403749_403749;
   reg _403750_403750 ; 
   reg __403750_403750;
   reg _403751_403751 ; 
   reg __403751_403751;
   reg _403752_403752 ; 
   reg __403752_403752;
   reg _403753_403753 ; 
   reg __403753_403753;
   reg _403754_403754 ; 
   reg __403754_403754;
   reg _403755_403755 ; 
   reg __403755_403755;
   reg _403756_403756 ; 
   reg __403756_403756;
   reg _403757_403757 ; 
   reg __403757_403757;
   reg _403758_403758 ; 
   reg __403758_403758;
   reg _403759_403759 ; 
   reg __403759_403759;
   reg _403760_403760 ; 
   reg __403760_403760;
   reg _403761_403761 ; 
   reg __403761_403761;
   reg _403762_403762 ; 
   reg __403762_403762;
   reg _403763_403763 ; 
   reg __403763_403763;
   reg _403764_403764 ; 
   reg __403764_403764;
   reg _403765_403765 ; 
   reg __403765_403765;
   reg _403766_403766 ; 
   reg __403766_403766;
   reg _403767_403767 ; 
   reg __403767_403767;
   reg _403768_403768 ; 
   reg __403768_403768;
   reg _403769_403769 ; 
   reg __403769_403769;
   reg _403770_403770 ; 
   reg __403770_403770;
   reg _403771_403771 ; 
   reg __403771_403771;
   reg _403772_403772 ; 
   reg __403772_403772;
   reg _403773_403773 ; 
   reg __403773_403773;
   reg _403774_403774 ; 
   reg __403774_403774;
   reg _403775_403775 ; 
   reg __403775_403775;
   reg _403776_403776 ; 
   reg __403776_403776;
   reg _403777_403777 ; 
   reg __403777_403777;
   reg _403778_403778 ; 
   reg __403778_403778;
   reg _403779_403779 ; 
   reg __403779_403779;
   reg _403780_403780 ; 
   reg __403780_403780;
   reg _403781_403781 ; 
   reg __403781_403781;
   reg _403782_403782 ; 
   reg __403782_403782;
   reg _403783_403783 ; 
   reg __403783_403783;
   reg _403784_403784 ; 
   reg __403784_403784;
   reg _403785_403785 ; 
   reg __403785_403785;
   reg _403786_403786 ; 
   reg __403786_403786;
   reg _403787_403787 ; 
   reg __403787_403787;
   reg _403788_403788 ; 
   reg __403788_403788;
   reg _403789_403789 ; 
   reg __403789_403789;
   reg _403790_403790 ; 
   reg __403790_403790;
   reg _403791_403791 ; 
   reg __403791_403791;
   reg _403792_403792 ; 
   reg __403792_403792;
   reg _403793_403793 ; 
   reg __403793_403793;
   reg _403794_403794 ; 
   reg __403794_403794;
   reg _403795_403795 ; 
   reg __403795_403795;
   reg _403796_403796 ; 
   reg __403796_403796;
   reg _403797_403797 ; 
   reg __403797_403797;
   reg _403798_403798 ; 
   reg __403798_403798;
   reg _403799_403799 ; 
   reg __403799_403799;
   reg _403800_403800 ; 
   reg __403800_403800;
   reg _403801_403801 ; 
   reg __403801_403801;
   reg _403802_403802 ; 
   reg __403802_403802;
   reg _403803_403803 ; 
   reg __403803_403803;
   reg _403804_403804 ; 
   reg __403804_403804;
   reg _403805_403805 ; 
   reg __403805_403805;
   reg _403806_403806 ; 
   reg __403806_403806;
   reg _403807_403807 ; 
   reg __403807_403807;
   reg _403808_403808 ; 
   reg __403808_403808;
   reg _403809_403809 ; 
   reg __403809_403809;
   reg _403810_403810 ; 
   reg __403810_403810;
   reg _403811_403811 ; 
   reg __403811_403811;
   reg _403812_403812 ; 
   reg __403812_403812;
   reg _403813_403813 ; 
   reg __403813_403813;
   reg _403814_403814 ; 
   reg __403814_403814;
   reg _403815_403815 ; 
   reg __403815_403815;
   reg _403816_403816 ; 
   reg __403816_403816;
   reg _403817_403817 ; 
   reg __403817_403817;
   reg _403818_403818 ; 
   reg __403818_403818;
   reg _403819_403819 ; 
   reg __403819_403819;
   reg _403820_403820 ; 
   reg __403820_403820;
   reg _403821_403821 ; 
   reg __403821_403821;
   reg _403822_403822 ; 
   reg __403822_403822;
   reg _403823_403823 ; 
   reg __403823_403823;
   reg _403824_403824 ; 
   reg __403824_403824;
   reg _403825_403825 ; 
   reg __403825_403825;
   reg _403826_403826 ; 
   reg __403826_403826;
   reg _403827_403827 ; 
   reg __403827_403827;
   reg _403828_403828 ; 
   reg __403828_403828;
   reg _403829_403829 ; 
   reg __403829_403829;
   reg _403830_403830 ; 
   reg __403830_403830;
   reg _403831_403831 ; 
   reg __403831_403831;
   reg _403832_403832 ; 
   reg __403832_403832;
   reg _403833_403833 ; 
   reg __403833_403833;
   reg _403834_403834 ; 
   reg __403834_403834;
   reg _403835_403835 ; 
   reg __403835_403835;
   reg _403836_403836 ; 
   reg __403836_403836;
   reg _403837_403837 ; 
   reg __403837_403837;
   reg _403838_403838 ; 
   reg __403838_403838;
   reg _403839_403839 ; 
   reg __403839_403839;
   reg _403840_403840 ; 
   reg __403840_403840;
   reg _403841_403841 ; 
   reg __403841_403841;
   reg _403842_403842 ; 
   reg __403842_403842;
   reg _403843_403843 ; 
   reg __403843_403843;
   reg _403844_403844 ; 
   reg __403844_403844;
   reg _403845_403845 ; 
   reg __403845_403845;
   reg _403846_403846 ; 
   reg __403846_403846;
   reg _403847_403847 ; 
   reg __403847_403847;
   reg _403848_403848 ; 
   reg __403848_403848;
   reg _403849_403849 ; 
   reg __403849_403849;
   reg _403850_403850 ; 
   reg __403850_403850;
   reg _403851_403851 ; 
   reg __403851_403851;
   reg _403852_403852 ; 
   reg __403852_403852;
   reg _403853_403853 ; 
   reg __403853_403853;
   reg _403854_403854 ; 
   reg __403854_403854;
   reg _403855_403855 ; 
   reg __403855_403855;
   reg _403856_403856 ; 
   reg __403856_403856;
   reg _403857_403857 ; 
   reg __403857_403857;
   reg _403858_403858 ; 
   reg __403858_403858;
   reg _403859_403859 ; 
   reg __403859_403859;
   reg _403860_403860 ; 
   reg __403860_403860;
   reg _403861_403861 ; 
   reg __403861_403861;
   reg _403862_403862 ; 
   reg __403862_403862;
   reg _403863_403863 ; 
   reg __403863_403863;
   reg _403864_403864 ; 
   reg __403864_403864;
   reg _403865_403865 ; 
   reg __403865_403865;
   reg _403866_403866 ; 
   reg __403866_403866;
   reg _403867_403867 ; 
   reg __403867_403867;
   reg _403868_403868 ; 
   reg __403868_403868;
   reg _403869_403869 ; 
   reg __403869_403869;
   reg _403870_403870 ; 
   reg __403870_403870;
   reg _403871_403871 ; 
   reg __403871_403871;
   reg _403872_403872 ; 
   reg __403872_403872;
   reg _403873_403873 ; 
   reg __403873_403873;
   reg _403874_403874 ; 
   reg __403874_403874;
   reg _403875_403875 ; 
   reg __403875_403875;
   reg _403876_403876 ; 
   reg __403876_403876;
   reg _403877_403877 ; 
   reg __403877_403877;
   reg _403878_403878 ; 
   reg __403878_403878;
   reg _403879_403879 ; 
   reg __403879_403879;
   reg _403880_403880 ; 
   reg __403880_403880;
   reg _403881_403881 ; 
   reg __403881_403881;
   reg _403882_403882 ; 
   reg __403882_403882;
   reg _403883_403883 ; 
   reg __403883_403883;
   reg _403884_403884 ; 
   reg __403884_403884;
   reg _403885_403885 ; 
   reg __403885_403885;
   reg _403886_403886 ; 
   reg __403886_403886;
   reg _403887_403887 ; 
   reg __403887_403887;
   reg _403888_403888 ; 
   reg __403888_403888;
   reg _403889_403889 ; 
   reg __403889_403889;
   reg _403890_403890 ; 
   reg __403890_403890;
   reg _403891_403891 ; 
   reg __403891_403891;
   reg _403892_403892 ; 
   reg __403892_403892;
   reg _403893_403893 ; 
   reg __403893_403893;
   reg _403894_403894 ; 
   reg __403894_403894;
   reg _403895_403895 ; 
   reg __403895_403895;
   reg _403896_403896 ; 
   reg __403896_403896;
   reg _403897_403897 ; 
   reg __403897_403897;
   reg _403898_403898 ; 
   reg __403898_403898;
   reg _403899_403899 ; 
   reg __403899_403899;
   reg _403900_403900 ; 
   reg __403900_403900;
   reg _403901_403901 ; 
   reg __403901_403901;
   reg _403902_403902 ; 
   reg __403902_403902;
   reg _403903_403903 ; 
   reg __403903_403903;
   reg _403904_403904 ; 
   reg __403904_403904;
   reg _403905_403905 ; 
   reg __403905_403905;
   reg _403906_403906 ; 
   reg __403906_403906;
   reg _403907_403907 ; 
   reg __403907_403907;
   reg _403908_403908 ; 
   reg __403908_403908;
   reg _403909_403909 ; 
   reg __403909_403909;
   reg _403910_403910 ; 
   reg __403910_403910;
   reg _403911_403911 ; 
   reg __403911_403911;
   reg _403912_403912 ; 
   reg __403912_403912;
   reg _403913_403913 ; 
   reg __403913_403913;
   reg _403914_403914 ; 
   reg __403914_403914;
   reg _403915_403915 ; 
   reg __403915_403915;
   reg _403916_403916 ; 
   reg __403916_403916;
   reg _403917_403917 ; 
   reg __403917_403917;
   reg _403918_403918 ; 
   reg __403918_403918;
   reg _403919_403919 ; 
   reg __403919_403919;
   reg _403920_403920 ; 
   reg __403920_403920;
   reg _403921_403921 ; 
   reg __403921_403921;
   reg _403922_403922 ; 
   reg __403922_403922;
   reg _403923_403923 ; 
   reg __403923_403923;
   reg _403924_403924 ; 
   reg __403924_403924;
   reg _403925_403925 ; 
   reg __403925_403925;
   reg _403926_403926 ; 
   reg __403926_403926;
   reg _403927_403927 ; 
   reg __403927_403927;
   reg _403928_403928 ; 
   reg __403928_403928;
   reg _403929_403929 ; 
   reg __403929_403929;
   reg _403930_403930 ; 
   reg __403930_403930;
   reg _403931_403931 ; 
   reg __403931_403931;
   reg _403932_403932 ; 
   reg __403932_403932;
   reg _403933_403933 ; 
   reg __403933_403933;
   reg _403934_403934 ; 
   reg __403934_403934;
   reg _403935_403935 ; 
   reg __403935_403935;
   reg _403936_403936 ; 
   reg __403936_403936;
   reg _403937_403937 ; 
   reg __403937_403937;
   reg _403938_403938 ; 
   reg __403938_403938;
   reg _403939_403939 ; 
   reg __403939_403939;
   reg _403940_403940 ; 
   reg __403940_403940;
   reg _403941_403941 ; 
   reg __403941_403941;
   reg _403942_403942 ; 
   reg __403942_403942;
   reg _403943_403943 ; 
   reg __403943_403943;
   reg _403944_403944 ; 
   reg __403944_403944;
   reg _403945_403945 ; 
   reg __403945_403945;
   reg _403946_403946 ; 
   reg __403946_403946;
   reg _403947_403947 ; 
   reg __403947_403947;
   reg _403948_403948 ; 
   reg __403948_403948;
   reg _403949_403949 ; 
   reg __403949_403949;
   reg _403950_403950 ; 
   reg __403950_403950;
   reg _403951_403951 ; 
   reg __403951_403951;
   reg _403952_403952 ; 
   reg __403952_403952;
   reg _403953_403953 ; 
   reg __403953_403953;
   reg _403954_403954 ; 
   reg __403954_403954;
   reg _403955_403955 ; 
   reg __403955_403955;
   reg _403956_403956 ; 
   reg __403956_403956;
   reg _403957_403957 ; 
   reg __403957_403957;
   reg _403958_403958 ; 
   reg __403958_403958;
   reg _403959_403959 ; 
   reg __403959_403959;
   reg _403960_403960 ; 
   reg __403960_403960;
   reg _403961_403961 ; 
   reg __403961_403961;
   reg _403962_403962 ; 
   reg __403962_403962;
   reg _403963_403963 ; 
   reg __403963_403963;
   reg _403964_403964 ; 
   reg __403964_403964;
   reg _403965_403965 ; 
   reg __403965_403965;
   reg _403966_403966 ; 
   reg __403966_403966;
   reg _403967_403967 ; 
   reg __403967_403967;
   reg _403968_403968 ; 
   reg __403968_403968;
   reg _403969_403969 ; 
   reg __403969_403969;
   reg _403970_403970 ; 
   reg __403970_403970;
   reg _403971_403971 ; 
   reg __403971_403971;
   reg _403972_403972 ; 
   reg __403972_403972;
   reg _403973_403973 ; 
   reg __403973_403973;
   reg _403974_403974 ; 
   reg __403974_403974;
   reg _403975_403975 ; 
   reg __403975_403975;
   reg _403976_403976 ; 
   reg __403976_403976;
   reg _403977_403977 ; 
   reg __403977_403977;
   reg _403978_403978 ; 
   reg __403978_403978;
   reg _403979_403979 ; 
   reg __403979_403979;
   reg _403980_403980 ; 
   reg __403980_403980;
   reg _403981_403981 ; 
   reg __403981_403981;
   reg _403982_403982 ; 
   reg __403982_403982;
   reg _403983_403983 ; 
   reg __403983_403983;
   reg _403984_403984 ; 
   reg __403984_403984;
   reg _403985_403985 ; 
   reg __403985_403985;
   reg _403986_403986 ; 
   reg __403986_403986;
   reg _403987_403987 ; 
   reg __403987_403987;
   reg _403988_403988 ; 
   reg __403988_403988;
   reg _403989_403989 ; 
   reg __403989_403989;
   reg _403990_403990 ; 
   reg __403990_403990;
   reg _403991_403991 ; 
   reg __403991_403991;
   reg _403992_403992 ; 
   reg __403992_403992;
   reg _403993_403993 ; 
   reg __403993_403993;
   reg _403994_403994 ; 
   reg __403994_403994;
   reg _403995_403995 ; 
   reg __403995_403995;
   reg _403996_403996 ; 
   reg __403996_403996;
   reg _403997_403997 ; 
   reg __403997_403997;
   reg _403998_403998 ; 
   reg __403998_403998;
   reg _403999_403999 ; 
   reg __403999_403999;
   reg _404000_404000 ; 
   reg __404000_404000;
   reg _404001_404001 ; 
   reg __404001_404001;
   reg _404002_404002 ; 
   reg __404002_404002;
   reg _404003_404003 ; 
   reg __404003_404003;
   reg _404004_404004 ; 
   reg __404004_404004;
   reg _404005_404005 ; 
   reg __404005_404005;
   reg _404006_404006 ; 
   reg __404006_404006;
   reg _404007_404007 ; 
   reg __404007_404007;
   reg _404008_404008 ; 
   reg __404008_404008;
   reg _404009_404009 ; 
   reg __404009_404009;
   reg _404010_404010 ; 
   reg __404010_404010;
   reg _404011_404011 ; 
   reg __404011_404011;
   reg _404012_404012 ; 
   reg __404012_404012;
   reg _404013_404013 ; 
   reg __404013_404013;
   reg _404014_404014 ; 
   reg __404014_404014;
   reg _404015_404015 ; 
   reg __404015_404015;
   reg _404016_404016 ; 
   reg __404016_404016;
   reg _404017_404017 ; 
   reg __404017_404017;
   reg _404018_404018 ; 
   reg __404018_404018;
   reg _404019_404019 ; 
   reg __404019_404019;
   reg _404020_404020 ; 
   reg __404020_404020;
   reg _404021_404021 ; 
   reg __404021_404021;
   reg _404022_404022 ; 
   reg __404022_404022;
   reg _404023_404023 ; 
   reg __404023_404023;
   reg _404024_404024 ; 
   reg __404024_404024;
   reg _404025_404025 ; 
   reg __404025_404025;
   reg _404026_404026 ; 
   reg __404026_404026;
   reg _404027_404027 ; 
   reg __404027_404027;
   reg _404028_404028 ; 
   reg __404028_404028;
   reg _404029_404029 ; 
   reg __404029_404029;
   reg _404030_404030 ; 
   reg __404030_404030;
   reg _404031_404031 ; 
   reg __404031_404031;
   reg _404032_404032 ; 
   reg __404032_404032;
   reg _404033_404033 ; 
   reg __404033_404033;
   reg _404034_404034 ; 
   reg __404034_404034;
   reg _404035_404035 ; 
   reg __404035_404035;
   reg _404036_404036 ; 
   reg __404036_404036;
   reg _404037_404037 ; 
   reg __404037_404037;
   reg _404038_404038 ; 
   reg __404038_404038;
   reg _404039_404039 ; 
   reg __404039_404039;
   reg _404040_404040 ; 
   reg __404040_404040;
   reg _404041_404041 ; 
   reg __404041_404041;
   reg _404042_404042 ; 
   reg __404042_404042;
   reg _404043_404043 ; 
   reg __404043_404043;
   reg _404044_404044 ; 
   reg __404044_404044;
   reg _404045_404045 ; 
   reg __404045_404045;
   reg _404046_404046 ; 
   reg __404046_404046;
   reg _404047_404047 ; 
   reg __404047_404047;
   reg _404048_404048 ; 
   reg __404048_404048;
   reg _404049_404049 ; 
   reg __404049_404049;
   reg _404050_404050 ; 
   reg __404050_404050;
   reg _404051_404051 ; 
   reg __404051_404051;
   reg _404052_404052 ; 
   reg __404052_404052;
   reg _404053_404053 ; 
   reg __404053_404053;
   reg _404054_404054 ; 
   reg __404054_404054;
   reg _404055_404055 ; 
   reg __404055_404055;
   reg _404056_404056 ; 
   reg __404056_404056;
   reg _404057_404057 ; 
   reg __404057_404057;
   reg _404058_404058 ; 
   reg __404058_404058;
   reg _404059_404059 ; 
   reg __404059_404059;
   reg _404060_404060 ; 
   reg __404060_404060;
   reg _404061_404061 ; 
   reg __404061_404061;
   reg _404062_404062 ; 
   reg __404062_404062;
   reg _404063_404063 ; 
   reg __404063_404063;
   reg _404064_404064 ; 
   reg __404064_404064;
   reg _404065_404065 ; 
   reg __404065_404065;
   reg _404066_404066 ; 
   reg __404066_404066;
   reg _404067_404067 ; 
   reg __404067_404067;
   reg _404068_404068 ; 
   reg __404068_404068;
   reg _404069_404069 ; 
   reg __404069_404069;
   reg _404070_404070 ; 
   reg __404070_404070;
   reg _404071_404071 ; 
   reg __404071_404071;
   reg _404072_404072 ; 
   reg __404072_404072;
   reg _404073_404073 ; 
   reg __404073_404073;
   reg _404074_404074 ; 
   reg __404074_404074;
   reg _404075_404075 ; 
   reg __404075_404075;
   reg _404076_404076 ; 
   reg __404076_404076;
   reg _404077_404077 ; 
   reg __404077_404077;
   reg _404078_404078 ; 
   reg __404078_404078;
   reg _404079_404079 ; 
   reg __404079_404079;
   reg _404080_404080 ; 
   reg __404080_404080;
   reg _404081_404081 ; 
   reg __404081_404081;
   reg _404082_404082 ; 
   reg __404082_404082;
   reg _404083_404083 ; 
   reg __404083_404083;
   reg _404084_404084 ; 
   reg __404084_404084;
   reg _404085_404085 ; 
   reg __404085_404085;
   reg _404086_404086 ; 
   reg __404086_404086;
   reg _404087_404087 ; 
   reg __404087_404087;
   reg _404088_404088 ; 
   reg __404088_404088;
   reg _404089_404089 ; 
   reg __404089_404089;
   reg _404090_404090 ; 
   reg __404090_404090;
   reg _404091_404091 ; 
   reg __404091_404091;
   reg _404092_404092 ; 
   reg __404092_404092;
   reg _404093_404093 ; 
   reg __404093_404093;
   reg _404094_404094 ; 
   reg __404094_404094;
   reg _404095_404095 ; 
   reg __404095_404095;
   reg _404096_404096 ; 
   reg __404096_404096;
   reg _404097_404097 ; 
   reg __404097_404097;
   reg _404098_404098 ; 
   reg __404098_404098;
   reg _404099_404099 ; 
   reg __404099_404099;
   reg _404100_404100 ; 
   reg __404100_404100;
   reg _404101_404101 ; 
   reg __404101_404101;
   reg _404102_404102 ; 
   reg __404102_404102;
   reg _404103_404103 ; 
   reg __404103_404103;
   reg _404104_404104 ; 
   reg __404104_404104;
   reg _404105_404105 ; 
   reg __404105_404105;
   reg _404106_404106 ; 
   reg __404106_404106;
   reg _404107_404107 ; 
   reg __404107_404107;
   reg _404108_404108 ; 
   reg __404108_404108;
   reg _404109_404109 ; 
   reg __404109_404109;
   reg _404110_404110 ; 
   reg __404110_404110;
   reg _404111_404111 ; 
   reg __404111_404111;
   reg _404112_404112 ; 
   reg __404112_404112;
   reg _404113_404113 ; 
   reg __404113_404113;
   reg _404114_404114 ; 
   reg __404114_404114;
   reg _404115_404115 ; 
   reg __404115_404115;
   reg _404116_404116 ; 
   reg __404116_404116;
   reg _404117_404117 ; 
   reg __404117_404117;
   reg _404118_404118 ; 
   reg __404118_404118;
   reg _404119_404119 ; 
   reg __404119_404119;
   reg _404120_404120 ; 
   reg __404120_404120;
   reg _404121_404121 ; 
   reg __404121_404121;
   reg _404122_404122 ; 
   reg __404122_404122;
   reg _404123_404123 ; 
   reg __404123_404123;
   reg _404124_404124 ; 
   reg __404124_404124;
   reg _404125_404125 ; 
   reg __404125_404125;
   reg _404126_404126 ; 
   reg __404126_404126;
   reg _404127_404127 ; 
   reg __404127_404127;
   reg _404128_404128 ; 
   reg __404128_404128;
   reg _404129_404129 ; 
   reg __404129_404129;
   reg _404130_404130 ; 
   reg __404130_404130;
   reg _404131_404131 ; 
   reg __404131_404131;
   reg _404132_404132 ; 
   reg __404132_404132;
   reg _404133_404133 ; 
   reg __404133_404133;
   reg _404134_404134 ; 
   reg __404134_404134;
   reg _404135_404135 ; 
   reg __404135_404135;
   reg _404136_404136 ; 
   reg __404136_404136;
   reg _404137_404137 ; 
   reg __404137_404137;
   reg _404138_404138 ; 
   reg __404138_404138;
   reg _404139_404139 ; 
   reg __404139_404139;
   reg _404140_404140 ; 
   reg __404140_404140;
   reg _404141_404141 ; 
   reg __404141_404141;
   reg _404142_404142 ; 
   reg __404142_404142;
   reg _404143_404143 ; 
   reg __404143_404143;
   reg _404144_404144 ; 
   reg __404144_404144;
   reg _404145_404145 ; 
   reg __404145_404145;
   reg _404146_404146 ; 
   reg __404146_404146;
   reg _404147_404147 ; 
   reg __404147_404147;
   reg _404148_404148 ; 
   reg __404148_404148;
   reg _404149_404149 ; 
   reg __404149_404149;
   reg _404150_404150 ; 
   reg __404150_404150;
   reg _404151_404151 ; 
   reg __404151_404151;
   reg _404152_404152 ; 
   reg __404152_404152;
   reg _404153_404153 ; 
   reg __404153_404153;
   reg _404154_404154 ; 
   reg __404154_404154;
   reg _404155_404155 ; 
   reg __404155_404155;
   reg _404156_404156 ; 
   reg __404156_404156;
   reg _404157_404157 ; 
   reg __404157_404157;
   reg _404158_404158 ; 
   reg __404158_404158;
   reg _404159_404159 ; 
   reg __404159_404159;
   reg _404160_404160 ; 
   reg __404160_404160;
   reg _404161_404161 ; 
   reg __404161_404161;
   reg _404162_404162 ; 
   reg __404162_404162;
   reg _404163_404163 ; 
   reg __404163_404163;
   reg _404164_404164 ; 
   reg __404164_404164;
   reg _404165_404165 ; 
   reg __404165_404165;
   reg _404166_404166 ; 
   reg __404166_404166;
   reg _404167_404167 ; 
   reg __404167_404167;
   reg _404168_404168 ; 
   reg __404168_404168;
   reg _404169_404169 ; 
   reg __404169_404169;
   reg _404170_404170 ; 
   reg __404170_404170;
   reg _404171_404171 ; 
   reg __404171_404171;
   reg _404172_404172 ; 
   reg __404172_404172;
   reg _404173_404173 ; 
   reg __404173_404173;
   reg _404174_404174 ; 
   reg __404174_404174;
   reg _404175_404175 ; 
   reg __404175_404175;
   reg _404176_404176 ; 
   reg __404176_404176;
   reg _404177_404177 ; 
   reg __404177_404177;
   reg _404178_404178 ; 
   reg __404178_404178;
   reg _404179_404179 ; 
   reg __404179_404179;
   reg _404180_404180 ; 
   reg __404180_404180;
   reg _404181_404181 ; 
   reg __404181_404181;
   reg _404182_404182 ; 
   reg __404182_404182;
   reg _404183_404183 ; 
   reg __404183_404183;
   reg _404184_404184 ; 
   reg __404184_404184;
   reg _404185_404185 ; 
   reg __404185_404185;
   reg _404186_404186 ; 
   reg __404186_404186;
   reg _404187_404187 ; 
   reg __404187_404187;
   reg _404188_404188 ; 
   reg __404188_404188;
   reg _404189_404189 ; 
   reg __404189_404189;
   reg _404190_404190 ; 
   reg __404190_404190;
   reg _404191_404191 ; 
   reg __404191_404191;
   reg _404192_404192 ; 
   reg __404192_404192;
   reg _404193_404193 ; 
   reg __404193_404193;
   reg _404194_404194 ; 
   reg __404194_404194;
   reg _404195_404195 ; 
   reg __404195_404195;
   reg _404196_404196 ; 
   reg __404196_404196;
   reg _404197_404197 ; 
   reg __404197_404197;
   reg _404198_404198 ; 
   reg __404198_404198;
   reg _404199_404199 ; 
   reg __404199_404199;
   reg _404200_404200 ; 
   reg __404200_404200;
   reg _404201_404201 ; 
   reg __404201_404201;
   reg _404202_404202 ; 
   reg __404202_404202;
   reg _404203_404203 ; 
   reg __404203_404203;
   reg _404204_404204 ; 
   reg __404204_404204;
   reg _404205_404205 ; 
   reg __404205_404205;
   reg _404206_404206 ; 
   reg __404206_404206;
   reg _404207_404207 ; 
   reg __404207_404207;
   reg _404208_404208 ; 
   reg __404208_404208;
   reg _404209_404209 ; 
   reg __404209_404209;
   reg _404210_404210 ; 
   reg __404210_404210;
   reg _404211_404211 ; 
   reg __404211_404211;
   reg _404212_404212 ; 
   reg __404212_404212;
   reg _404213_404213 ; 
   reg __404213_404213;
   reg _404214_404214 ; 
   reg __404214_404214;
   reg _404215_404215 ; 
   reg __404215_404215;
   reg _404216_404216 ; 
   reg __404216_404216;
   reg _404217_404217 ; 
   reg __404217_404217;
   reg _404218_404218 ; 
   reg __404218_404218;
   reg _404219_404219 ; 
   reg __404219_404219;
   reg _404220_404220 ; 
   reg __404220_404220;
   reg _404221_404221 ; 
   reg __404221_404221;
   reg _404222_404222 ; 
   reg __404222_404222;
   reg _404223_404223 ; 
   reg __404223_404223;
   reg _404224_404224 ; 
   reg __404224_404224;
   reg _404225_404225 ; 
   reg __404225_404225;
   reg _404226_404226 ; 
   reg __404226_404226;
   reg _404227_404227 ; 
   reg __404227_404227;
   reg _404228_404228 ; 
   reg __404228_404228;
   reg _404229_404229 ; 
   reg __404229_404229;
   reg _404230_404230 ; 
   reg __404230_404230;
   reg _404231_404231 ; 
   reg __404231_404231;
   reg _404232_404232 ; 
   reg __404232_404232;
   reg _404233_404233 ; 
   reg __404233_404233;
   reg _404234_404234 ; 
   reg __404234_404234;
   reg _404235_404235 ; 
   reg __404235_404235;
   reg _404236_404236 ; 
   reg __404236_404236;
   reg _404237_404237 ; 
   reg __404237_404237;
   reg _404238_404238 ; 
   reg __404238_404238;
   reg _404239_404239 ; 
   reg __404239_404239;
   reg _404240_404240 ; 
   reg __404240_404240;
   reg _404241_404241 ; 
   reg __404241_404241;
   reg _404242_404242 ; 
   reg __404242_404242;
   reg _404243_404243 ; 
   reg __404243_404243;
   reg _404244_404244 ; 
   reg __404244_404244;
   reg _404245_404245 ; 
   reg __404245_404245;
   reg _404246_404246 ; 
   reg __404246_404246;
   reg _404247_404247 ; 
   reg __404247_404247;
   reg _404248_404248 ; 
   reg __404248_404248;
   reg _404249_404249 ; 
   reg __404249_404249;
   reg _404250_404250 ; 
   reg __404250_404250;
   reg _404251_404251 ; 
   reg __404251_404251;
   reg _404252_404252 ; 
   reg __404252_404252;
   reg _404253_404253 ; 
   reg __404253_404253;
   reg _404254_404254 ; 
   reg __404254_404254;
   reg _404255_404255 ; 
   reg __404255_404255;
   reg _404256_404256 ; 
   reg __404256_404256;
   reg _404257_404257 ; 
   reg __404257_404257;
   reg _404258_404258 ; 
   reg __404258_404258;
   reg _404259_404259 ; 
   reg __404259_404259;
   reg _404260_404260 ; 
   reg __404260_404260;
   reg _404261_404261 ; 
   reg __404261_404261;
   reg _404262_404262 ; 
   reg __404262_404262;
   reg _404263_404263 ; 
   reg __404263_404263;
   reg _404264_404264 ; 
   reg __404264_404264;
   reg _404265_404265 ; 
   reg __404265_404265;
   reg _404266_404266 ; 
   reg __404266_404266;
   reg _404267_404267 ; 
   reg __404267_404267;
   reg _404268_404268 ; 
   reg __404268_404268;
   reg _404269_404269 ; 
   reg __404269_404269;
   reg _404270_404270 ; 
   reg __404270_404270;
   reg _404271_404271 ; 
   reg __404271_404271;
   reg _404272_404272 ; 
   reg __404272_404272;
   reg _404273_404273 ; 
   reg __404273_404273;
   reg _404274_404274 ; 
   reg __404274_404274;
   reg _404275_404275 ; 
   reg __404275_404275;
   reg _404276_404276 ; 
   reg __404276_404276;
   reg _404277_404277 ; 
   reg __404277_404277;
   reg _404278_404278 ; 
   reg __404278_404278;
   reg _404279_404279 ; 
   reg __404279_404279;
   reg _404280_404280 ; 
   reg __404280_404280;
   reg _404281_404281 ; 
   reg __404281_404281;
   reg _404282_404282 ; 
   reg __404282_404282;
   reg _404283_404283 ; 
   reg __404283_404283;
   reg _404284_404284 ; 
   reg __404284_404284;
   reg _404285_404285 ; 
   reg __404285_404285;
   reg _404286_404286 ; 
   reg __404286_404286;
   reg _404287_404287 ; 
   reg __404287_404287;
   reg _404288_404288 ; 
   reg __404288_404288;
   reg _404289_404289 ; 
   reg __404289_404289;
   reg _404290_404290 ; 
   reg __404290_404290;
   reg _404291_404291 ; 
   reg __404291_404291;
   reg _404292_404292 ; 
   reg __404292_404292;
   reg _404293_404293 ; 
   reg __404293_404293;
   reg _404294_404294 ; 
   reg __404294_404294;
   reg _404295_404295 ; 
   reg __404295_404295;
   reg _404296_404296 ; 
   reg __404296_404296;
   reg _404297_404297 ; 
   reg __404297_404297;
   reg _404298_404298 ; 
   reg __404298_404298;
   reg _404299_404299 ; 
   reg __404299_404299;
   reg _404300_404300 ; 
   reg __404300_404300;
   reg _404301_404301 ; 
   reg __404301_404301;
   reg _404302_404302 ; 
   reg __404302_404302;
   reg _404303_404303 ; 
   reg __404303_404303;
   reg _404304_404304 ; 
   reg __404304_404304;
   reg _404305_404305 ; 
   reg __404305_404305;
   reg _404306_404306 ; 
   reg __404306_404306;
   reg _404307_404307 ; 
   reg __404307_404307;
   reg _404308_404308 ; 
   reg __404308_404308;
   reg _404309_404309 ; 
   reg __404309_404309;
   reg _404310_404310 ; 
   reg __404310_404310;
   reg _404311_404311 ; 
   reg __404311_404311;
   reg _404312_404312 ; 
   reg __404312_404312;
   reg _404313_404313 ; 
   reg __404313_404313;
   reg _404314_404314 ; 
   reg __404314_404314;
   reg _404315_404315 ; 
   reg __404315_404315;
   reg _404316_404316 ; 
   reg __404316_404316;
   reg _404317_404317 ; 
   reg __404317_404317;
   reg _404318_404318 ; 
   reg __404318_404318;
   reg _404319_404319 ; 
   reg __404319_404319;
   reg _404320_404320 ; 
   reg __404320_404320;
   reg _404321_404321 ; 
   reg __404321_404321;
   reg _404322_404322 ; 
   reg __404322_404322;
   reg _404323_404323 ; 
   reg __404323_404323;
   reg _404324_404324 ; 
   reg __404324_404324;
   reg _404325_404325 ; 
   reg __404325_404325;
   reg _404326_404326 ; 
   reg __404326_404326;
   reg _404327_404327 ; 
   reg __404327_404327;
   reg _404328_404328 ; 
   reg __404328_404328;
   reg _404329_404329 ; 
   reg __404329_404329;
   reg _404330_404330 ; 
   reg __404330_404330;
   reg _404331_404331 ; 
   reg __404331_404331;
   reg _404332_404332 ; 
   reg __404332_404332;
   reg _404333_404333 ; 
   reg __404333_404333;
   reg _404334_404334 ; 
   reg __404334_404334;
   reg _404335_404335 ; 
   reg __404335_404335;
   reg _404336_404336 ; 
   reg __404336_404336;
   reg _404337_404337 ; 
   reg __404337_404337;
   reg _404338_404338 ; 
   reg __404338_404338;
   reg _404339_404339 ; 
   reg __404339_404339;
   reg _404340_404340 ; 
   reg __404340_404340;
   reg _404341_404341 ; 
   reg __404341_404341;
   reg _404342_404342 ; 
   reg __404342_404342;
   reg _404343_404343 ; 
   reg __404343_404343;
   reg _404344_404344 ; 
   reg __404344_404344;
   reg _404345_404345 ; 
   reg __404345_404345;
   reg _404346_404346 ; 
   reg __404346_404346;
   reg _404347_404347 ; 
   reg __404347_404347;
   reg _404348_404348 ; 
   reg __404348_404348;
   reg _404349_404349 ; 
   reg __404349_404349;
   reg _404350_404350 ; 
   reg __404350_404350;
   reg _404351_404351 ; 
   reg __404351_404351;
   reg _404352_404352 ; 
   reg __404352_404352;
   reg _404353_404353 ; 
   reg __404353_404353;
   reg _404354_404354 ; 
   reg __404354_404354;
   reg _404355_404355 ; 
   reg __404355_404355;
   reg _404356_404356 ; 
   reg __404356_404356;
   reg _404357_404357 ; 
   reg __404357_404357;
   reg _404358_404358 ; 
   reg __404358_404358;
   reg _404359_404359 ; 
   reg __404359_404359;
   reg _404360_404360 ; 
   reg __404360_404360;
   reg _404361_404361 ; 
   reg __404361_404361;
   reg _404362_404362 ; 
   reg __404362_404362;
   reg _404363_404363 ; 
   reg __404363_404363;
   reg _404364_404364 ; 
   reg __404364_404364;
   reg _404365_404365 ; 
   reg __404365_404365;
   reg _404366_404366 ; 
   reg __404366_404366;
   reg _404367_404367 ; 
   reg __404367_404367;
   reg _404368_404368 ; 
   reg __404368_404368;
   reg _404369_404369 ; 
   reg __404369_404369;
   reg _404370_404370 ; 
   reg __404370_404370;
   reg _404371_404371 ; 
   reg __404371_404371;
   reg _404372_404372 ; 
   reg __404372_404372;
   reg _404373_404373 ; 
   reg __404373_404373;
   reg _404374_404374 ; 
   reg __404374_404374;
   reg _404375_404375 ; 
   reg __404375_404375;
   reg _404376_404376 ; 
   reg __404376_404376;
   reg _404377_404377 ; 
   reg __404377_404377;
   reg _404378_404378 ; 
   reg __404378_404378;
   reg _404379_404379 ; 
   reg __404379_404379;
   reg _404380_404380 ; 
   reg __404380_404380;
   reg _404381_404381 ; 
   reg __404381_404381;
   reg _404382_404382 ; 
   reg __404382_404382;
   reg _404383_404383 ; 
   reg __404383_404383;
   reg _404384_404384 ; 
   reg __404384_404384;
   reg _404385_404385 ; 
   reg __404385_404385;
   reg _404386_404386 ; 
   reg __404386_404386;
   reg _404387_404387 ; 
   reg __404387_404387;
   reg _404388_404388 ; 
   reg __404388_404388;
   reg _404389_404389 ; 
   reg __404389_404389;
   reg _404390_404390 ; 
   reg __404390_404390;
   reg _404391_404391 ; 
   reg __404391_404391;
   reg _404392_404392 ; 
   reg __404392_404392;
   reg _404393_404393 ; 
   reg __404393_404393;
   reg _404394_404394 ; 
   reg __404394_404394;
   reg _404395_404395 ; 
   reg __404395_404395;
   reg _404396_404396 ; 
   reg __404396_404396;
   reg _404397_404397 ; 
   reg __404397_404397;
   reg _404398_404398 ; 
   reg __404398_404398;
   reg _404399_404399 ; 
   reg __404399_404399;
   reg _404400_404400 ; 
   reg __404400_404400;
   reg _404401_404401 ; 
   reg __404401_404401;
   reg _404402_404402 ; 
   reg __404402_404402;
   reg _404403_404403 ; 
   reg __404403_404403;
   reg _404404_404404 ; 
   reg __404404_404404;
   reg _404405_404405 ; 
   reg __404405_404405;
   reg _404406_404406 ; 
   reg __404406_404406;
   reg _404407_404407 ; 
   reg __404407_404407;
   reg _404408_404408 ; 
   reg __404408_404408;
   reg _404409_404409 ; 
   reg __404409_404409;
   reg _404410_404410 ; 
   reg __404410_404410;
   reg _404411_404411 ; 
   reg __404411_404411;
   reg _404412_404412 ; 
   reg __404412_404412;
   reg _404413_404413 ; 
   reg __404413_404413;
   reg _404414_404414 ; 
   reg __404414_404414;
   reg _404415_404415 ; 
   reg __404415_404415;
   reg _404416_404416 ; 
   reg __404416_404416;
   reg _404417_404417 ; 
   reg __404417_404417;
   reg _404418_404418 ; 
   reg __404418_404418;
   reg _404419_404419 ; 
   reg __404419_404419;
   reg _404420_404420 ; 
   reg __404420_404420;
   reg _404421_404421 ; 
   reg __404421_404421;
   reg _404422_404422 ; 
   reg __404422_404422;
   reg _404423_404423 ; 
   reg __404423_404423;
   reg _404424_404424 ; 
   reg __404424_404424;
   reg _404425_404425 ; 
   reg __404425_404425;
   reg _404426_404426 ; 
   reg __404426_404426;
   reg _404427_404427 ; 
   reg __404427_404427;
   reg _404428_404428 ; 
   reg __404428_404428;
   reg _404429_404429 ; 
   reg __404429_404429;
   reg _404430_404430 ; 
   reg __404430_404430;
   reg _404431_404431 ; 
   reg __404431_404431;
   reg _404432_404432 ; 
   reg __404432_404432;
   reg _404433_404433 ; 
   reg __404433_404433;
   reg _404434_404434 ; 
   reg __404434_404434;
   reg _404435_404435 ; 
   reg __404435_404435;
   reg _404436_404436 ; 
   reg __404436_404436;
   reg _404437_404437 ; 
   reg __404437_404437;
   reg _404438_404438 ; 
   reg __404438_404438;
   reg _404439_404439 ; 
   reg __404439_404439;
   reg _404440_404440 ; 
   reg __404440_404440;
   reg _404441_404441 ; 
   reg __404441_404441;
   reg _404442_404442 ; 
   reg __404442_404442;
   reg _404443_404443 ; 
   reg __404443_404443;
   reg _404444_404444 ; 
   reg __404444_404444;
   reg _404445_404445 ; 
   reg __404445_404445;
   reg _404446_404446 ; 
   reg __404446_404446;
   reg _404447_404447 ; 
   reg __404447_404447;
   reg _404448_404448 ; 
   reg __404448_404448;
   reg _404449_404449 ; 
   reg __404449_404449;
   reg _404450_404450 ; 
   reg __404450_404450;
   reg _404451_404451 ; 
   reg __404451_404451;
   reg _404452_404452 ; 
   reg __404452_404452;
   reg _404453_404453 ; 
   reg __404453_404453;
   reg _404454_404454 ; 
   reg __404454_404454;
   reg _404455_404455 ; 
   reg __404455_404455;
   reg _404456_404456 ; 
   reg __404456_404456;
   reg _404457_404457 ; 
   reg __404457_404457;
   reg _404458_404458 ; 
   reg __404458_404458;
   reg _404459_404459 ; 
   reg __404459_404459;
   reg _404460_404460 ; 
   reg __404460_404460;
   reg _404461_404461 ; 
   reg __404461_404461;
   reg _404462_404462 ; 
   reg __404462_404462;
   reg _404463_404463 ; 
   reg __404463_404463;
   reg _404464_404464 ; 
   reg __404464_404464;
   reg _404465_404465 ; 
   reg __404465_404465;
   reg _404466_404466 ; 
   reg __404466_404466;
   reg _404467_404467 ; 
   reg __404467_404467;
   reg _404468_404468 ; 
   reg __404468_404468;
   reg _404469_404469 ; 
   reg __404469_404469;
   reg _404470_404470 ; 
   reg __404470_404470;
   reg _404471_404471 ; 
   reg __404471_404471;
   reg _404472_404472 ; 
   reg __404472_404472;
   reg _404473_404473 ; 
   reg __404473_404473;
   reg _404474_404474 ; 
   reg __404474_404474;
   reg _404475_404475 ; 
   reg __404475_404475;
   reg _404476_404476 ; 
   reg __404476_404476;
   reg _404477_404477 ; 
   reg __404477_404477;
   reg _404478_404478 ; 
   reg __404478_404478;
   reg _404479_404479 ; 
   reg __404479_404479;
   reg _404480_404480 ; 
   reg __404480_404480;
   reg _404481_404481 ; 
   reg __404481_404481;
   reg _404482_404482 ; 
   reg __404482_404482;
   reg _404483_404483 ; 
   reg __404483_404483;
   reg _404484_404484 ; 
   reg __404484_404484;
   reg _404485_404485 ; 
   reg __404485_404485;
   reg _404486_404486 ; 
   reg __404486_404486;
   reg _404487_404487 ; 
   reg __404487_404487;
   reg _404488_404488 ; 
   reg __404488_404488;
   reg _404489_404489 ; 
   reg __404489_404489;
   reg _404490_404490 ; 
   reg __404490_404490;
   reg _404491_404491 ; 
   reg __404491_404491;
   reg _404492_404492 ; 
   reg __404492_404492;
   reg _404493_404493 ; 
   reg __404493_404493;
   reg _404494_404494 ; 
   reg __404494_404494;
   reg _404495_404495 ; 
   reg __404495_404495;
   reg _404496_404496 ; 
   reg __404496_404496;
   reg _404497_404497 ; 
   reg __404497_404497;
   reg _404498_404498 ; 
   reg __404498_404498;
   reg _404499_404499 ; 
   reg __404499_404499;
   reg _404500_404500 ; 
   reg __404500_404500;
   reg _404501_404501 ; 
   reg __404501_404501;
   reg _404502_404502 ; 
   reg __404502_404502;
   reg _404503_404503 ; 
   reg __404503_404503;
   reg _404504_404504 ; 
   reg __404504_404504;
   reg _404505_404505 ; 
   reg __404505_404505;
   reg _404506_404506 ; 
   reg __404506_404506;
   reg _404507_404507 ; 
   reg __404507_404507;
   reg _404508_404508 ; 
   reg __404508_404508;
   reg _404509_404509 ; 
   reg __404509_404509;
   reg _404510_404510 ; 
   reg __404510_404510;
   reg _404511_404511 ; 
   reg __404511_404511;
   reg _404512_404512 ; 
   reg __404512_404512;
   reg _404513_404513 ; 
   reg __404513_404513;
   reg _404514_404514 ; 
   reg __404514_404514;
   reg _404515_404515 ; 
   reg __404515_404515;
   reg _404516_404516 ; 
   reg __404516_404516;
   reg _404517_404517 ; 
   reg __404517_404517;
   reg _404518_404518 ; 
   reg __404518_404518;
   reg _404519_404519 ; 
   reg __404519_404519;
   reg _404520_404520 ; 
   reg __404520_404520;
   reg _404521_404521 ; 
   reg __404521_404521;
   reg _404522_404522 ; 
   reg __404522_404522;
   reg _404523_404523 ; 
   reg __404523_404523;
   reg _404524_404524 ; 
   reg __404524_404524;
   reg _404525_404525 ; 
   reg __404525_404525;
   reg _404526_404526 ; 
   reg __404526_404526;
   reg _404527_404527 ; 
   reg __404527_404527;
   reg _404528_404528 ; 
   reg __404528_404528;
   reg _404529_404529 ; 
   reg __404529_404529;
   reg _404530_404530 ; 
   reg __404530_404530;
   reg _404531_404531 ; 
   reg __404531_404531;
   reg _404532_404532 ; 
   reg __404532_404532;
   reg _404533_404533 ; 
   reg __404533_404533;
   reg _404534_404534 ; 
   reg __404534_404534;
   reg _404535_404535 ; 
   reg __404535_404535;
   reg _404536_404536 ; 
   reg __404536_404536;
   reg _404537_404537 ; 
   reg __404537_404537;
   reg _404538_404538 ; 
   reg __404538_404538;
   reg _404539_404539 ; 
   reg __404539_404539;
   reg _404540_404540 ; 
   reg __404540_404540;
   reg _404541_404541 ; 
   reg __404541_404541;
   reg _404542_404542 ; 
   reg __404542_404542;
   reg _404543_404543 ; 
   reg __404543_404543;
   reg _404544_404544 ; 
   reg __404544_404544;
   reg _404545_404545 ; 
   reg __404545_404545;
   reg _404546_404546 ; 
   reg __404546_404546;
   reg _404547_404547 ; 
   reg __404547_404547;
   reg _404548_404548 ; 
   reg __404548_404548;
   reg _404549_404549 ; 
   reg __404549_404549;
   reg _404550_404550 ; 
   reg __404550_404550;
   reg _404551_404551 ; 
   reg __404551_404551;
   reg _404552_404552 ; 
   reg __404552_404552;
   reg _404553_404553 ; 
   reg __404553_404553;
   reg _404554_404554 ; 
   reg __404554_404554;
   reg _404555_404555 ; 
   reg __404555_404555;
   reg _404556_404556 ; 
   reg __404556_404556;
   reg _404557_404557 ; 
   reg __404557_404557;
   reg _404558_404558 ; 
   reg __404558_404558;
   reg _404559_404559 ; 
   reg __404559_404559;
   reg _404560_404560 ; 
   reg __404560_404560;
   reg _404561_404561 ; 
   reg __404561_404561;
   reg _404562_404562 ; 
   reg __404562_404562;
   reg _404563_404563 ; 
   reg __404563_404563;
   reg _404564_404564 ; 
   reg __404564_404564;
   reg _404565_404565 ; 
   reg __404565_404565;
   reg _404566_404566 ; 
   reg __404566_404566;
   reg _404567_404567 ; 
   reg __404567_404567;
   reg _404568_404568 ; 
   reg __404568_404568;
   reg _404569_404569 ; 
   reg __404569_404569;
   reg _404570_404570 ; 
   reg __404570_404570;
   reg _404571_404571 ; 
   reg __404571_404571;
   reg _404572_404572 ; 
   reg __404572_404572;
   reg _404573_404573 ; 
   reg __404573_404573;
   reg _404574_404574 ; 
   reg __404574_404574;
   reg _404575_404575 ; 
   reg __404575_404575;
   reg _404576_404576 ; 
   reg __404576_404576;
   reg _404577_404577 ; 
   reg __404577_404577;
   reg _404578_404578 ; 
   reg __404578_404578;
   reg _404579_404579 ; 
   reg __404579_404579;
   reg _404580_404580 ; 
   reg __404580_404580;
   reg _404581_404581 ; 
   reg __404581_404581;
   reg _404582_404582 ; 
   reg __404582_404582;
   reg _404583_404583 ; 
   reg __404583_404583;
   reg _404584_404584 ; 
   reg __404584_404584;
   reg _404585_404585 ; 
   reg __404585_404585;
   reg _404586_404586 ; 
   reg __404586_404586;
   reg _404587_404587 ; 
   reg __404587_404587;
   reg _404588_404588 ; 
   reg __404588_404588;
   reg _404589_404589 ; 
   reg __404589_404589;
   reg _404590_404590 ; 
   reg __404590_404590;
   reg _404591_404591 ; 
   reg __404591_404591;
   reg _404592_404592 ; 
   reg __404592_404592;
   reg _404593_404593 ; 
   reg __404593_404593;
   reg _404594_404594 ; 
   reg __404594_404594;
   reg _404595_404595 ; 
   reg __404595_404595;
   reg _404596_404596 ; 
   reg __404596_404596;
   reg _404597_404597 ; 
   reg __404597_404597;
   reg _404598_404598 ; 
   reg __404598_404598;
   reg _404599_404599 ; 
   reg __404599_404599;
   reg _404600_404600 ; 
   reg __404600_404600;
   reg _404601_404601 ; 
   reg __404601_404601;
   reg _404602_404602 ; 
   reg __404602_404602;
   reg _404603_404603 ; 
   reg __404603_404603;
   reg _404604_404604 ; 
   reg __404604_404604;
   reg _404605_404605 ; 
   reg __404605_404605;
   reg _404606_404606 ; 
   reg __404606_404606;
   reg _404607_404607 ; 
   reg __404607_404607;
   reg _404608_404608 ; 
   reg __404608_404608;
   reg _404609_404609 ; 
   reg __404609_404609;
   reg _404610_404610 ; 
   reg __404610_404610;
   reg _404611_404611 ; 
   reg __404611_404611;
   reg _404612_404612 ; 
   reg __404612_404612;
   reg _404613_404613 ; 
   reg __404613_404613;
   reg _404614_404614 ; 
   reg __404614_404614;
   reg _404615_404615 ; 
   reg __404615_404615;
   reg _404616_404616 ; 
   reg __404616_404616;
   reg _404617_404617 ; 
   reg __404617_404617;
   reg _404618_404618 ; 
   reg __404618_404618;
   reg _404619_404619 ; 
   reg __404619_404619;
   reg _404620_404620 ; 
   reg __404620_404620;
   reg _404621_404621 ; 
   reg __404621_404621;
   reg _404622_404622 ; 
   reg __404622_404622;
   reg _404623_404623 ; 
   reg __404623_404623;
   reg _404624_404624 ; 
   reg __404624_404624;
   reg _404625_404625 ; 
   reg __404625_404625;
   reg _404626_404626 ; 
   reg __404626_404626;
   reg _404627_404627 ; 
   reg __404627_404627;
   reg _404628_404628 ; 
   reg __404628_404628;
   reg _404629_404629 ; 
   reg __404629_404629;
   reg _404630_404630 ; 
   reg __404630_404630;
   reg _404631_404631 ; 
   reg __404631_404631;
   reg _404632_404632 ; 
   reg __404632_404632;
   reg _404633_404633 ; 
   reg __404633_404633;
   reg _404634_404634 ; 
   reg __404634_404634;
   reg _404635_404635 ; 
   reg __404635_404635;
   reg _404636_404636 ; 
   reg __404636_404636;
   reg _404637_404637 ; 
   reg __404637_404637;
   reg _404638_404638 ; 
   reg __404638_404638;
   reg _404639_404639 ; 
   reg __404639_404639;
   reg _404640_404640 ; 
   reg __404640_404640;
   reg _404641_404641 ; 
   reg __404641_404641;
   reg _404642_404642 ; 
   reg __404642_404642;
   reg _404643_404643 ; 
   reg __404643_404643;
   reg _404644_404644 ; 
   reg __404644_404644;
   reg _404645_404645 ; 
   reg __404645_404645;
   reg _404646_404646 ; 
   reg __404646_404646;
   reg _404647_404647 ; 
   reg __404647_404647;
   reg _404648_404648 ; 
   reg __404648_404648;
   reg _404649_404649 ; 
   reg __404649_404649;
   reg _404650_404650 ; 
   reg __404650_404650;
   reg _404651_404651 ; 
   reg __404651_404651;
   reg _404652_404652 ; 
   reg __404652_404652;
   reg _404653_404653 ; 
   reg __404653_404653;
   reg _404654_404654 ; 
   reg __404654_404654;
   reg _404655_404655 ; 
   reg __404655_404655;
   reg _404656_404656 ; 
   reg __404656_404656;
   reg _404657_404657 ; 
   reg __404657_404657;
   reg _404658_404658 ; 
   reg __404658_404658;
   reg _404659_404659 ; 
   reg __404659_404659;
   reg _404660_404660 ; 
   reg __404660_404660;
   reg _404661_404661 ; 
   reg __404661_404661;
   reg _404662_404662 ; 
   reg __404662_404662;
   reg _404663_404663 ; 
   reg __404663_404663;
   reg _404664_404664 ; 
   reg __404664_404664;
   reg _404665_404665 ; 
   reg __404665_404665;
   reg _404666_404666 ; 
   reg __404666_404666;
   reg _404667_404667 ; 
   reg __404667_404667;
   reg _404668_404668 ; 
   reg __404668_404668;
   reg _404669_404669 ; 
   reg __404669_404669;
   reg _404670_404670 ; 
   reg __404670_404670;
   reg _404671_404671 ; 
   reg __404671_404671;
   reg _404672_404672 ; 
   reg __404672_404672;
   reg _404673_404673 ; 
   reg __404673_404673;
   reg _404674_404674 ; 
   reg __404674_404674;
   reg _404675_404675 ; 
   reg __404675_404675;
   reg _404676_404676 ; 
   reg __404676_404676;
   reg _404677_404677 ; 
   reg __404677_404677;
   reg _404678_404678 ; 
   reg __404678_404678;
   reg _404679_404679 ; 
   reg __404679_404679;
   reg _404680_404680 ; 
   reg __404680_404680;
   reg _404681_404681 ; 
   reg __404681_404681;
   reg _404682_404682 ; 
   reg __404682_404682;
   reg _404683_404683 ; 
   reg __404683_404683;
   reg _404684_404684 ; 
   reg __404684_404684;
   reg _404685_404685 ; 
   reg __404685_404685;
   reg _404686_404686 ; 
   reg __404686_404686;
   reg _404687_404687 ; 
   reg __404687_404687;
   reg _404688_404688 ; 
   reg __404688_404688;
   reg _404689_404689 ; 
   reg __404689_404689;
   reg _404690_404690 ; 
   reg __404690_404690;
   reg _404691_404691 ; 
   reg __404691_404691;
   reg _404692_404692 ; 
   reg __404692_404692;
   reg _404693_404693 ; 
   reg __404693_404693;
   reg _404694_404694 ; 
   reg __404694_404694;
   reg _404695_404695 ; 
   reg __404695_404695;
   reg _404696_404696 ; 
   reg __404696_404696;
   reg _404697_404697 ; 
   reg __404697_404697;
   reg _404698_404698 ; 
   reg __404698_404698;
   reg _404699_404699 ; 
   reg __404699_404699;
   reg _404700_404700 ; 
   reg __404700_404700;
   reg _404701_404701 ; 
   reg __404701_404701;
   reg _404702_404702 ; 
   reg __404702_404702;
   reg _404703_404703 ; 
   reg __404703_404703;
   reg _404704_404704 ; 
   reg __404704_404704;
   reg _404705_404705 ; 
   reg __404705_404705;
   reg _404706_404706 ; 
   reg __404706_404706;
   reg _404707_404707 ; 
   reg __404707_404707;
   reg _404708_404708 ; 
   reg __404708_404708;
   reg _404709_404709 ; 
   reg __404709_404709;
   reg _404710_404710 ; 
   reg __404710_404710;
   reg _404711_404711 ; 
   reg __404711_404711;
   reg _404712_404712 ; 
   reg __404712_404712;
   reg _404713_404713 ; 
   reg __404713_404713;
   reg _404714_404714 ; 
   reg __404714_404714;
   reg _404715_404715 ; 
   reg __404715_404715;
   reg _404716_404716 ; 
   reg __404716_404716;
   reg _404717_404717 ; 
   reg __404717_404717;
   reg _404718_404718 ; 
   reg __404718_404718;
   reg _404719_404719 ; 
   reg __404719_404719;
   reg _404720_404720 ; 
   reg __404720_404720;
   reg _404721_404721 ; 
   reg __404721_404721;
   reg _404722_404722 ; 
   reg __404722_404722;
   reg _404723_404723 ; 
   reg __404723_404723;
   reg _404724_404724 ; 
   reg __404724_404724;
   reg _404725_404725 ; 
   reg __404725_404725;
   reg _404726_404726 ; 
   reg __404726_404726;
   reg _404727_404727 ; 
   reg __404727_404727;
   reg _404728_404728 ; 
   reg __404728_404728;
   reg _404729_404729 ; 
   reg __404729_404729;
   reg _404730_404730 ; 
   reg __404730_404730;
   reg _404731_404731 ; 
   reg __404731_404731;
   reg _404732_404732 ; 
   reg __404732_404732;
   reg _404733_404733 ; 
   reg __404733_404733;
   reg _404734_404734 ; 
   reg __404734_404734;
   reg _404735_404735 ; 
   reg __404735_404735;
   reg _404736_404736 ; 
   reg __404736_404736;
   reg _404737_404737 ; 
   reg __404737_404737;
   reg _404738_404738 ; 
   reg __404738_404738;
   reg _404739_404739 ; 
   reg __404739_404739;
   reg _404740_404740 ; 
   reg __404740_404740;
   reg _404741_404741 ; 
   reg __404741_404741;
   reg _404742_404742 ; 
   reg __404742_404742;
   reg _404743_404743 ; 
   reg __404743_404743;
   reg _404744_404744 ; 
   reg __404744_404744;
   reg _404745_404745 ; 
   reg __404745_404745;
   reg _404746_404746 ; 
   reg __404746_404746;
   reg _404747_404747 ; 
   reg __404747_404747;
   reg _404748_404748 ; 
   reg __404748_404748;
   reg _404749_404749 ; 
   reg __404749_404749;
   reg _404750_404750 ; 
   reg __404750_404750;
   reg _404751_404751 ; 
   reg __404751_404751;
   reg _404752_404752 ; 
   reg __404752_404752;
   reg _404753_404753 ; 
   reg __404753_404753;
   reg _404754_404754 ; 
   reg __404754_404754;
   reg _404755_404755 ; 
   reg __404755_404755;
   reg _404756_404756 ; 
   reg __404756_404756;
   reg _404757_404757 ; 
   reg __404757_404757;
   reg _404758_404758 ; 
   reg __404758_404758;
   reg _404759_404759 ; 
   reg __404759_404759;
   reg _404760_404760 ; 
   reg __404760_404760;
   reg _404761_404761 ; 
   reg __404761_404761;
   reg _404762_404762 ; 
   reg __404762_404762;
   reg _404763_404763 ; 
   reg __404763_404763;
   reg _404764_404764 ; 
   reg __404764_404764;
   reg _404765_404765 ; 
   reg __404765_404765;
   reg _404766_404766 ; 
   reg __404766_404766;
   reg _404767_404767 ; 
   reg __404767_404767;
   reg _404768_404768 ; 
   reg __404768_404768;
   reg _404769_404769 ; 
   reg __404769_404769;
   reg _404770_404770 ; 
   reg __404770_404770;
   reg _404771_404771 ; 
   reg __404771_404771;
   reg _404772_404772 ; 
   reg __404772_404772;
   reg _404773_404773 ; 
   reg __404773_404773;
   reg _404774_404774 ; 
   reg __404774_404774;
   reg _404775_404775 ; 
   reg __404775_404775;
   reg _404776_404776 ; 
   reg __404776_404776;
   reg _404777_404777 ; 
   reg __404777_404777;
   reg _404778_404778 ; 
   reg __404778_404778;
   reg _404779_404779 ; 
   reg __404779_404779;
   reg _404780_404780 ; 
   reg __404780_404780;
   reg _404781_404781 ; 
   reg __404781_404781;
   reg _404782_404782 ; 
   reg __404782_404782;
   reg _404783_404783 ; 
   reg __404783_404783;
   reg _404784_404784 ; 
   reg __404784_404784;
   reg _404785_404785 ; 
   reg __404785_404785;
   reg _404786_404786 ; 
   reg __404786_404786;
   reg _404787_404787 ; 
   reg __404787_404787;
   reg _404788_404788 ; 
   reg __404788_404788;
   reg _404789_404789 ; 
   reg __404789_404789;
   reg _404790_404790 ; 
   reg __404790_404790;
   reg _404791_404791 ; 
   reg __404791_404791;
   reg _404792_404792 ; 
   reg __404792_404792;
   reg _404793_404793 ; 
   reg __404793_404793;
   reg _404794_404794 ; 
   reg __404794_404794;
   reg _404795_404795 ; 
   reg __404795_404795;
   reg _404796_404796 ; 
   reg __404796_404796;
   reg _404797_404797 ; 
   reg __404797_404797;
   reg _404798_404798 ; 
   reg __404798_404798;
   reg _404799_404799 ; 
   reg __404799_404799;
   reg _404800_404800 ; 
   reg __404800_404800;
   reg _404801_404801 ; 
   reg __404801_404801;
   reg _404802_404802 ; 
   reg __404802_404802;
   reg _404803_404803 ; 
   reg __404803_404803;
   reg _404804_404804 ; 
   reg __404804_404804;
   reg _404805_404805 ; 
   reg __404805_404805;
   reg _404806_404806 ; 
   reg __404806_404806;
   reg _404807_404807 ; 
   reg __404807_404807;
   reg _404808_404808 ; 
   reg __404808_404808;
   reg _404809_404809 ; 
   reg __404809_404809;
   reg _404810_404810 ; 
   reg __404810_404810;
   reg _404811_404811 ; 
   reg __404811_404811;
   reg _404812_404812 ; 
   reg __404812_404812;
   reg _404813_404813 ; 
   reg __404813_404813;
   reg _404814_404814 ; 
   reg __404814_404814;
   reg _404815_404815 ; 
   reg __404815_404815;
   reg _404816_404816 ; 
   reg __404816_404816;
   reg _404817_404817 ; 
   reg __404817_404817;
   reg _404818_404818 ; 
   reg __404818_404818;
   reg _404819_404819 ; 
   reg __404819_404819;
   reg _404820_404820 ; 
   reg __404820_404820;
   reg _404821_404821 ; 
   reg __404821_404821;
   reg _404822_404822 ; 
   reg __404822_404822;
   reg _404823_404823 ; 
   reg __404823_404823;
   reg _404824_404824 ; 
   reg __404824_404824;
   reg _404825_404825 ; 
   reg __404825_404825;
   reg _404826_404826 ; 
   reg __404826_404826;
   reg _404827_404827 ; 
   reg __404827_404827;
   reg _404828_404828 ; 
   reg __404828_404828;
   reg _404829_404829 ; 
   reg __404829_404829;
   reg _404830_404830 ; 
   reg __404830_404830;
   reg _404831_404831 ; 
   reg __404831_404831;
   reg _404832_404832 ; 
   reg __404832_404832;
   reg _404833_404833 ; 
   reg __404833_404833;
   reg _404834_404834 ; 
   reg __404834_404834;
   reg _404835_404835 ; 
   reg __404835_404835;
   reg _404836_404836 ; 
   reg __404836_404836;
   reg _404837_404837 ; 
   reg __404837_404837;
   reg _404838_404838 ; 
   reg __404838_404838;
   reg _404839_404839 ; 
   reg __404839_404839;
   reg _404840_404840 ; 
   reg __404840_404840;
   reg _404841_404841 ; 
   reg __404841_404841;
   reg _404842_404842 ; 
   reg __404842_404842;
   reg _404843_404843 ; 
   reg __404843_404843;
   reg _404844_404844 ; 
   reg __404844_404844;
   reg _404845_404845 ; 
   reg __404845_404845;
   reg _404846_404846 ; 
   reg __404846_404846;
   reg _404847_404847 ; 
   reg __404847_404847;
   reg _404848_404848 ; 
   reg __404848_404848;
   reg _404849_404849 ; 
   reg __404849_404849;
   reg _404850_404850 ; 
   reg __404850_404850;
   reg _404851_404851 ; 
   reg __404851_404851;
   reg _404852_404852 ; 
   reg __404852_404852;
   reg _404853_404853 ; 
   reg __404853_404853;
   reg _404854_404854 ; 
   reg __404854_404854;
   reg _404855_404855 ; 
   reg __404855_404855;
   reg _404856_404856 ; 
   reg __404856_404856;
   reg _404857_404857 ; 
   reg __404857_404857;
   reg _404858_404858 ; 
   reg __404858_404858;
   reg _404859_404859 ; 
   reg __404859_404859;
   reg _404860_404860 ; 
   reg __404860_404860;
   reg _404861_404861 ; 
   reg __404861_404861;
   reg _404862_404862 ; 
   reg __404862_404862;
   reg _404863_404863 ; 
   reg __404863_404863;
   reg _404864_404864 ; 
   reg __404864_404864;
   reg _404865_404865 ; 
   reg __404865_404865;
   reg _404866_404866 ; 
   reg __404866_404866;
   reg _404867_404867 ; 
   reg __404867_404867;
   reg _404868_404868 ; 
   reg __404868_404868;
   reg _404869_404869 ; 
   reg __404869_404869;
   reg _404870_404870 ; 
   reg __404870_404870;
   reg _404871_404871 ; 
   reg __404871_404871;
   reg _404872_404872 ; 
   reg __404872_404872;
   reg _404873_404873 ; 
   reg __404873_404873;
   reg _404874_404874 ; 
   reg __404874_404874;
   reg _404875_404875 ; 
   reg __404875_404875;
   reg _404876_404876 ; 
   reg __404876_404876;
   reg _404877_404877 ; 
   reg __404877_404877;
   reg _404878_404878 ; 
   reg __404878_404878;
   reg _404879_404879 ; 
   reg __404879_404879;
   reg _404880_404880 ; 
   reg __404880_404880;
   reg _404881_404881 ; 
   reg __404881_404881;
   reg _404882_404882 ; 
   reg __404882_404882;
   reg _404883_404883 ; 
   reg __404883_404883;
   reg _404884_404884 ; 
   reg __404884_404884;
   reg _404885_404885 ; 
   reg __404885_404885;
   reg _404886_404886 ; 
   reg __404886_404886;
   reg _404887_404887 ; 
   reg __404887_404887;
   reg _404888_404888 ; 
   reg __404888_404888;
   reg _404889_404889 ; 
   reg __404889_404889;
   reg _404890_404890 ; 
   reg __404890_404890;
   reg _404891_404891 ; 
   reg __404891_404891;
   reg _404892_404892 ; 
   reg __404892_404892;
   reg _404893_404893 ; 
   reg __404893_404893;
   reg _404894_404894 ; 
   reg __404894_404894;
   reg _404895_404895 ; 
   reg __404895_404895;
   reg _404896_404896 ; 
   reg __404896_404896;
   reg _404897_404897 ; 
   reg __404897_404897;
   reg _404898_404898 ; 
   reg __404898_404898;
   reg _404899_404899 ; 
   reg __404899_404899;
   reg _404900_404900 ; 
   reg __404900_404900;
   reg _404901_404901 ; 
   reg __404901_404901;
   reg _404902_404902 ; 
   reg __404902_404902;
   reg _404903_404903 ; 
   reg __404903_404903;
   reg _404904_404904 ; 
   reg __404904_404904;
   reg _404905_404905 ; 
   reg __404905_404905;
   reg _404906_404906 ; 
   reg __404906_404906;
   reg _404907_404907 ; 
   reg __404907_404907;
   reg _404908_404908 ; 
   reg __404908_404908;
   reg _404909_404909 ; 
   reg __404909_404909;
   reg _404910_404910 ; 
   reg __404910_404910;
   reg _404911_404911 ; 
   reg __404911_404911;
   reg _404912_404912 ; 
   reg __404912_404912;
   reg _404913_404913 ; 
   reg __404913_404913;
   reg _404914_404914 ; 
   reg __404914_404914;
   reg _404915_404915 ; 
   reg __404915_404915;
   reg _404916_404916 ; 
   reg __404916_404916;
   reg _404917_404917 ; 
   reg __404917_404917;
   reg _404918_404918 ; 
   reg __404918_404918;
   reg _404919_404919 ; 
   reg __404919_404919;
   reg _404920_404920 ; 
   reg __404920_404920;
   reg _404921_404921 ; 
   reg __404921_404921;
   reg _404922_404922 ; 
   reg __404922_404922;
   reg _404923_404923 ; 
   reg __404923_404923;
   reg _404924_404924 ; 
   reg __404924_404924;
   reg _404925_404925 ; 
   reg __404925_404925;
   reg _404926_404926 ; 
   reg __404926_404926;
   reg _404927_404927 ; 
   reg __404927_404927;
   reg _404928_404928 ; 
   reg __404928_404928;
   reg _404929_404929 ; 
   reg __404929_404929;
   reg _404930_404930 ; 
   reg __404930_404930;
   reg _404931_404931 ; 
   reg __404931_404931;
   reg _404932_404932 ; 
   reg __404932_404932;
   reg _404933_404933 ; 
   reg __404933_404933;
   reg _404934_404934 ; 
   reg __404934_404934;
   reg _404935_404935 ; 
   reg __404935_404935;
   reg _404936_404936 ; 
   reg __404936_404936;
   reg _404937_404937 ; 
   reg __404937_404937;
   reg _404938_404938 ; 
   reg __404938_404938;
   reg _404939_404939 ; 
   reg __404939_404939;
   reg _404940_404940 ; 
   reg __404940_404940;
   reg _404941_404941 ; 
   reg __404941_404941;
   reg _404942_404942 ; 
   reg __404942_404942;
   reg _404943_404943 ; 
   reg __404943_404943;
   reg _404944_404944 ; 
   reg __404944_404944;
   reg _404945_404945 ; 
   reg __404945_404945;
   reg _404946_404946 ; 
   reg __404946_404946;
   reg _404947_404947 ; 
   reg __404947_404947;
   reg _404948_404948 ; 
   reg __404948_404948;
   reg _404949_404949 ; 
   reg __404949_404949;
   reg _404950_404950 ; 
   reg __404950_404950;
   reg _404951_404951 ; 
   reg __404951_404951;
   reg _404952_404952 ; 
   reg __404952_404952;
   reg _404953_404953 ; 
   reg __404953_404953;
   reg _404954_404954 ; 
   reg __404954_404954;
   reg _404955_404955 ; 
   reg __404955_404955;
   reg _404956_404956 ; 
   reg __404956_404956;
   reg _404957_404957 ; 
   reg __404957_404957;
   reg _404958_404958 ; 
   reg __404958_404958;
   reg _404959_404959 ; 
   reg __404959_404959;
   reg _404960_404960 ; 
   reg __404960_404960;
   reg _404961_404961 ; 
   reg __404961_404961;
   reg _404962_404962 ; 
   reg __404962_404962;
   reg _404963_404963 ; 
   reg __404963_404963;
   reg _404964_404964 ; 
   reg __404964_404964;
   reg _404965_404965 ; 
   reg __404965_404965;
   reg _404966_404966 ; 
   reg __404966_404966;
   reg _404967_404967 ; 
   reg __404967_404967;
   reg _404968_404968 ; 
   reg __404968_404968;
   reg _404969_404969 ; 
   reg __404969_404969;
   reg _404970_404970 ; 
   reg __404970_404970;
   reg _404971_404971 ; 
   reg __404971_404971;
   reg _404972_404972 ; 
   reg __404972_404972;
   reg _404973_404973 ; 
   reg __404973_404973;
   reg _404974_404974 ; 
   reg __404974_404974;
   reg _404975_404975 ; 
   reg __404975_404975;
   reg _404976_404976 ; 
   reg __404976_404976;
   reg _404977_404977 ; 
   reg __404977_404977;
   reg _404978_404978 ; 
   reg __404978_404978;
   reg _404979_404979 ; 
   reg __404979_404979;
   reg _404980_404980 ; 
   reg __404980_404980;
   reg _404981_404981 ; 
   reg __404981_404981;
   reg _404982_404982 ; 
   reg __404982_404982;
   reg _404983_404983 ; 
   reg __404983_404983;
   reg _404984_404984 ; 
   reg __404984_404984;
   reg _404985_404985 ; 
   reg __404985_404985;
   reg _404986_404986 ; 
   reg __404986_404986;
   reg _404987_404987 ; 
   reg __404987_404987;
   reg _404988_404988 ; 
   reg __404988_404988;
   reg _404989_404989 ; 
   reg __404989_404989;
   reg _404990_404990 ; 
   reg __404990_404990;
   reg _404991_404991 ; 
   reg __404991_404991;
   reg _404992_404992 ; 
   reg __404992_404992;
   reg _404993_404993 ; 
   reg __404993_404993;
   reg _404994_404994 ; 
   reg __404994_404994;
   reg _404995_404995 ; 
   reg __404995_404995;
   reg _404996_404996 ; 
   reg __404996_404996;
   reg _404997_404997 ; 
   reg __404997_404997;
   reg _404998_404998 ; 
   reg __404998_404998;
   reg _404999_404999 ; 
   reg __404999_404999;
   reg _405000_405000 ; 
   reg __405000_405000;
   reg _405001_405001 ; 
   reg __405001_405001;
   reg _405002_405002 ; 
   reg __405002_405002;
   reg _405003_405003 ; 
   reg __405003_405003;
   reg _405004_405004 ; 
   reg __405004_405004;
   reg _405005_405005 ; 
   reg __405005_405005;
   reg _405006_405006 ; 
   reg __405006_405006;
   reg _405007_405007 ; 
   reg __405007_405007;
   reg _405008_405008 ; 
   reg __405008_405008;
   reg _405009_405009 ; 
   reg __405009_405009;
   reg _405010_405010 ; 
   reg __405010_405010;
   reg _405011_405011 ; 
   reg __405011_405011;
   reg _405012_405012 ; 
   reg __405012_405012;
   reg _405013_405013 ; 
   reg __405013_405013;
   reg _405014_405014 ; 
   reg __405014_405014;
   reg _405015_405015 ; 
   reg __405015_405015;
   reg _405016_405016 ; 
   reg __405016_405016;
   reg _405017_405017 ; 
   reg __405017_405017;
   reg _405018_405018 ; 
   reg __405018_405018;
   reg _405019_405019 ; 
   reg __405019_405019;
   reg _405020_405020 ; 
   reg __405020_405020;
   reg _405021_405021 ; 
   reg __405021_405021;
   reg _405022_405022 ; 
   reg __405022_405022;
   reg _405023_405023 ; 
   reg __405023_405023;
   reg _405024_405024 ; 
   reg __405024_405024;
   reg _405025_405025 ; 
   reg __405025_405025;
   reg _405026_405026 ; 
   reg __405026_405026;
   reg _405027_405027 ; 
   reg __405027_405027;
   reg _405028_405028 ; 
   reg __405028_405028;
   reg _405029_405029 ; 
   reg __405029_405029;
   reg _405030_405030 ; 
   reg __405030_405030;
   reg _405031_405031 ; 
   reg __405031_405031;
   reg _405032_405032 ; 
   reg __405032_405032;
   reg _405033_405033 ; 
   reg __405033_405033;
   reg _405034_405034 ; 
   reg __405034_405034;
   reg _405035_405035 ; 
   reg __405035_405035;
   reg _405036_405036 ; 
   reg __405036_405036;
   reg _405037_405037 ; 
   reg __405037_405037;
   reg _405038_405038 ; 
   reg __405038_405038;
   reg _405039_405039 ; 
   reg __405039_405039;
   reg _405040_405040 ; 
   reg __405040_405040;
   reg _405041_405041 ; 
   reg __405041_405041;
   reg _405042_405042 ; 
   reg __405042_405042;
   reg _405043_405043 ; 
   reg __405043_405043;
   reg _405044_405044 ; 
   reg __405044_405044;
   reg _405045_405045 ; 
   reg __405045_405045;
   reg _405046_405046 ; 
   reg __405046_405046;
   reg _405047_405047 ; 
   reg __405047_405047;
   reg _405048_405048 ; 
   reg __405048_405048;
   reg _405049_405049 ; 
   reg __405049_405049;
   reg _405050_405050 ; 
   reg __405050_405050;
   reg _405051_405051 ; 
   reg __405051_405051;
   reg _405052_405052 ; 
   reg __405052_405052;
   reg _405053_405053 ; 
   reg __405053_405053;
   reg _405054_405054 ; 
   reg __405054_405054;
   reg _405055_405055 ; 
   reg __405055_405055;
   reg _405056_405056 ; 
   reg __405056_405056;
   reg _405057_405057 ; 
   reg __405057_405057;
   reg _405058_405058 ; 
   reg __405058_405058;
   reg _405059_405059 ; 
   reg __405059_405059;
   reg _405060_405060 ; 
   reg __405060_405060;
   reg _405061_405061 ; 
   reg __405061_405061;
   reg _405062_405062 ; 
   reg __405062_405062;
   reg _405063_405063 ; 
   reg __405063_405063;
   reg _405064_405064 ; 
   reg __405064_405064;
   reg _405065_405065 ; 
   reg __405065_405065;
   reg _405066_405066 ; 
   reg __405066_405066;
   reg _405067_405067 ; 
   reg __405067_405067;
   reg _405068_405068 ; 
   reg __405068_405068;
   reg _405069_405069 ; 
   reg __405069_405069;
   reg _405070_405070 ; 
   reg __405070_405070;
   reg _405071_405071 ; 
   reg __405071_405071;
   reg _405072_405072 ; 
   reg __405072_405072;
   reg _405073_405073 ; 
   reg __405073_405073;
   reg _405074_405074 ; 
   reg __405074_405074;
   reg _405075_405075 ; 
   reg __405075_405075;
   reg _405076_405076 ; 
   reg __405076_405076;
   reg _405077_405077 ; 
   reg __405077_405077;
   reg _405078_405078 ; 
   reg __405078_405078;
   reg _405079_405079 ; 
   reg __405079_405079;
   reg _405080_405080 ; 
   reg __405080_405080;
   reg _405081_405081 ; 
   reg __405081_405081;
   reg _405082_405082 ; 
   reg __405082_405082;
   reg _405083_405083 ; 
   reg __405083_405083;
   reg _405084_405084 ; 
   reg __405084_405084;
   reg _405085_405085 ; 
   reg __405085_405085;
   reg _405086_405086 ; 
   reg __405086_405086;
   reg _405087_405087 ; 
   reg __405087_405087;
   reg _405088_405088 ; 
   reg __405088_405088;
   reg _405089_405089 ; 
   reg __405089_405089;
   reg _405090_405090 ; 
   reg __405090_405090;
   reg _405091_405091 ; 
   reg __405091_405091;
   reg _405092_405092 ; 
   reg __405092_405092;
   reg _405093_405093 ; 
   reg __405093_405093;
   reg _405094_405094 ; 
   reg __405094_405094;
   reg _405095_405095 ; 
   reg __405095_405095;
   reg _405096_405096 ; 
   reg __405096_405096;
   reg _405097_405097 ; 
   reg __405097_405097;
   reg _405098_405098 ; 
   reg __405098_405098;
   reg _405099_405099 ; 
   reg __405099_405099;
   reg _405100_405100 ; 
   reg __405100_405100;
   reg _405101_405101 ; 
   reg __405101_405101;
   reg _405102_405102 ; 
   reg __405102_405102;
   reg _405103_405103 ; 
   reg __405103_405103;
   reg _405104_405104 ; 
   reg __405104_405104;
   reg _405105_405105 ; 
   reg __405105_405105;
   reg _405106_405106 ; 
   reg __405106_405106;
   reg _405107_405107 ; 
   reg __405107_405107;
   reg _405108_405108 ; 
   reg __405108_405108;
   reg _405109_405109 ; 
   reg __405109_405109;
   reg _405110_405110 ; 
   reg __405110_405110;
   reg _405111_405111 ; 
   reg __405111_405111;
   reg _405112_405112 ; 
   reg __405112_405112;
   reg _405113_405113 ; 
   reg __405113_405113;
   reg _405114_405114 ; 
   reg __405114_405114;
   reg _405115_405115 ; 
   reg __405115_405115;
   reg _405116_405116 ; 
   reg __405116_405116;
   reg _405117_405117 ; 
   reg __405117_405117;
   reg _405118_405118 ; 
   reg __405118_405118;
   reg _405119_405119 ; 
   reg __405119_405119;
   reg _405120_405120 ; 
   reg __405120_405120;
   reg _405121_405121 ; 
   reg __405121_405121;
   reg _405122_405122 ; 
   reg __405122_405122;
   reg _405123_405123 ; 
   reg __405123_405123;
   reg _405124_405124 ; 
   reg __405124_405124;
   reg _405125_405125 ; 
   reg __405125_405125;
   reg _405126_405126 ; 
   reg __405126_405126;
   reg _405127_405127 ; 
   reg __405127_405127;
   reg _405128_405128 ; 
   reg __405128_405128;
   reg _405129_405129 ; 
   reg __405129_405129;
   reg _405130_405130 ; 
   reg __405130_405130;
   reg _405131_405131 ; 
   reg __405131_405131;
   reg _405132_405132 ; 
   reg __405132_405132;
   reg _405133_405133 ; 
   reg __405133_405133;
   reg _405134_405134 ; 
   reg __405134_405134;
   reg _405135_405135 ; 
   reg __405135_405135;
   reg _405136_405136 ; 
   reg __405136_405136;
   reg _405137_405137 ; 
   reg __405137_405137;
   reg _405138_405138 ; 
   reg __405138_405138;
   reg _405139_405139 ; 
   reg __405139_405139;
   reg _405140_405140 ; 
   reg __405140_405140;
   reg _405141_405141 ; 
   reg __405141_405141;
   reg _405142_405142 ; 
   reg __405142_405142;
   reg _405143_405143 ; 
   reg __405143_405143;
   reg _405144_405144 ; 
   reg __405144_405144;
   reg _405145_405145 ; 
   reg __405145_405145;
   reg _405146_405146 ; 
   reg __405146_405146;
   reg _405147_405147 ; 
   reg __405147_405147;
   reg _405148_405148 ; 
   reg __405148_405148;
   reg _405149_405149 ; 
   reg __405149_405149;
   reg _405150_405150 ; 
   reg __405150_405150;
   reg _405151_405151 ; 
   reg __405151_405151;
   reg _405152_405152 ; 
   reg __405152_405152;
   reg _405153_405153 ; 
   reg __405153_405153;
   reg _405154_405154 ; 
   reg __405154_405154;
   reg _405155_405155 ; 
   reg __405155_405155;
   reg _405156_405156 ; 
   reg __405156_405156;
   reg _405157_405157 ; 
   reg __405157_405157;
   reg _405158_405158 ; 
   reg __405158_405158;
   reg _405159_405159 ; 
   reg __405159_405159;
   reg _405160_405160 ; 
   reg __405160_405160;
   reg _405161_405161 ; 
   reg __405161_405161;
   reg _405162_405162 ; 
   reg __405162_405162;
   reg _405163_405163 ; 
   reg __405163_405163;
   reg _405164_405164 ; 
   reg __405164_405164;
   reg _405165_405165 ; 
   reg __405165_405165;
   reg _405166_405166 ; 
   reg __405166_405166;
   reg _405167_405167 ; 
   reg __405167_405167;
   reg _405168_405168 ; 
   reg __405168_405168;
   reg _405169_405169 ; 
   reg __405169_405169;
   reg _405170_405170 ; 
   reg __405170_405170;
   reg _405171_405171 ; 
   reg __405171_405171;
   reg _405172_405172 ; 
   reg __405172_405172;
   reg _405173_405173 ; 
   reg __405173_405173;
   reg _405174_405174 ; 
   reg __405174_405174;
   reg _405175_405175 ; 
   reg __405175_405175;
   reg _405176_405176 ; 
   reg __405176_405176;
   reg _405177_405177 ; 
   reg __405177_405177;
   reg _405178_405178 ; 
   reg __405178_405178;
   reg _405179_405179 ; 
   reg __405179_405179;
   reg _405180_405180 ; 
   reg __405180_405180;
   reg _405181_405181 ; 
   reg __405181_405181;
   reg _405182_405182 ; 
   reg __405182_405182;
   reg _405183_405183 ; 
   reg __405183_405183;
   reg _405184_405184 ; 
   reg __405184_405184;
   reg _405185_405185 ; 
   reg __405185_405185;
   reg _405186_405186 ; 
   reg __405186_405186;
   reg _405187_405187 ; 
   reg __405187_405187;
   reg _405188_405188 ; 
   reg __405188_405188;
   reg _405189_405189 ; 
   reg __405189_405189;
   reg _405190_405190 ; 
   reg __405190_405190;
   reg _405191_405191 ; 
   reg __405191_405191;
   reg _405192_405192 ; 
   reg __405192_405192;
   reg _405193_405193 ; 
   reg __405193_405193;
   reg _405194_405194 ; 
   reg __405194_405194;
   reg _405195_405195 ; 
   reg __405195_405195;
   reg _405196_405196 ; 
   reg __405196_405196;
   reg _405197_405197 ; 
   reg __405197_405197;
   reg _405198_405198 ; 
   reg __405198_405198;
   reg _405199_405199 ; 
   reg __405199_405199;
   reg _405200_405200 ; 
   reg __405200_405200;
   reg _405201_405201 ; 
   reg __405201_405201;
   reg _405202_405202 ; 
   reg __405202_405202;
   reg _405203_405203 ; 
   reg __405203_405203;
   reg _405204_405204 ; 
   reg __405204_405204;
   reg _405205_405205 ; 
   reg __405205_405205;
   reg _405206_405206 ; 
   reg __405206_405206;
   reg _405207_405207 ; 
   reg __405207_405207;
   reg _405208_405208 ; 
   reg __405208_405208;
   reg _405209_405209 ; 
   reg __405209_405209;
   reg _405210_405210 ; 
   reg __405210_405210;
   reg _405211_405211 ; 
   reg __405211_405211;
   reg _405212_405212 ; 
   reg __405212_405212;
   reg _405213_405213 ; 
   reg __405213_405213;
   reg _405214_405214 ; 
   reg __405214_405214;
   reg _405215_405215 ; 
   reg __405215_405215;
   reg _405216_405216 ; 
   reg __405216_405216;
   reg _405217_405217 ; 
   reg __405217_405217;
   reg _405218_405218 ; 
   reg __405218_405218;
   reg _405219_405219 ; 
   reg __405219_405219;
   reg _405220_405220 ; 
   reg __405220_405220;
   reg _405221_405221 ; 
   reg __405221_405221;
   reg _405222_405222 ; 
   reg __405222_405222;
   reg _405223_405223 ; 
   reg __405223_405223;
   reg _405224_405224 ; 
   reg __405224_405224;
   reg _405225_405225 ; 
   reg __405225_405225;
   reg _405226_405226 ; 
   reg __405226_405226;
   reg _405227_405227 ; 
   reg __405227_405227;
   reg _405228_405228 ; 
   reg __405228_405228;
   reg _405229_405229 ; 
   reg __405229_405229;
   reg _405230_405230 ; 
   reg __405230_405230;
   reg _405231_405231 ; 
   reg __405231_405231;
   reg _405232_405232 ; 
   reg __405232_405232;
   reg _405233_405233 ; 
   reg __405233_405233;
   reg _405234_405234 ; 
   reg __405234_405234;
   reg _405235_405235 ; 
   reg __405235_405235;
   reg _405236_405236 ; 
   reg __405236_405236;
   reg _405237_405237 ; 
   reg __405237_405237;
   reg _405238_405238 ; 
   reg __405238_405238;
   reg _405239_405239 ; 
   reg __405239_405239;
   reg _405240_405240 ; 
   reg __405240_405240;
   reg _405241_405241 ; 
   reg __405241_405241;
   reg _405242_405242 ; 
   reg __405242_405242;
   reg _405243_405243 ; 
   reg __405243_405243;
   reg _405244_405244 ; 
   reg __405244_405244;
   reg _405245_405245 ; 
   reg __405245_405245;
   reg _405246_405246 ; 
   reg __405246_405246;
   reg _405247_405247 ; 
   reg __405247_405247;
   reg _405248_405248 ; 
   reg __405248_405248;
   reg _405249_405249 ; 
   reg __405249_405249;
   reg _405250_405250 ; 
   reg __405250_405250;
   reg _405251_405251 ; 
   reg __405251_405251;
   reg _405252_405252 ; 
   reg __405252_405252;
   reg _405253_405253 ; 
   reg __405253_405253;
   reg _405254_405254 ; 
   reg __405254_405254;
   reg _405255_405255 ; 
   reg __405255_405255;
   reg _405256_405256 ; 
   reg __405256_405256;
   reg _405257_405257 ; 
   reg __405257_405257;
   reg _405258_405258 ; 
   reg __405258_405258;
   reg _405259_405259 ; 
   reg __405259_405259;
   reg _405260_405260 ; 
   reg __405260_405260;
   reg _405261_405261 ; 
   reg __405261_405261;
   reg _405262_405262 ; 
   reg __405262_405262;
   reg _405263_405263 ; 
   reg __405263_405263;
   reg _405264_405264 ; 
   reg __405264_405264;
   reg _405265_405265 ; 
   reg __405265_405265;
   reg _405266_405266 ; 
   reg __405266_405266;
   reg _405267_405267 ; 
   reg __405267_405267;
   reg _405268_405268 ; 
   reg __405268_405268;
   reg _405269_405269 ; 
   reg __405269_405269;
   reg _405270_405270 ; 
   reg __405270_405270;
   reg _405271_405271 ; 
   reg __405271_405271;
   reg _405272_405272 ; 
   reg __405272_405272;
   reg _405273_405273 ; 
   reg __405273_405273;
   reg _405274_405274 ; 
   reg __405274_405274;
   reg _405275_405275 ; 
   reg __405275_405275;
   reg _405276_405276 ; 
   reg __405276_405276;
   reg _405277_405277 ; 
   reg __405277_405277;
   reg _405278_405278 ; 
   reg __405278_405278;
   reg _405279_405279 ; 
   reg __405279_405279;
   reg _405280_405280 ; 
   reg __405280_405280;
   reg _405281_405281 ; 
   reg __405281_405281;
   reg _405282_405282 ; 
   reg __405282_405282;
   reg _405283_405283 ; 
   reg __405283_405283;
   reg _405284_405284 ; 
   reg __405284_405284;
   reg _405285_405285 ; 
   reg __405285_405285;
   reg _405286_405286 ; 
   reg __405286_405286;
   reg _405287_405287 ; 
   reg __405287_405287;
   reg _405288_405288 ; 
   reg __405288_405288;
   reg _405289_405289 ; 
   reg __405289_405289;
   reg _405290_405290 ; 
   reg __405290_405290;
   reg _405291_405291 ; 
   reg __405291_405291;
   reg _405292_405292 ; 
   reg __405292_405292;
   reg _405293_405293 ; 
   reg __405293_405293;
   reg _405294_405294 ; 
   reg __405294_405294;
   reg _405295_405295 ; 
   reg __405295_405295;
   reg _405296_405296 ; 
   reg __405296_405296;
   reg _405297_405297 ; 
   reg __405297_405297;
   reg _405298_405298 ; 
   reg __405298_405298;
   reg _405299_405299 ; 
   reg __405299_405299;
   reg _405300_405300 ; 
   reg __405300_405300;
   reg _405301_405301 ; 
   reg __405301_405301;
   reg _405302_405302 ; 
   reg __405302_405302;
   reg _405303_405303 ; 
   reg __405303_405303;
   reg _405304_405304 ; 
   reg __405304_405304;
   reg _405305_405305 ; 
   reg __405305_405305;
   reg _405306_405306 ; 
   reg __405306_405306;
   reg _405307_405307 ; 
   reg __405307_405307;
   reg _405308_405308 ; 
   reg __405308_405308;
   reg _405309_405309 ; 
   reg __405309_405309;
   reg _405310_405310 ; 
   reg __405310_405310;
   reg _405311_405311 ; 
   reg __405311_405311;
   reg _405312_405312 ; 
   reg __405312_405312;
   reg _405313_405313 ; 
   reg __405313_405313;
   reg _405314_405314 ; 
   reg __405314_405314;
   reg _405315_405315 ; 
   reg __405315_405315;
   reg _405316_405316 ; 
   reg __405316_405316;
   reg _405317_405317 ; 
   reg __405317_405317;
   reg _405318_405318 ; 
   reg __405318_405318;
   reg _405319_405319 ; 
   reg __405319_405319;
   reg _405320_405320 ; 
   reg __405320_405320;
   reg _405321_405321 ; 
   reg __405321_405321;
   reg _405322_405322 ; 
   reg __405322_405322;
   reg _405323_405323 ; 
   reg __405323_405323;
   reg _405324_405324 ; 
   reg __405324_405324;
   reg _405325_405325 ; 
   reg __405325_405325;
   reg _405326_405326 ; 
   reg __405326_405326;
   reg _405327_405327 ; 
   reg __405327_405327;
   reg _405328_405328 ; 
   reg __405328_405328;
   reg _405329_405329 ; 
   reg __405329_405329;
   reg _405330_405330 ; 
   reg __405330_405330;
   reg _405331_405331 ; 
   reg __405331_405331;
   reg _405332_405332 ; 
   reg __405332_405332;
   reg _405333_405333 ; 
   reg __405333_405333;
   reg _405334_405334 ; 
   reg __405334_405334;
   reg _405335_405335 ; 
   reg __405335_405335;
   reg _405336_405336 ; 
   reg __405336_405336;
   reg _405337_405337 ; 
   reg __405337_405337;
   reg _405338_405338 ; 
   reg __405338_405338;
   reg _405339_405339 ; 
   reg __405339_405339;
   reg _405340_405340 ; 
   reg __405340_405340;
   reg _405341_405341 ; 
   reg __405341_405341;
   reg _405342_405342 ; 
   reg __405342_405342;
   reg _405343_405343 ; 
   reg __405343_405343;
   reg _405344_405344 ; 
   reg __405344_405344;
   reg _405345_405345 ; 
   reg __405345_405345;
   reg _405346_405346 ; 
   reg __405346_405346;
   reg _405347_405347 ; 
   reg __405347_405347;
   reg _405348_405348 ; 
   reg __405348_405348;
   reg _405349_405349 ; 
   reg __405349_405349;
   reg _405350_405350 ; 
   reg __405350_405350;
   reg _405351_405351 ; 
   reg __405351_405351;
   reg _405352_405352 ; 
   reg __405352_405352;
   reg _405353_405353 ; 
   reg __405353_405353;
   reg _405354_405354 ; 
   reg __405354_405354;
   reg _405355_405355 ; 
   reg __405355_405355;
   reg _405356_405356 ; 
   reg __405356_405356;
   reg _405357_405357 ; 
   reg __405357_405357;
   reg _405358_405358 ; 
   reg __405358_405358;
   reg _405359_405359 ; 
   reg __405359_405359;
   reg _405360_405360 ; 
   reg __405360_405360;
   reg _405361_405361 ; 
   reg __405361_405361;
   reg _405362_405362 ; 
   reg __405362_405362;
   reg _405363_405363 ; 
   reg __405363_405363;
   reg _405364_405364 ; 
   reg __405364_405364;
   reg _405365_405365 ; 
   reg __405365_405365;
   reg _405366_405366 ; 
   reg __405366_405366;
   reg _405367_405367 ; 
   reg __405367_405367;
   reg _405368_405368 ; 
   reg __405368_405368;
   reg _405369_405369 ; 
   reg __405369_405369;
   reg _405370_405370 ; 
   reg __405370_405370;
   reg _405371_405371 ; 
   reg __405371_405371;
   reg _405372_405372 ; 
   reg __405372_405372;
   reg _405373_405373 ; 
   reg __405373_405373;
   reg _405374_405374 ; 
   reg __405374_405374;
   reg _405375_405375 ; 
   reg __405375_405375;
   reg _405376_405376 ; 
   reg __405376_405376;
   reg _405377_405377 ; 
   reg __405377_405377;
   reg _405378_405378 ; 
   reg __405378_405378;
   reg _405379_405379 ; 
   reg __405379_405379;
   reg _405380_405380 ; 
   reg __405380_405380;
   reg _405381_405381 ; 
   reg __405381_405381;
   reg _405382_405382 ; 
   reg __405382_405382;
   reg _405383_405383 ; 
   reg __405383_405383;
   reg _405384_405384 ; 
   reg __405384_405384;
   reg _405385_405385 ; 
   reg __405385_405385;
   reg _405386_405386 ; 
   reg __405386_405386;
   reg _405387_405387 ; 
   reg __405387_405387;
   reg _405388_405388 ; 
   reg __405388_405388;
   reg _405389_405389 ; 
   reg __405389_405389;
   reg _405390_405390 ; 
   reg __405390_405390;
   reg _405391_405391 ; 
   reg __405391_405391;
   reg _405392_405392 ; 
   reg __405392_405392;
   reg _405393_405393 ; 
   reg __405393_405393;
   reg _405394_405394 ; 
   reg __405394_405394;
   reg _405395_405395 ; 
   reg __405395_405395;
   reg _405396_405396 ; 
   reg __405396_405396;
   reg _405397_405397 ; 
   reg __405397_405397;
   reg _405398_405398 ; 
   reg __405398_405398;
   reg _405399_405399 ; 
   reg __405399_405399;
   reg _405400_405400 ; 
   reg __405400_405400;
   reg _405401_405401 ; 
   reg __405401_405401;
   reg _405402_405402 ; 
   reg __405402_405402;
   reg _405403_405403 ; 
   reg __405403_405403;
   reg _405404_405404 ; 
   reg __405404_405404;
   reg _405405_405405 ; 
   reg __405405_405405;
   reg _405406_405406 ; 
   reg __405406_405406;
   reg _405407_405407 ; 
   reg __405407_405407;
   reg _405408_405408 ; 
   reg __405408_405408;
   reg _405409_405409 ; 
   reg __405409_405409;
   reg _405410_405410 ; 
   reg __405410_405410;
   reg _405411_405411 ; 
   reg __405411_405411;
   reg _405412_405412 ; 
   reg __405412_405412;
   reg _405413_405413 ; 
   reg __405413_405413;
   reg _405414_405414 ; 
   reg __405414_405414;
   reg _405415_405415 ; 
   reg __405415_405415;
   reg _405416_405416 ; 
   reg __405416_405416;
   reg _405417_405417 ; 
   reg __405417_405417;
   reg _405418_405418 ; 
   reg __405418_405418;
   reg _405419_405419 ; 
   reg __405419_405419;
   reg _405420_405420 ; 
   reg __405420_405420;
   reg _405421_405421 ; 
   reg __405421_405421;
   reg _405422_405422 ; 
   reg __405422_405422;
   reg _405423_405423 ; 
   reg __405423_405423;
   reg _405424_405424 ; 
   reg __405424_405424;
   reg _405425_405425 ; 
   reg __405425_405425;
   reg _405426_405426 ; 
   reg __405426_405426;
   reg _405427_405427 ; 
   reg __405427_405427;
   reg _405428_405428 ; 
   reg __405428_405428;
   reg _405429_405429 ; 
   reg __405429_405429;
   reg _405430_405430 ; 
   reg __405430_405430;
   reg _405431_405431 ; 
   reg __405431_405431;
   reg _405432_405432 ; 
   reg __405432_405432;
   reg _405433_405433 ; 
   reg __405433_405433;
   reg _405434_405434 ; 
   reg __405434_405434;
   reg _405435_405435 ; 
   reg __405435_405435;
   reg _405436_405436 ; 
   reg __405436_405436;
   reg _405437_405437 ; 
   reg __405437_405437;
   reg _405438_405438 ; 
   reg __405438_405438;
   reg _405439_405439 ; 
   reg __405439_405439;
   reg _405440_405440 ; 
   reg __405440_405440;
   reg _405441_405441 ; 
   reg __405441_405441;
   reg _405442_405442 ; 
   reg __405442_405442;
   reg _405443_405443 ; 
   reg __405443_405443;
   reg _405444_405444 ; 
   reg __405444_405444;
   reg _405445_405445 ; 
   reg __405445_405445;
   reg _405446_405446 ; 
   reg __405446_405446;
   reg _405447_405447 ; 
   reg __405447_405447;
   reg _405448_405448 ; 
   reg __405448_405448;
   reg _405449_405449 ; 
   reg __405449_405449;
   reg _405450_405450 ; 
   reg __405450_405450;
   reg _405451_405451 ; 
   reg __405451_405451;
   reg _405452_405452 ; 
   reg __405452_405452;
   reg _405453_405453 ; 
   reg __405453_405453;
   reg _405454_405454 ; 
   reg __405454_405454;
   reg _405455_405455 ; 
   reg __405455_405455;
   reg _405456_405456 ; 
   reg __405456_405456;
   reg _405457_405457 ; 
   reg __405457_405457;
   reg _405458_405458 ; 
   reg __405458_405458;
   reg _405459_405459 ; 
   reg __405459_405459;
   reg _405460_405460 ; 
   reg __405460_405460;
   reg _405461_405461 ; 
   reg __405461_405461;
   reg _405462_405462 ; 
   reg __405462_405462;
   reg _405463_405463 ; 
   reg __405463_405463;
   reg _405464_405464 ; 
   reg __405464_405464;
   reg _405465_405465 ; 
   reg __405465_405465;
   reg _405466_405466 ; 
   reg __405466_405466;
   reg _405467_405467 ; 
   reg __405467_405467;
   reg _405468_405468 ; 
   reg __405468_405468;
   reg _405469_405469 ; 
   reg __405469_405469;
   reg _405470_405470 ; 
   reg __405470_405470;
   reg _405471_405471 ; 
   reg __405471_405471;
   reg _405472_405472 ; 
   reg __405472_405472;
   reg _405473_405473 ; 
   reg __405473_405473;
   reg _405474_405474 ; 
   reg __405474_405474;
   reg _405475_405475 ; 
   reg __405475_405475;
   reg _405476_405476 ; 
   reg __405476_405476;
   reg _405477_405477 ; 
   reg __405477_405477;
   reg _405478_405478 ; 
   reg __405478_405478;
   reg _405479_405479 ; 
   reg __405479_405479;
   reg _405480_405480 ; 
   reg __405480_405480;
   reg _405481_405481 ; 
   reg __405481_405481;
   reg _405482_405482 ; 
   reg __405482_405482;
   reg _405483_405483 ; 
   reg __405483_405483;
   reg _405484_405484 ; 
   reg __405484_405484;
   reg _405485_405485 ; 
   reg __405485_405485;
   reg _405486_405486 ; 
   reg __405486_405486;
   reg _405487_405487 ; 
   reg __405487_405487;
   reg _405488_405488 ; 
   reg __405488_405488;
   reg _405489_405489 ; 
   reg __405489_405489;
   reg _405490_405490 ; 
   reg __405490_405490;
   reg _405491_405491 ; 
   reg __405491_405491;
   reg _405492_405492 ; 
   reg __405492_405492;
   reg _405493_405493 ; 
   reg __405493_405493;
   reg _405494_405494 ; 
   reg __405494_405494;
   reg _405495_405495 ; 
   reg __405495_405495;
   reg _405496_405496 ; 
   reg __405496_405496;
   reg _405497_405497 ; 
   reg __405497_405497;
   reg _405498_405498 ; 
   reg __405498_405498;
   reg _405499_405499 ; 
   reg __405499_405499;
   reg _405500_405500 ; 
   reg __405500_405500;
   reg _405501_405501 ; 
   reg __405501_405501;
   reg _405502_405502 ; 
   reg __405502_405502;
   reg _405503_405503 ; 
   reg __405503_405503;
   reg _405504_405504 ; 
   reg __405504_405504;
   reg _405505_405505 ; 
   reg __405505_405505;
   reg _405506_405506 ; 
   reg __405506_405506;
   reg _405507_405507 ; 
   reg __405507_405507;
   reg _405508_405508 ; 
   reg __405508_405508;
   reg _405509_405509 ; 
   reg __405509_405509;
   reg _405510_405510 ; 
   reg __405510_405510;
   reg _405511_405511 ; 
   reg __405511_405511;
   reg _405512_405512 ; 
   reg __405512_405512;
   reg _405513_405513 ; 
   reg __405513_405513;
   reg _405514_405514 ; 
   reg __405514_405514;
   reg _405515_405515 ; 
   reg __405515_405515;
   reg _405516_405516 ; 
   reg __405516_405516;
   reg _405517_405517 ; 
   reg __405517_405517;
   reg _405518_405518 ; 
   reg __405518_405518;
   reg _405519_405519 ; 
   reg __405519_405519;
   reg _405520_405520 ; 
   reg __405520_405520;
   reg _405521_405521 ; 
   reg __405521_405521;
   reg _405522_405522 ; 
   reg __405522_405522;
   reg _405523_405523 ; 
   reg __405523_405523;
   reg _405524_405524 ; 
   reg __405524_405524;
   reg _405525_405525 ; 
   reg __405525_405525;
   reg _405526_405526 ; 
   reg __405526_405526;
   reg _405527_405527 ; 
   reg __405527_405527;
   reg _405528_405528 ; 
   reg __405528_405528;
   reg _405529_405529 ; 
   reg __405529_405529;
   reg _405530_405530 ; 
   reg __405530_405530;
   reg _405531_405531 ; 
   reg __405531_405531;
   reg _405532_405532 ; 
   reg __405532_405532;
   reg _405533_405533 ; 
   reg __405533_405533;
   reg _405534_405534 ; 
   reg __405534_405534;
   reg _405535_405535 ; 
   reg __405535_405535;
   reg _405536_405536 ; 
   reg __405536_405536;
   reg _405537_405537 ; 
   reg __405537_405537;
   reg _405538_405538 ; 
   reg __405538_405538;
   reg _405539_405539 ; 
   reg __405539_405539;
   reg _405540_405540 ; 
   reg __405540_405540;
   reg _405541_405541 ; 
   reg __405541_405541;
   reg _405542_405542 ; 
   reg __405542_405542;
   reg _405543_405543 ; 
   reg __405543_405543;
   reg _405544_405544 ; 
   reg __405544_405544;
   reg _405545_405545 ; 
   reg __405545_405545;
   reg _405546_405546 ; 
   reg __405546_405546;
   reg _405547_405547 ; 
   reg __405547_405547;
   reg _405548_405548 ; 
   reg __405548_405548;
   reg _405549_405549 ; 
   reg __405549_405549;
   reg _405550_405550 ; 
   reg __405550_405550;
   reg _405551_405551 ; 
   reg __405551_405551;
   reg _405552_405552 ; 
   reg __405552_405552;
   reg _405553_405553 ; 
   reg __405553_405553;
   reg _405554_405554 ; 
   reg __405554_405554;
   reg _405555_405555 ; 
   reg __405555_405555;
   reg _405556_405556 ; 
   reg __405556_405556;
   reg _405557_405557 ; 
   reg __405557_405557;
   reg _405558_405558 ; 
   reg __405558_405558;
   reg _405559_405559 ; 
   reg __405559_405559;
   reg _405560_405560 ; 
   reg __405560_405560;
   reg _405561_405561 ; 
   reg __405561_405561;
   reg _405562_405562 ; 
   reg __405562_405562;
   reg _405563_405563 ; 
   reg __405563_405563;
   reg _405564_405564 ; 
   reg __405564_405564;
   reg _405565_405565 ; 
   reg __405565_405565;
   reg _405566_405566 ; 
   reg __405566_405566;
   reg _405567_405567 ; 
   reg __405567_405567;
   reg _405568_405568 ; 
   reg __405568_405568;
   reg _405569_405569 ; 
   reg __405569_405569;
   reg _405570_405570 ; 
   reg __405570_405570;
   reg _405571_405571 ; 
   reg __405571_405571;
   reg _405572_405572 ; 
   reg __405572_405572;
   reg _405573_405573 ; 
   reg __405573_405573;
   reg _405574_405574 ; 
   reg __405574_405574;
   reg _405575_405575 ; 
   reg __405575_405575;
   reg _405576_405576 ; 
   reg __405576_405576;
   reg _405577_405577 ; 
   reg __405577_405577;
   reg _405578_405578 ; 
   reg __405578_405578;
   reg _405579_405579 ; 
   reg __405579_405579;
   reg _405580_405580 ; 
   reg __405580_405580;
   reg _405581_405581 ; 
   reg __405581_405581;
   reg _405582_405582 ; 
   reg __405582_405582;
   reg _405583_405583 ; 
   reg __405583_405583;
   reg _405584_405584 ; 
   reg __405584_405584;
   reg _405585_405585 ; 
   reg __405585_405585;
   reg _405586_405586 ; 
   reg __405586_405586;
   reg _405587_405587 ; 
   reg __405587_405587;
   reg _405588_405588 ; 
   reg __405588_405588;
   reg _405589_405589 ; 
   reg __405589_405589;
   reg _405590_405590 ; 
   reg __405590_405590;
   reg _405591_405591 ; 
   reg __405591_405591;
   reg _405592_405592 ; 
   reg __405592_405592;
   reg _405593_405593 ; 
   reg __405593_405593;
   reg _405594_405594 ; 
   reg __405594_405594;
   reg _405595_405595 ; 
   reg __405595_405595;
   reg _405596_405596 ; 
   reg __405596_405596;
   reg _405597_405597 ; 
   reg __405597_405597;
   reg _405598_405598 ; 
   reg __405598_405598;
   reg _405599_405599 ; 
   reg __405599_405599;
   reg _405600_405600 ; 
   reg __405600_405600;
   reg _405601_405601 ; 
   reg __405601_405601;
   reg _405602_405602 ; 
   reg __405602_405602;
   reg _405603_405603 ; 
   reg __405603_405603;
   reg _405604_405604 ; 
   reg __405604_405604;
   reg _405605_405605 ; 
   reg __405605_405605;
   reg _405606_405606 ; 
   reg __405606_405606;
   reg _405607_405607 ; 
   reg __405607_405607;
   reg _405608_405608 ; 
   reg __405608_405608;
   reg _405609_405609 ; 
   reg __405609_405609;
   reg _405610_405610 ; 
   reg __405610_405610;
   reg _405611_405611 ; 
   reg __405611_405611;
   reg _405612_405612 ; 
   reg __405612_405612;
   reg _405613_405613 ; 
   reg __405613_405613;
   reg _405614_405614 ; 
   reg __405614_405614;
   reg _405615_405615 ; 
   reg __405615_405615;
   reg _405616_405616 ; 
   reg __405616_405616;
   reg _405617_405617 ; 
   reg __405617_405617;
   reg _405618_405618 ; 
   reg __405618_405618;
   reg _405619_405619 ; 
   reg __405619_405619;
   reg _405620_405620 ; 
   reg __405620_405620;
   reg _405621_405621 ; 
   reg __405621_405621;
   reg _405622_405622 ; 
   reg __405622_405622;
   reg _405623_405623 ; 
   reg __405623_405623;
   reg _405624_405624 ; 
   reg __405624_405624;
   reg _405625_405625 ; 
   reg __405625_405625;
   reg _405626_405626 ; 
   reg __405626_405626;
   reg _405627_405627 ; 
   reg __405627_405627;
   reg _405628_405628 ; 
   reg __405628_405628;
   reg _405629_405629 ; 
   reg __405629_405629;
   reg _405630_405630 ; 
   reg __405630_405630;
   reg _405631_405631 ; 
   reg __405631_405631;
   reg _405632_405632 ; 
   reg __405632_405632;
   reg _405633_405633 ; 
   reg __405633_405633;
   reg _405634_405634 ; 
   reg __405634_405634;
   reg _405635_405635 ; 
   reg __405635_405635;
   reg _405636_405636 ; 
   reg __405636_405636;
   reg _405637_405637 ; 
   reg __405637_405637;
   reg _405638_405638 ; 
   reg __405638_405638;
   reg _405639_405639 ; 
   reg __405639_405639;
   reg _405640_405640 ; 
   reg __405640_405640;
   reg _405641_405641 ; 
   reg __405641_405641;
   reg _405642_405642 ; 
   reg __405642_405642;
   reg _405643_405643 ; 
   reg __405643_405643;
   reg _405644_405644 ; 
   reg __405644_405644;
   reg _405645_405645 ; 
   reg __405645_405645;
   reg _405646_405646 ; 
   reg __405646_405646;
   reg _405647_405647 ; 
   reg __405647_405647;
   reg _405648_405648 ; 
   reg __405648_405648;
   reg _405649_405649 ; 
   reg __405649_405649;
   reg _405650_405650 ; 
   reg __405650_405650;
   reg _405651_405651 ; 
   reg __405651_405651;
   reg _405652_405652 ; 
   reg __405652_405652;
   reg _405653_405653 ; 
   reg __405653_405653;
   reg _405654_405654 ; 
   reg __405654_405654;
   reg _405655_405655 ; 
   reg __405655_405655;
   reg _405656_405656 ; 
   reg __405656_405656;
   reg _405657_405657 ; 
   reg __405657_405657;
   reg _405658_405658 ; 
   reg __405658_405658;
   reg _405659_405659 ; 
   reg __405659_405659;
   reg _405660_405660 ; 
   reg __405660_405660;
   reg _405661_405661 ; 
   reg __405661_405661;
   reg _405662_405662 ; 
   reg __405662_405662;
   reg _405663_405663 ; 
   reg __405663_405663;
   reg _405664_405664 ; 
   reg __405664_405664;
   reg _405665_405665 ; 
   reg __405665_405665;
   reg _405666_405666 ; 
   reg __405666_405666;
   reg _405667_405667 ; 
   reg __405667_405667;
   reg _405668_405668 ; 
   reg __405668_405668;
   reg _405669_405669 ; 
   reg __405669_405669;
   reg _405670_405670 ; 
   reg __405670_405670;
   reg _405671_405671 ; 
   reg __405671_405671;
   reg _405672_405672 ; 
   reg __405672_405672;
   reg _405673_405673 ; 
   reg __405673_405673;
   reg _405674_405674 ; 
   reg __405674_405674;
   reg _405675_405675 ; 
   reg __405675_405675;
   reg _405676_405676 ; 
   reg __405676_405676;
   reg _405677_405677 ; 
   reg __405677_405677;
   reg _405678_405678 ; 
   reg __405678_405678;
   reg _405679_405679 ; 
   reg __405679_405679;
   reg _405680_405680 ; 
   reg __405680_405680;
   reg _405681_405681 ; 
   reg __405681_405681;
   reg _405682_405682 ; 
   reg __405682_405682;
   reg _405683_405683 ; 
   reg __405683_405683;
   reg _405684_405684 ; 
   reg __405684_405684;
   reg _405685_405685 ; 
   reg __405685_405685;
   reg _405686_405686 ; 
   reg __405686_405686;
   reg _405687_405687 ; 
   reg __405687_405687;
   reg _405688_405688 ; 
   reg __405688_405688;
   reg _405689_405689 ; 
   reg __405689_405689;
   reg _405690_405690 ; 
   reg __405690_405690;
   reg _405691_405691 ; 
   reg __405691_405691;
   reg _405692_405692 ; 
   reg __405692_405692;
   reg _405693_405693 ; 
   reg __405693_405693;
   reg _405694_405694 ; 
   reg __405694_405694;
   reg _405695_405695 ; 
   reg __405695_405695;
   reg _405696_405696 ; 
   reg __405696_405696;
   reg _405697_405697 ; 
   reg __405697_405697;
   reg _405698_405698 ; 
   reg __405698_405698;
   reg _405699_405699 ; 
   reg __405699_405699;
   reg _405700_405700 ; 
   reg __405700_405700;
   reg _405701_405701 ; 
   reg __405701_405701;
   reg _405702_405702 ; 
   reg __405702_405702;
   reg _405703_405703 ; 
   reg __405703_405703;
   reg _405704_405704 ; 
   reg __405704_405704;
   reg _405705_405705 ; 
   reg __405705_405705;
   reg _405706_405706 ; 
   reg __405706_405706;
   reg _405707_405707 ; 
   reg __405707_405707;
   reg _405708_405708 ; 
   reg __405708_405708;
   reg _405709_405709 ; 
   reg __405709_405709;
   reg _405710_405710 ; 
   reg __405710_405710;
   reg _405711_405711 ; 
   reg __405711_405711;
   reg _405712_405712 ; 
   reg __405712_405712;
   reg _405713_405713 ; 
   reg __405713_405713;
   reg _405714_405714 ; 
   reg __405714_405714;
   reg _405715_405715 ; 
   reg __405715_405715;
   reg _405716_405716 ; 
   reg __405716_405716;
   reg _405717_405717 ; 
   reg __405717_405717;
   reg _405718_405718 ; 
   reg __405718_405718;
   reg _405719_405719 ; 
   reg __405719_405719;
   reg _405720_405720 ; 
   reg __405720_405720;
   reg _405721_405721 ; 
   reg __405721_405721;
   reg _405722_405722 ; 
   reg __405722_405722;
   reg _405723_405723 ; 
   reg __405723_405723;
   reg _405724_405724 ; 
   reg __405724_405724;
   reg _405725_405725 ; 
   reg __405725_405725;
   reg _405726_405726 ; 
   reg __405726_405726;
   reg _405727_405727 ; 
   reg __405727_405727;
   reg _405728_405728 ; 
   reg __405728_405728;
   reg _405729_405729 ; 
   reg __405729_405729;
   reg _405730_405730 ; 
   reg __405730_405730;
   reg _405731_405731 ; 
   reg __405731_405731;
   reg _405732_405732 ; 
   reg __405732_405732;
   reg _405733_405733 ; 
   reg __405733_405733;
   reg _405734_405734 ; 
   reg __405734_405734;
   reg _405735_405735 ; 
   reg __405735_405735;
   reg _405736_405736 ; 
   reg __405736_405736;
   reg _405737_405737 ; 
   reg __405737_405737;
   reg _405738_405738 ; 
   reg __405738_405738;
   reg _405739_405739 ; 
   reg __405739_405739;
   reg _405740_405740 ; 
   reg __405740_405740;
   reg _405741_405741 ; 
   reg __405741_405741;
   reg _405742_405742 ; 
   reg __405742_405742;
   reg _405743_405743 ; 
   reg __405743_405743;
   reg _405744_405744 ; 
   reg __405744_405744;
   reg _405745_405745 ; 
   reg __405745_405745;
   reg _405746_405746 ; 
   reg __405746_405746;
   reg _405747_405747 ; 
   reg __405747_405747;
   reg _405748_405748 ; 
   reg __405748_405748;
   reg _405749_405749 ; 
   reg __405749_405749;
   reg _405750_405750 ; 
   reg __405750_405750;
   reg _405751_405751 ; 
   reg __405751_405751;
   reg _405752_405752 ; 
   reg __405752_405752;
   reg _405753_405753 ; 
   reg __405753_405753;
   reg _405754_405754 ; 
   reg __405754_405754;
   reg _405755_405755 ; 
   reg __405755_405755;
   reg _405756_405756 ; 
   reg __405756_405756;
   reg _405757_405757 ; 
   reg __405757_405757;
   reg _405758_405758 ; 
   reg __405758_405758;
   reg _405759_405759 ; 
   reg __405759_405759;
   reg _405760_405760 ; 
   reg __405760_405760;
   reg _405761_405761 ; 
   reg __405761_405761;
   reg _405762_405762 ; 
   reg __405762_405762;
   reg _405763_405763 ; 
   reg __405763_405763;
   reg _405764_405764 ; 
   reg __405764_405764;
   reg _405765_405765 ; 
   reg __405765_405765;
   reg _405766_405766 ; 
   reg __405766_405766;
   reg _405767_405767 ; 
   reg __405767_405767;
   reg _405768_405768 ; 
   reg __405768_405768;
   reg _405769_405769 ; 
   reg __405769_405769;
   reg _405770_405770 ; 
   reg __405770_405770;
   reg _405771_405771 ; 
   reg __405771_405771;
   reg _405772_405772 ; 
   reg __405772_405772;
   reg _405773_405773 ; 
   reg __405773_405773;
   reg _405774_405774 ; 
   reg __405774_405774;
   reg _405775_405775 ; 
   reg __405775_405775;
   reg _405776_405776 ; 
   reg __405776_405776;
   reg _405777_405777 ; 
   reg __405777_405777;
   reg _405778_405778 ; 
   reg __405778_405778;
   reg _405779_405779 ; 
   reg __405779_405779;
   reg _405780_405780 ; 
   reg __405780_405780;
   reg _405781_405781 ; 
   reg __405781_405781;
   reg _405782_405782 ; 
   reg __405782_405782;
   reg _405783_405783 ; 
   reg __405783_405783;
   reg _405784_405784 ; 
   reg __405784_405784;
   reg _405785_405785 ; 
   reg __405785_405785;
   reg _405786_405786 ; 
   reg __405786_405786;
   reg _405787_405787 ; 
   reg __405787_405787;
   reg _405788_405788 ; 
   reg __405788_405788;
   reg _405789_405789 ; 
   reg __405789_405789;
   reg _405790_405790 ; 
   reg __405790_405790;
   reg _405791_405791 ; 
   reg __405791_405791;
   reg _405792_405792 ; 
   reg __405792_405792;
   reg _405793_405793 ; 
   reg __405793_405793;
   reg _405794_405794 ; 
   reg __405794_405794;
   reg _405795_405795 ; 
   reg __405795_405795;
   reg _405796_405796 ; 
   reg __405796_405796;
   reg _405797_405797 ; 
   reg __405797_405797;
   reg _405798_405798 ; 
   reg __405798_405798;
   reg _405799_405799 ; 
   reg __405799_405799;
   reg _405800_405800 ; 
   reg __405800_405800;
   reg _405801_405801 ; 
   reg __405801_405801;
   reg _405802_405802 ; 
   reg __405802_405802;
   reg _405803_405803 ; 
   reg __405803_405803;
   reg _405804_405804 ; 
   reg __405804_405804;
   reg _405805_405805 ; 
   reg __405805_405805;
   reg _405806_405806 ; 
   reg __405806_405806;
   reg _405807_405807 ; 
   reg __405807_405807;
   reg _405808_405808 ; 
   reg __405808_405808;
   reg _405809_405809 ; 
   reg __405809_405809;
   reg _405810_405810 ; 
   reg __405810_405810;
   reg _405811_405811 ; 
   reg __405811_405811;
   reg _405812_405812 ; 
   reg __405812_405812;
   reg _405813_405813 ; 
   reg __405813_405813;
   reg _405814_405814 ; 
   reg __405814_405814;
   reg _405815_405815 ; 
   reg __405815_405815;
   reg _405816_405816 ; 
   reg __405816_405816;
   reg _405817_405817 ; 
   reg __405817_405817;
   reg _405818_405818 ; 
   reg __405818_405818;
   reg _405819_405819 ; 
   reg __405819_405819;
   reg _405820_405820 ; 
   reg __405820_405820;
   reg _405821_405821 ; 
   reg __405821_405821;
   reg _405822_405822 ; 
   reg __405822_405822;
   reg _405823_405823 ; 
   reg __405823_405823;
   reg _405824_405824 ; 
   reg __405824_405824;
   reg _405825_405825 ; 
   reg __405825_405825;
   reg _405826_405826 ; 
   reg __405826_405826;
   reg _405827_405827 ; 
   reg __405827_405827;
   reg _405828_405828 ; 
   reg __405828_405828;
   reg _405829_405829 ; 
   reg __405829_405829;
   reg _405830_405830 ; 
   reg __405830_405830;
   reg _405831_405831 ; 
   reg __405831_405831;
   reg _405832_405832 ; 
   reg __405832_405832;
   reg _405833_405833 ; 
   reg __405833_405833;
   reg _405834_405834 ; 
   reg __405834_405834;
   reg _405835_405835 ; 
   reg __405835_405835;
   reg _405836_405836 ; 
   reg __405836_405836;
   reg _405837_405837 ; 
   reg __405837_405837;
   reg _405838_405838 ; 
   reg __405838_405838;
   reg _405839_405839 ; 
   reg __405839_405839;
   reg _405840_405840 ; 
   reg __405840_405840;
   reg _405841_405841 ; 
   reg __405841_405841;
   reg _405842_405842 ; 
   reg __405842_405842;
   reg _405843_405843 ; 
   reg __405843_405843;
   reg _405844_405844 ; 
   reg __405844_405844;
   reg _405845_405845 ; 
   reg __405845_405845;
   reg _405846_405846 ; 
   reg __405846_405846;
   reg _405847_405847 ; 
   reg __405847_405847;
   reg _405848_405848 ; 
   reg __405848_405848;
   reg _405849_405849 ; 
   reg __405849_405849;
   reg _405850_405850 ; 
   reg __405850_405850;
   reg _405851_405851 ; 
   reg __405851_405851;
   reg _405852_405852 ; 
   reg __405852_405852;
   reg _405853_405853 ; 
   reg __405853_405853;
   reg _405854_405854 ; 
   reg __405854_405854;
   reg _405855_405855 ; 
   reg __405855_405855;
   reg _405856_405856 ; 
   reg __405856_405856;
   reg _405857_405857 ; 
   reg __405857_405857;
   reg _405858_405858 ; 
   reg __405858_405858;
   reg _405859_405859 ; 
   reg __405859_405859;
   reg _405860_405860 ; 
   reg __405860_405860;
   reg _405861_405861 ; 
   reg __405861_405861;
   reg _405862_405862 ; 
   reg __405862_405862;
   reg _405863_405863 ; 
   reg __405863_405863;
   reg _405864_405864 ; 
   reg __405864_405864;
   reg _405865_405865 ; 
   reg __405865_405865;
   reg _405866_405866 ; 
   reg __405866_405866;
   reg _405867_405867 ; 
   reg __405867_405867;
   reg _405868_405868 ; 
   reg __405868_405868;
   reg _405869_405869 ; 
   reg __405869_405869;
   reg _405870_405870 ; 
   reg __405870_405870;
   reg _405871_405871 ; 
   reg __405871_405871;
   reg _405872_405872 ; 
   reg __405872_405872;
   reg _405873_405873 ; 
   reg __405873_405873;
   reg _405874_405874 ; 
   reg __405874_405874;
   reg _405875_405875 ; 
   reg __405875_405875;
   reg _405876_405876 ; 
   reg __405876_405876;
   reg _405877_405877 ; 
   reg __405877_405877;
   reg _405878_405878 ; 
   reg __405878_405878;
   reg _405879_405879 ; 
   reg __405879_405879;
   reg _405880_405880 ; 
   reg __405880_405880;
   reg _405881_405881 ; 
   reg __405881_405881;
   reg _405882_405882 ; 
   reg __405882_405882;
   reg _405883_405883 ; 
   reg __405883_405883;
   reg _405884_405884 ; 
   reg __405884_405884;
   reg _405885_405885 ; 
   reg __405885_405885;
   reg _405886_405886 ; 
   reg __405886_405886;
   reg _405887_405887 ; 
   reg __405887_405887;
   reg _405888_405888 ; 
   reg __405888_405888;
   reg _405889_405889 ; 
   reg __405889_405889;
   reg _405890_405890 ; 
   reg __405890_405890;
   reg _405891_405891 ; 
   reg __405891_405891;
   reg _405892_405892 ; 
   reg __405892_405892;
   reg _405893_405893 ; 
   reg __405893_405893;
   reg _405894_405894 ; 
   reg __405894_405894;
   reg _405895_405895 ; 
   reg __405895_405895;
   reg _405896_405896 ; 
   reg __405896_405896;
   reg _405897_405897 ; 
   reg __405897_405897;
   reg _405898_405898 ; 
   reg __405898_405898;
   reg _405899_405899 ; 
   reg __405899_405899;
   reg _405900_405900 ; 
   reg __405900_405900;
   reg _405901_405901 ; 
   reg __405901_405901;
   reg _405902_405902 ; 
   reg __405902_405902;
   reg _405903_405903 ; 
   reg __405903_405903;
   reg _405904_405904 ; 
   reg __405904_405904;
   reg _405905_405905 ; 
   reg __405905_405905;
   reg _405906_405906 ; 
   reg __405906_405906;
   reg _405907_405907 ; 
   reg __405907_405907;
   reg _405908_405908 ; 
   reg __405908_405908;
   reg _405909_405909 ; 
   reg __405909_405909;
   reg _405910_405910 ; 
   reg __405910_405910;
   reg _405911_405911 ; 
   reg __405911_405911;
   reg _405912_405912 ; 
   reg __405912_405912;
   reg _405913_405913 ; 
   reg __405913_405913;
   reg _405914_405914 ; 
   reg __405914_405914;
   reg _405915_405915 ; 
   reg __405915_405915;
   reg _405916_405916 ; 
   reg __405916_405916;
   reg _405917_405917 ; 
   reg __405917_405917;
   reg _405918_405918 ; 
   reg __405918_405918;
   reg _405919_405919 ; 
   reg __405919_405919;
   reg _405920_405920 ; 
   reg __405920_405920;
   reg _405921_405921 ; 
   reg __405921_405921;
   reg _405922_405922 ; 
   reg __405922_405922;
   reg _405923_405923 ; 
   reg __405923_405923;
   reg _405924_405924 ; 
   reg __405924_405924;
   reg _405925_405925 ; 
   reg __405925_405925;
   reg _405926_405926 ; 
   reg __405926_405926;
   reg _405927_405927 ; 
   reg __405927_405927;
   reg _405928_405928 ; 
   reg __405928_405928;
   reg _405929_405929 ; 
   reg __405929_405929;
   reg _405930_405930 ; 
   reg __405930_405930;
   reg _405931_405931 ; 
   reg __405931_405931;
   reg _405932_405932 ; 
   reg __405932_405932;
   reg _405933_405933 ; 
   reg __405933_405933;
   reg _405934_405934 ; 
   reg __405934_405934;
   reg _405935_405935 ; 
   reg __405935_405935;
   reg _405936_405936 ; 
   reg __405936_405936;
   reg _405937_405937 ; 
   reg __405937_405937;
   reg _405938_405938 ; 
   reg __405938_405938;
   reg _405939_405939 ; 
   reg __405939_405939;
   reg _405940_405940 ; 
   reg __405940_405940;
   reg _405941_405941 ; 
   reg __405941_405941;
   reg _405942_405942 ; 
   reg __405942_405942;
   reg _405943_405943 ; 
   reg __405943_405943;
   reg _405944_405944 ; 
   reg __405944_405944;
   reg _405945_405945 ; 
   reg __405945_405945;
   reg _405946_405946 ; 
   reg __405946_405946;
   reg _405947_405947 ; 
   reg __405947_405947;
   reg _405948_405948 ; 
   reg __405948_405948;
   reg _405949_405949 ; 
   reg __405949_405949;
   reg _405950_405950 ; 
   reg __405950_405950;
   reg _405951_405951 ; 
   reg __405951_405951;
   reg _405952_405952 ; 
   reg __405952_405952;
   reg _405953_405953 ; 
   reg __405953_405953;
   reg _405954_405954 ; 
   reg __405954_405954;
   reg _405955_405955 ; 
   reg __405955_405955;
   reg _405956_405956 ; 
   reg __405956_405956;
   reg _405957_405957 ; 
   reg __405957_405957;
   reg _405958_405958 ; 
   reg __405958_405958;
   reg _405959_405959 ; 
   reg __405959_405959;
   reg _405960_405960 ; 
   reg __405960_405960;
   reg _405961_405961 ; 
   reg __405961_405961;
   reg _405962_405962 ; 
   reg __405962_405962;
   reg _405963_405963 ; 
   reg __405963_405963;
   reg _405964_405964 ; 
   reg __405964_405964;
   reg _405965_405965 ; 
   reg __405965_405965;
   reg _405966_405966 ; 
   reg __405966_405966;
   reg _405967_405967 ; 
   reg __405967_405967;
   reg _405968_405968 ; 
   reg __405968_405968;
   reg _405969_405969 ; 
   reg __405969_405969;
   reg _405970_405970 ; 
   reg __405970_405970;
   reg _405971_405971 ; 
   reg __405971_405971;
   reg _405972_405972 ; 
   reg __405972_405972;
   reg _405973_405973 ; 
   reg __405973_405973;
   reg _405974_405974 ; 
   reg __405974_405974;
   reg _405975_405975 ; 
   reg __405975_405975;
   reg _405976_405976 ; 
   reg __405976_405976;
   reg _405977_405977 ; 
   reg __405977_405977;
   reg _405978_405978 ; 
   reg __405978_405978;
   reg _405979_405979 ; 
   reg __405979_405979;
   reg _405980_405980 ; 
   reg __405980_405980;
   reg _405981_405981 ; 
   reg __405981_405981;
   reg _405982_405982 ; 
   reg __405982_405982;
   reg _405983_405983 ; 
   reg __405983_405983;
   reg _405984_405984 ; 
   reg __405984_405984;
   reg _405985_405985 ; 
   reg __405985_405985;
   reg _405986_405986 ; 
   reg __405986_405986;
   reg _405987_405987 ; 
   reg __405987_405987;
   reg _405988_405988 ; 
   reg __405988_405988;
   reg _405989_405989 ; 
   reg __405989_405989;
   reg _405990_405990 ; 
   reg __405990_405990;
   reg _405991_405991 ; 
   reg __405991_405991;
   reg _405992_405992 ; 
   reg __405992_405992;
   reg _405993_405993 ; 
   reg __405993_405993;
   reg _405994_405994 ; 
   reg __405994_405994;
   reg _405995_405995 ; 
   reg __405995_405995;
   reg _405996_405996 ; 
   reg __405996_405996;
   reg _405997_405997 ; 
   reg __405997_405997;
   reg _405998_405998 ; 
   reg __405998_405998;
   reg _405999_405999 ; 
   reg __405999_405999;
   reg _406000_406000 ; 
   reg __406000_406000;
   reg _406001_406001 ; 
   reg __406001_406001;
   reg _406002_406002 ; 
   reg __406002_406002;
   reg _406003_406003 ; 
   reg __406003_406003;
   reg _406004_406004 ; 
   reg __406004_406004;
   reg _406005_406005 ; 
   reg __406005_406005;
   reg _406006_406006 ; 
   reg __406006_406006;
   reg _406007_406007 ; 
   reg __406007_406007;
   reg _406008_406008 ; 
   reg __406008_406008;
   reg _406009_406009 ; 
   reg __406009_406009;
   reg _406010_406010 ; 
   reg __406010_406010;
   reg _406011_406011 ; 
   reg __406011_406011;
   reg _406012_406012 ; 
   reg __406012_406012;
   reg _406013_406013 ; 
   reg __406013_406013;
   reg _406014_406014 ; 
   reg __406014_406014;
   reg _406015_406015 ; 
   reg __406015_406015;
   reg _406016_406016 ; 
   reg __406016_406016;
   reg _406017_406017 ; 
   reg __406017_406017;
   reg _406018_406018 ; 
   reg __406018_406018;
   reg _406019_406019 ; 
   reg __406019_406019;
   reg _406020_406020 ; 
   reg __406020_406020;
   reg _406021_406021 ; 
   reg __406021_406021;
   reg _406022_406022 ; 
   reg __406022_406022;
   reg _406023_406023 ; 
   reg __406023_406023;
   reg _406024_406024 ; 
   reg __406024_406024;
   reg _406025_406025 ; 
   reg __406025_406025;
   reg _406026_406026 ; 
   reg __406026_406026;
   reg _406027_406027 ; 
   reg __406027_406027;
   reg _406028_406028 ; 
   reg __406028_406028;
   reg _406029_406029 ; 
   reg __406029_406029;
   reg _406030_406030 ; 
   reg __406030_406030;
   reg _406031_406031 ; 
   reg __406031_406031;
   reg _406032_406032 ; 
   reg __406032_406032;
   reg _406033_406033 ; 
   reg __406033_406033;
   reg _406034_406034 ; 
   reg __406034_406034;
   reg _406035_406035 ; 
   reg __406035_406035;
   reg _406036_406036 ; 
   reg __406036_406036;
   reg _406037_406037 ; 
   reg __406037_406037;
   reg _406038_406038 ; 
   reg __406038_406038;
   reg _406039_406039 ; 
   reg __406039_406039;
   reg _406040_406040 ; 
   reg __406040_406040;
   reg _406041_406041 ; 
   reg __406041_406041;
   reg _406042_406042 ; 
   reg __406042_406042;
   reg _406043_406043 ; 
   reg __406043_406043;
   reg _406044_406044 ; 
   reg __406044_406044;
   reg _406045_406045 ; 
   reg __406045_406045;
   reg _406046_406046 ; 
   reg __406046_406046;
   reg _406047_406047 ; 
   reg __406047_406047;
   reg _406048_406048 ; 
   reg __406048_406048;
   reg _406049_406049 ; 
   reg __406049_406049;
   reg _406050_406050 ; 
   reg __406050_406050;
   reg _406051_406051 ; 
   reg __406051_406051;
   reg _406052_406052 ; 
   reg __406052_406052;
   reg _406053_406053 ; 
   reg __406053_406053;
   reg _406054_406054 ; 
   reg __406054_406054;
   reg _406055_406055 ; 
   reg __406055_406055;
   reg _406056_406056 ; 
   reg __406056_406056;
   reg _406057_406057 ; 
   reg __406057_406057;
   reg _406058_406058 ; 
   reg __406058_406058;
   reg _406059_406059 ; 
   reg __406059_406059;
   reg _406060_406060 ; 
   reg __406060_406060;
   reg _406061_406061 ; 
   reg __406061_406061;
   reg _406062_406062 ; 
   reg __406062_406062;
   reg _406063_406063 ; 
   reg __406063_406063;
   reg _406064_406064 ; 
   reg __406064_406064;
   reg _406065_406065 ; 
   reg __406065_406065;
   reg _406066_406066 ; 
   reg __406066_406066;
   reg _406067_406067 ; 
   reg __406067_406067;
   reg _406068_406068 ; 
   reg __406068_406068;
   reg _406069_406069 ; 
   reg __406069_406069;
   reg _406070_406070 ; 
   reg __406070_406070;
   reg _406071_406071 ; 
   reg __406071_406071;
   reg _406072_406072 ; 
   reg __406072_406072;
   reg _406073_406073 ; 
   reg __406073_406073;
   reg _406074_406074 ; 
   reg __406074_406074;
   reg _406075_406075 ; 
   reg __406075_406075;
   reg _406076_406076 ; 
   reg __406076_406076;
   reg _406077_406077 ; 
   reg __406077_406077;
   reg _406078_406078 ; 
   reg __406078_406078;
   reg _406079_406079 ; 
   reg __406079_406079;
   reg _406080_406080 ; 
   reg __406080_406080;
   reg _406081_406081 ; 
   reg __406081_406081;
   reg _406082_406082 ; 
   reg __406082_406082;
   reg _406083_406083 ; 
   reg __406083_406083;
   reg _406084_406084 ; 
   reg __406084_406084;
   reg _406085_406085 ; 
   reg __406085_406085;
   reg _406086_406086 ; 
   reg __406086_406086;
   reg _406087_406087 ; 
   reg __406087_406087;
   reg _406088_406088 ; 
   reg __406088_406088;
   reg _406089_406089 ; 
   reg __406089_406089;
   reg _406090_406090 ; 
   reg __406090_406090;
   reg _406091_406091 ; 
   reg __406091_406091;
   reg _406092_406092 ; 
   reg __406092_406092;
   reg _406093_406093 ; 
   reg __406093_406093;
   reg _406094_406094 ; 
   reg __406094_406094;
   reg _406095_406095 ; 
   reg __406095_406095;
   reg _406096_406096 ; 
   reg __406096_406096;
   reg _406097_406097 ; 
   reg __406097_406097;
   reg _406098_406098 ; 
   reg __406098_406098;
   reg _406099_406099 ; 
   reg __406099_406099;
   reg _406100_406100 ; 
   reg __406100_406100;
   reg _406101_406101 ; 
   reg __406101_406101;
   reg _406102_406102 ; 
   reg __406102_406102;
   reg _406103_406103 ; 
   reg __406103_406103;
   reg _406104_406104 ; 
   reg __406104_406104;
   reg _406105_406105 ; 
   reg __406105_406105;
   reg _406106_406106 ; 
   reg __406106_406106;
   reg _406107_406107 ; 
   reg __406107_406107;
   reg _406108_406108 ; 
   reg __406108_406108;
   reg _406109_406109 ; 
   reg __406109_406109;
   reg _406110_406110 ; 
   reg __406110_406110;
   reg _406111_406111 ; 
   reg __406111_406111;
   reg _406112_406112 ; 
   reg __406112_406112;
   reg _406113_406113 ; 
   reg __406113_406113;
   reg _406114_406114 ; 
   reg __406114_406114;
   reg _406115_406115 ; 
   reg __406115_406115;
   reg _406116_406116 ; 
   reg __406116_406116;
   reg _406117_406117 ; 
   reg __406117_406117;
   reg _406118_406118 ; 
   reg __406118_406118;
   reg _406119_406119 ; 
   reg __406119_406119;
   reg _406120_406120 ; 
   reg __406120_406120;
   reg _406121_406121 ; 
   reg __406121_406121;
   reg _406122_406122 ; 
   reg __406122_406122;
   reg _406123_406123 ; 
   reg __406123_406123;
   reg _406124_406124 ; 
   reg __406124_406124;
   reg _406125_406125 ; 
   reg __406125_406125;
   reg _406126_406126 ; 
   reg __406126_406126;
   reg _406127_406127 ; 
   reg __406127_406127;
   reg _406128_406128 ; 
   reg __406128_406128;
   reg _406129_406129 ; 
   reg __406129_406129;
   reg _406130_406130 ; 
   reg __406130_406130;
   reg _406131_406131 ; 
   reg __406131_406131;
   reg _406132_406132 ; 
   reg __406132_406132;
   reg _406133_406133 ; 
   reg __406133_406133;
   reg _406134_406134 ; 
   reg __406134_406134;
   reg _406135_406135 ; 
   reg __406135_406135;
   reg _406136_406136 ; 
   reg __406136_406136;
   reg _406137_406137 ; 
   reg __406137_406137;
   reg _406138_406138 ; 
   reg __406138_406138;
   reg _406139_406139 ; 
   reg __406139_406139;
   reg _406140_406140 ; 
   reg __406140_406140;
   reg _406141_406141 ; 
   reg __406141_406141;
   reg _406142_406142 ; 
   reg __406142_406142;
   reg _406143_406143 ; 
   reg __406143_406143;
   reg _406144_406144 ; 
   reg __406144_406144;
   reg _406145_406145 ; 
   reg __406145_406145;
   reg _406146_406146 ; 
   reg __406146_406146;
   reg _406147_406147 ; 
   reg __406147_406147;
   reg _406148_406148 ; 
   reg __406148_406148;
   reg _406149_406149 ; 
   reg __406149_406149;
   reg _406150_406150 ; 
   reg __406150_406150;
   reg _406151_406151 ; 
   reg __406151_406151;
   reg _406152_406152 ; 
   reg __406152_406152;
   reg _406153_406153 ; 
   reg __406153_406153;
   reg _406154_406154 ; 
   reg __406154_406154;
   reg _406155_406155 ; 
   reg __406155_406155;
   reg _406156_406156 ; 
   reg __406156_406156;
   reg _406157_406157 ; 
   reg __406157_406157;
   reg _406158_406158 ; 
   reg __406158_406158;
   reg _406159_406159 ; 
   reg __406159_406159;
   reg _406160_406160 ; 
   reg __406160_406160;
   reg _406161_406161 ; 
   reg __406161_406161;
   reg _406162_406162 ; 
   reg __406162_406162;
   reg _406163_406163 ; 
   reg __406163_406163;
   reg _406164_406164 ; 
   reg __406164_406164;
   reg _406165_406165 ; 
   reg __406165_406165;
   reg _406166_406166 ; 
   reg __406166_406166;
   reg _406167_406167 ; 
   reg __406167_406167;
   reg _406168_406168 ; 
   reg __406168_406168;
   reg _406169_406169 ; 
   reg __406169_406169;
   reg _406170_406170 ; 
   reg __406170_406170;
   reg _406171_406171 ; 
   reg __406171_406171;
   reg _406172_406172 ; 
   reg __406172_406172;
   reg _406173_406173 ; 
   reg __406173_406173;
   reg _406174_406174 ; 
   reg __406174_406174;
   reg _406175_406175 ; 
   reg __406175_406175;
   reg _406176_406176 ; 
   reg __406176_406176;
   reg _406177_406177 ; 
   reg __406177_406177;
   reg _406178_406178 ; 
   reg __406178_406178;
   reg _406179_406179 ; 
   reg __406179_406179;
   reg _406180_406180 ; 
   reg __406180_406180;
   reg _406181_406181 ; 
   reg __406181_406181;
   reg _406182_406182 ; 
   reg __406182_406182;
   reg _406183_406183 ; 
   reg __406183_406183;
   reg _406184_406184 ; 
   reg __406184_406184;
   reg _406185_406185 ; 
   reg __406185_406185;
   reg _406186_406186 ; 
   reg __406186_406186;
   reg _406187_406187 ; 
   reg __406187_406187;
   reg _406188_406188 ; 
   reg __406188_406188;
   reg _406189_406189 ; 
   reg __406189_406189;
   reg _406190_406190 ; 
   reg __406190_406190;
   reg _406191_406191 ; 
   reg __406191_406191;
   reg _406192_406192 ; 
   reg __406192_406192;
   reg _406193_406193 ; 
   reg __406193_406193;
   reg _406194_406194 ; 
   reg __406194_406194;
   reg _406195_406195 ; 
   reg __406195_406195;
   reg _406196_406196 ; 
   reg __406196_406196;
   reg _406197_406197 ; 
   reg __406197_406197;
   reg _406198_406198 ; 
   reg __406198_406198;
   reg _406199_406199 ; 
   reg __406199_406199;
   reg _406200_406200 ; 
   reg __406200_406200;
   reg _406201_406201 ; 
   reg __406201_406201;
   reg _406202_406202 ; 
   reg __406202_406202;
   reg _406203_406203 ; 
   reg __406203_406203;
   reg _406204_406204 ; 
   reg __406204_406204;
   reg _406205_406205 ; 
   reg __406205_406205;
   reg _406206_406206 ; 
   reg __406206_406206;
   reg _406207_406207 ; 
   reg __406207_406207;
   reg _406208_406208 ; 
   reg __406208_406208;
   reg _406209_406209 ; 
   reg __406209_406209;
   reg _406210_406210 ; 
   reg __406210_406210;
   reg _406211_406211 ; 
   reg __406211_406211;
   reg _406212_406212 ; 
   reg __406212_406212;
   reg _406213_406213 ; 
   reg __406213_406213;
   reg _406214_406214 ; 
   reg __406214_406214;
   reg _406215_406215 ; 
   reg __406215_406215;
   reg _406216_406216 ; 
   reg __406216_406216;
   reg _406217_406217 ; 
   reg __406217_406217;
   reg _406218_406218 ; 
   reg __406218_406218;
   reg _406219_406219 ; 
   reg __406219_406219;
   reg _406220_406220 ; 
   reg __406220_406220;
   reg _406221_406221 ; 
   reg __406221_406221;
   reg _406222_406222 ; 
   reg __406222_406222;
   reg _406223_406223 ; 
   reg __406223_406223;
   reg _406224_406224 ; 
   reg __406224_406224;
   reg _406225_406225 ; 
   reg __406225_406225;
   reg _406226_406226 ; 
   reg __406226_406226;
   reg _406227_406227 ; 
   reg __406227_406227;
   reg _406228_406228 ; 
   reg __406228_406228;
   reg _406229_406229 ; 
   reg __406229_406229;
   reg _406230_406230 ; 
   reg __406230_406230;
   reg _406231_406231 ; 
   reg __406231_406231;
   reg _406232_406232 ; 
   reg __406232_406232;
   reg _406233_406233 ; 
   reg __406233_406233;
   reg _406234_406234 ; 
   reg __406234_406234;
   reg _406235_406235 ; 
   reg __406235_406235;
   reg _406236_406236 ; 
   reg __406236_406236;
   reg _406237_406237 ; 
   reg __406237_406237;
   reg _406238_406238 ; 
   reg __406238_406238;
   reg _406239_406239 ; 
   reg __406239_406239;
   reg _406240_406240 ; 
   reg __406240_406240;
   reg _406241_406241 ; 
   reg __406241_406241;
   reg _406242_406242 ; 
   reg __406242_406242;
   reg _406243_406243 ; 
   reg __406243_406243;
   reg _406244_406244 ; 
   reg __406244_406244;
   reg _406245_406245 ; 
   reg __406245_406245;
   reg _406246_406246 ; 
   reg __406246_406246;
   reg _406247_406247 ; 
   reg __406247_406247;
   reg _406248_406248 ; 
   reg __406248_406248;
   reg _406249_406249 ; 
   reg __406249_406249;
   reg _406250_406250 ; 
   reg __406250_406250;
   reg _406251_406251 ; 
   reg __406251_406251;
   reg _406252_406252 ; 
   reg __406252_406252;
   reg _406253_406253 ; 
   reg __406253_406253;
   reg _406254_406254 ; 
   reg __406254_406254;
   reg _406255_406255 ; 
   reg __406255_406255;
   reg _406256_406256 ; 
   reg __406256_406256;
   reg _406257_406257 ; 
   reg __406257_406257;
   reg _406258_406258 ; 
   reg __406258_406258;
   reg _406259_406259 ; 
   reg __406259_406259;
   reg _406260_406260 ; 
   reg __406260_406260;
   reg _406261_406261 ; 
   reg __406261_406261;
   reg _406262_406262 ; 
   reg __406262_406262;
   reg _406263_406263 ; 
   reg __406263_406263;
   reg _406264_406264 ; 
   reg __406264_406264;
   reg _406265_406265 ; 
   reg __406265_406265;
   reg _406266_406266 ; 
   reg __406266_406266;
   reg _406267_406267 ; 
   reg __406267_406267;
   reg _406268_406268 ; 
   reg __406268_406268;
   reg _406269_406269 ; 
   reg __406269_406269;
   reg _406270_406270 ; 
   reg __406270_406270;
   reg _406271_406271 ; 
   reg __406271_406271;
   reg _406272_406272 ; 
   reg __406272_406272;
   reg _406273_406273 ; 
   reg __406273_406273;
   reg _406274_406274 ; 
   reg __406274_406274;
   reg _406275_406275 ; 
   reg __406275_406275;
   reg _406276_406276 ; 
   reg __406276_406276;
   reg _406277_406277 ; 
   reg __406277_406277;
   reg _406278_406278 ; 
   reg __406278_406278;
   reg _406279_406279 ; 
   reg __406279_406279;
   reg _406280_406280 ; 
   reg __406280_406280;
   reg _406281_406281 ; 
   reg __406281_406281;
   reg _406282_406282 ; 
   reg __406282_406282;
   reg _406283_406283 ; 
   reg __406283_406283;
   reg _406284_406284 ; 
   reg __406284_406284;
   reg _406285_406285 ; 
   reg __406285_406285;
   reg _406286_406286 ; 
   reg __406286_406286;
   reg _406287_406287 ; 
   reg __406287_406287;
   reg _406288_406288 ; 
   reg __406288_406288;
   reg _406289_406289 ; 
   reg __406289_406289;
   reg _406290_406290 ; 
   reg __406290_406290;
   reg _406291_406291 ; 
   reg __406291_406291;
   reg _406292_406292 ; 
   reg __406292_406292;
   reg _406293_406293 ; 
   reg __406293_406293;
   reg _406294_406294 ; 
   reg __406294_406294;
   reg _406295_406295 ; 
   reg __406295_406295;
   reg _406296_406296 ; 
   reg __406296_406296;
   reg _406297_406297 ; 
   reg __406297_406297;
   reg _406298_406298 ; 
   reg __406298_406298;
   reg _406299_406299 ; 
   reg __406299_406299;
   reg _406300_406300 ; 
   reg __406300_406300;
   reg _406301_406301 ; 
   reg __406301_406301;
   reg _406302_406302 ; 
   reg __406302_406302;
   reg _406303_406303 ; 
   reg __406303_406303;
   reg _406304_406304 ; 
   reg __406304_406304;
   reg _406305_406305 ; 
   reg __406305_406305;
   reg _406306_406306 ; 
   reg __406306_406306;
   reg _406307_406307 ; 
   reg __406307_406307;
   reg _406308_406308 ; 
   reg __406308_406308;
   reg _406309_406309 ; 
   reg __406309_406309;
   reg _406310_406310 ; 
   reg __406310_406310;
   reg _406311_406311 ; 
   reg __406311_406311;
   reg _406312_406312 ; 
   reg __406312_406312;
   reg _406313_406313 ; 
   reg __406313_406313;
   reg _406314_406314 ; 
   reg __406314_406314;
   reg _406315_406315 ; 
   reg __406315_406315;
   reg _406316_406316 ; 
   reg __406316_406316;
   reg _406317_406317 ; 
   reg __406317_406317;
   reg _406318_406318 ; 
   reg __406318_406318;
   reg _406319_406319 ; 
   reg __406319_406319;
   reg _406320_406320 ; 
   reg __406320_406320;
   reg _406321_406321 ; 
   reg __406321_406321;
   reg _406322_406322 ; 
   reg __406322_406322;
   reg _406323_406323 ; 
   reg __406323_406323;
   reg _406324_406324 ; 
   reg __406324_406324;
   reg _406325_406325 ; 
   reg __406325_406325;
   reg _406326_406326 ; 
   reg __406326_406326;
   reg _406327_406327 ; 
   reg __406327_406327;
   reg _406328_406328 ; 
   reg __406328_406328;
   reg _406329_406329 ; 
   reg __406329_406329;
   reg _406330_406330 ; 
   reg __406330_406330;
   reg _406331_406331 ; 
   reg __406331_406331;
   reg _406332_406332 ; 
   reg __406332_406332;
   reg _406333_406333 ; 
   reg __406333_406333;
   reg _406334_406334 ; 
   reg __406334_406334;
   reg _406335_406335 ; 
   reg __406335_406335;
   reg _406336_406336 ; 
   reg __406336_406336;
   reg _406337_406337 ; 
   reg __406337_406337;
   reg _406338_406338 ; 
   reg __406338_406338;
   reg _406339_406339 ; 
   reg __406339_406339;
   reg _406340_406340 ; 
   reg __406340_406340;
   reg _406341_406341 ; 
   reg __406341_406341;
   reg _406342_406342 ; 
   reg __406342_406342;
   reg _406343_406343 ; 
   reg __406343_406343;
   reg _406344_406344 ; 
   reg __406344_406344;
   reg _406345_406345 ; 
   reg __406345_406345;
   reg _406346_406346 ; 
   reg __406346_406346;
   reg _406347_406347 ; 
   reg __406347_406347;
   reg _406348_406348 ; 
   reg __406348_406348;
   reg _406349_406349 ; 
   reg __406349_406349;
   reg _406350_406350 ; 
   reg __406350_406350;
   reg _406351_406351 ; 
   reg __406351_406351;
   reg _406352_406352 ; 
   reg __406352_406352;
   reg _406353_406353 ; 
   reg __406353_406353;
   reg _406354_406354 ; 
   reg __406354_406354;
   reg _406355_406355 ; 
   reg __406355_406355;
   reg _406356_406356 ; 
   reg __406356_406356;
   reg _406357_406357 ; 
   reg __406357_406357;
   reg _406358_406358 ; 
   reg __406358_406358;
   reg _406359_406359 ; 
   reg __406359_406359;
   reg _406360_406360 ; 
   reg __406360_406360;
   reg _406361_406361 ; 
   reg __406361_406361;
   reg _406362_406362 ; 
   reg __406362_406362;
   reg _406363_406363 ; 
   reg __406363_406363;
   reg _406364_406364 ; 
   reg __406364_406364;
   reg _406365_406365 ; 
   reg __406365_406365;
   reg _406366_406366 ; 
   reg __406366_406366;
   reg _406367_406367 ; 
   reg __406367_406367;
   reg _406368_406368 ; 
   reg __406368_406368;
   reg _406369_406369 ; 
   reg __406369_406369;
   reg _406370_406370 ; 
   reg __406370_406370;
   reg _406371_406371 ; 
   reg __406371_406371;
   reg _406372_406372 ; 
   reg __406372_406372;
   reg _406373_406373 ; 
   reg __406373_406373;
   reg _406374_406374 ; 
   reg __406374_406374;
   reg _406375_406375 ; 
   reg __406375_406375;
   reg _406376_406376 ; 
   reg __406376_406376;
   reg _406377_406377 ; 
   reg __406377_406377;
   reg _406378_406378 ; 
   reg __406378_406378;
   reg _406379_406379 ; 
   reg __406379_406379;
   reg _406380_406380 ; 
   reg __406380_406380;
   reg _406381_406381 ; 
   reg __406381_406381;
   reg _406382_406382 ; 
   reg __406382_406382;
   reg _406383_406383 ; 
   reg __406383_406383;
   reg _406384_406384 ; 
   reg __406384_406384;
   reg _406385_406385 ; 
   reg __406385_406385;
   reg _406386_406386 ; 
   reg __406386_406386;
   reg _406387_406387 ; 
   reg __406387_406387;
   reg _406388_406388 ; 
   reg __406388_406388;
   reg _406389_406389 ; 
   reg __406389_406389;
   reg _406390_406390 ; 
   reg __406390_406390;
   reg _406391_406391 ; 
   reg __406391_406391;
   reg _406392_406392 ; 
   reg __406392_406392;
   reg _406393_406393 ; 
   reg __406393_406393;
   reg _406394_406394 ; 
   reg __406394_406394;
   reg _406395_406395 ; 
   reg __406395_406395;
   reg _406396_406396 ; 
   reg __406396_406396;
   reg _406397_406397 ; 
   reg __406397_406397;
   reg _406398_406398 ; 
   reg __406398_406398;
   reg _406399_406399 ; 
   reg __406399_406399;
   reg _406400_406400 ; 
   reg __406400_406400;
   reg _406401_406401 ; 
   reg __406401_406401;
   reg _406402_406402 ; 
   reg __406402_406402;
   reg _406403_406403 ; 
   reg __406403_406403;
   reg _406404_406404 ; 
   reg __406404_406404;
   reg _406405_406405 ; 
   reg __406405_406405;
   reg _406406_406406 ; 
   reg __406406_406406;
   reg _406407_406407 ; 
   reg __406407_406407;
   reg _406408_406408 ; 
   reg __406408_406408;
   reg _406409_406409 ; 
   reg __406409_406409;
   reg _406410_406410 ; 
   reg __406410_406410;
   reg _406411_406411 ; 
   reg __406411_406411;
   reg _406412_406412 ; 
   reg __406412_406412;
   reg _406413_406413 ; 
   reg __406413_406413;
   reg _406414_406414 ; 
   reg __406414_406414;
   reg _406415_406415 ; 
   reg __406415_406415;
   reg _406416_406416 ; 
   reg __406416_406416;
   reg _406417_406417 ; 
   reg __406417_406417;
   reg _406418_406418 ; 
   reg __406418_406418;
   reg _406419_406419 ; 
   reg __406419_406419;
   reg _406420_406420 ; 
   reg __406420_406420;
   reg _406421_406421 ; 
   reg __406421_406421;
   reg _406422_406422 ; 
   reg __406422_406422;
   reg _406423_406423 ; 
   reg __406423_406423;
   reg _406424_406424 ; 
   reg __406424_406424;
   reg _406425_406425 ; 
   reg __406425_406425;
   reg _406426_406426 ; 
   reg __406426_406426;
   reg _406427_406427 ; 
   reg __406427_406427;
   reg _406428_406428 ; 
   reg __406428_406428;
   reg _406429_406429 ; 
   reg __406429_406429;
   reg _406430_406430 ; 
   reg __406430_406430;
   reg _406431_406431 ; 
   reg __406431_406431;
   reg _406432_406432 ; 
   reg __406432_406432;
   reg _406433_406433 ; 
   reg __406433_406433;
   reg _406434_406434 ; 
   reg __406434_406434;
   reg _406435_406435 ; 
   reg __406435_406435;
   reg _406436_406436 ; 
   reg __406436_406436;
   reg _406437_406437 ; 
   reg __406437_406437;
   reg _406438_406438 ; 
   reg __406438_406438;
   reg _406439_406439 ; 
   reg __406439_406439;
   reg _406440_406440 ; 
   reg __406440_406440;
   reg _406441_406441 ; 
   reg __406441_406441;
   reg _406442_406442 ; 
   reg __406442_406442;
   reg _406443_406443 ; 
   reg __406443_406443;
   reg _406444_406444 ; 
   reg __406444_406444;
   reg _406445_406445 ; 
   reg __406445_406445;
   reg _406446_406446 ; 
   reg __406446_406446;
   reg _406447_406447 ; 
   reg __406447_406447;
   reg _406448_406448 ; 
   reg __406448_406448;
   reg _406449_406449 ; 
   reg __406449_406449;
   reg _406450_406450 ; 
   reg __406450_406450;
   reg _406451_406451 ; 
   reg __406451_406451;
   reg _406452_406452 ; 
   reg __406452_406452;
   reg _406453_406453 ; 
   reg __406453_406453;
   reg _406454_406454 ; 
   reg __406454_406454;
   reg _406455_406455 ; 
   reg __406455_406455;
   reg _406456_406456 ; 
   reg __406456_406456;
   reg _406457_406457 ; 
   reg __406457_406457;
   reg _406458_406458 ; 
   reg __406458_406458;
   reg _406459_406459 ; 
   reg __406459_406459;
   reg _406460_406460 ; 
   reg __406460_406460;
   reg _406461_406461 ; 
   reg __406461_406461;
   reg _406462_406462 ; 
   reg __406462_406462;
   reg _406463_406463 ; 
   reg __406463_406463;
   reg _406464_406464 ; 
   reg __406464_406464;
   reg _406465_406465 ; 
   reg __406465_406465;
   reg _406466_406466 ; 
   reg __406466_406466;
   reg _406467_406467 ; 
   reg __406467_406467;
   reg _406468_406468 ; 
   reg __406468_406468;
   reg _406469_406469 ; 
   reg __406469_406469;
   reg _406470_406470 ; 
   reg __406470_406470;
   reg _406471_406471 ; 
   reg __406471_406471;
   reg _406472_406472 ; 
   reg __406472_406472;
   reg _406473_406473 ; 
   reg __406473_406473;
   reg _406474_406474 ; 
   reg __406474_406474;
   reg _406475_406475 ; 
   reg __406475_406475;
   reg _406476_406476 ; 
   reg __406476_406476;
   reg _406477_406477 ; 
   reg __406477_406477;
   reg _406478_406478 ; 
   reg __406478_406478;
   reg _406479_406479 ; 
   reg __406479_406479;
   reg _406480_406480 ; 
   reg __406480_406480;
   reg _406481_406481 ; 
   reg __406481_406481;
   reg _406482_406482 ; 
   reg __406482_406482;
   reg _406483_406483 ; 
   reg __406483_406483;
   reg _406484_406484 ; 
   reg __406484_406484;
   reg _406485_406485 ; 
   reg __406485_406485;
   reg _406486_406486 ; 
   reg __406486_406486;
   reg _406487_406487 ; 
   reg __406487_406487;
   reg _406488_406488 ; 
   reg __406488_406488;
   reg _406489_406489 ; 
   reg __406489_406489;
   reg _406490_406490 ; 
   reg __406490_406490;
   reg _406491_406491 ; 
   reg __406491_406491;
   reg _406492_406492 ; 
   reg __406492_406492;
   reg _406493_406493 ; 
   reg __406493_406493;
   reg _406494_406494 ; 
   reg __406494_406494;
   reg _406495_406495 ; 
   reg __406495_406495;
   reg _406496_406496 ; 
   reg __406496_406496;
   reg _406497_406497 ; 
   reg __406497_406497;
   reg _406498_406498 ; 
   reg __406498_406498;
   reg _406499_406499 ; 
   reg __406499_406499;
   reg _406500_406500 ; 
   reg __406500_406500;
   reg _406501_406501 ; 
   reg __406501_406501;
   reg _406502_406502 ; 
   reg __406502_406502;
   reg _406503_406503 ; 
   reg __406503_406503;
   reg _406504_406504 ; 
   reg __406504_406504;
   reg _406505_406505 ; 
   reg __406505_406505;
   reg _406506_406506 ; 
   reg __406506_406506;
   reg _406507_406507 ; 
   reg __406507_406507;
   reg _406508_406508 ; 
   reg __406508_406508;
   reg _406509_406509 ; 
   reg __406509_406509;
   reg _406510_406510 ; 
   reg __406510_406510;
   reg _406511_406511 ; 
   reg __406511_406511;
   reg _406512_406512 ; 
   reg __406512_406512;
   reg _406513_406513 ; 
   reg __406513_406513;
   reg _406514_406514 ; 
   reg __406514_406514;
   reg _406515_406515 ; 
   reg __406515_406515;
   reg _406516_406516 ; 
   reg __406516_406516;
   reg _406517_406517 ; 
   reg __406517_406517;
   reg _406518_406518 ; 
   reg __406518_406518;
   reg _406519_406519 ; 
   reg __406519_406519;
   reg _406520_406520 ; 
   reg __406520_406520;
   reg _406521_406521 ; 
   reg __406521_406521;
   reg _406522_406522 ; 
   reg __406522_406522;
   reg _406523_406523 ; 
   reg __406523_406523;
   reg _406524_406524 ; 
   reg __406524_406524;
   reg _406525_406525 ; 
   reg __406525_406525;
   reg _406526_406526 ; 
   reg __406526_406526;
   reg _406527_406527 ; 
   reg __406527_406527;
   reg _406528_406528 ; 
   reg __406528_406528;
   reg _406529_406529 ; 
   reg __406529_406529;
   reg _406530_406530 ; 
   reg __406530_406530;
   reg _406531_406531 ; 
   reg __406531_406531;
   reg _406532_406532 ; 
   reg __406532_406532;
   reg _406533_406533 ; 
   reg __406533_406533;
   reg _406534_406534 ; 
   reg __406534_406534;
   reg _406535_406535 ; 
   reg __406535_406535;
   reg _406536_406536 ; 
   reg __406536_406536;
   reg _406537_406537 ; 
   reg __406537_406537;
   reg _406538_406538 ; 
   reg __406538_406538;
   reg _406539_406539 ; 
   reg __406539_406539;
   reg _406540_406540 ; 
   reg __406540_406540;
   reg _406541_406541 ; 
   reg __406541_406541;
   reg _406542_406542 ; 
   reg __406542_406542;
   reg _406543_406543 ; 
   reg __406543_406543;
   reg _406544_406544 ; 
   reg __406544_406544;
   reg _406545_406545 ; 
   reg __406545_406545;
   reg _406546_406546 ; 
   reg __406546_406546;
   reg _406547_406547 ; 
   reg __406547_406547;
   reg _406548_406548 ; 
   reg __406548_406548;
   reg _406549_406549 ; 
   reg __406549_406549;
   reg _406550_406550 ; 
   reg __406550_406550;
   reg _406551_406551 ; 
   reg __406551_406551;
   reg _406552_406552 ; 
   reg __406552_406552;
   reg _406553_406553 ; 
   reg __406553_406553;
   reg _406554_406554 ; 
   reg __406554_406554;
   reg _406555_406555 ; 
   reg __406555_406555;
   reg _406556_406556 ; 
   reg __406556_406556;
   reg _406557_406557 ; 
   reg __406557_406557;
   reg _406558_406558 ; 
   reg __406558_406558;
   reg _406559_406559 ; 
   reg __406559_406559;
   reg _406560_406560 ; 
   reg __406560_406560;
   reg _406561_406561 ; 
   reg __406561_406561;
   reg _406562_406562 ; 
   reg __406562_406562;
   reg _406563_406563 ; 
   reg __406563_406563;
   reg _406564_406564 ; 
   reg __406564_406564;
   reg _406565_406565 ; 
   reg __406565_406565;
   reg _406566_406566 ; 
   reg __406566_406566;
   reg _406567_406567 ; 
   reg __406567_406567;
   reg _406568_406568 ; 
   reg __406568_406568;
   reg _406569_406569 ; 
   reg __406569_406569;
   reg _406570_406570 ; 
   reg __406570_406570;
   reg _406571_406571 ; 
   reg __406571_406571;
   reg _406572_406572 ; 
   reg __406572_406572;
   reg _406573_406573 ; 
   reg __406573_406573;
   reg _406574_406574 ; 
   reg __406574_406574;
   reg _406575_406575 ; 
   reg __406575_406575;
   reg _406576_406576 ; 
   reg __406576_406576;
   reg _406577_406577 ; 
   reg __406577_406577;
   reg _406578_406578 ; 
   reg __406578_406578;
   reg _406579_406579 ; 
   reg __406579_406579;
   reg _406580_406580 ; 
   reg __406580_406580;
   reg _406581_406581 ; 
   reg __406581_406581;
   reg _406582_406582 ; 
   reg __406582_406582;
   reg _406583_406583 ; 
   reg __406583_406583;
   reg _406584_406584 ; 
   reg __406584_406584;
   reg _406585_406585 ; 
   reg __406585_406585;
   reg _406586_406586 ; 
   reg __406586_406586;
   reg _406587_406587 ; 
   reg __406587_406587;
   reg _406588_406588 ; 
   reg __406588_406588;
   reg _406589_406589 ; 
   reg __406589_406589;
   reg _406590_406590 ; 
   reg __406590_406590;
   reg _406591_406591 ; 
   reg __406591_406591;
   reg _406592_406592 ; 
   reg __406592_406592;
   reg _406593_406593 ; 
   reg __406593_406593;
   reg _406594_406594 ; 
   reg __406594_406594;
   reg _406595_406595 ; 
   reg __406595_406595;
   reg _406596_406596 ; 
   reg __406596_406596;
   reg _406597_406597 ; 
   reg __406597_406597;
   reg _406598_406598 ; 
   reg __406598_406598;
   reg _406599_406599 ; 
   reg __406599_406599;
   reg _406600_406600 ; 
   reg __406600_406600;
   reg _406601_406601 ; 
   reg __406601_406601;
   reg _406602_406602 ; 
   reg __406602_406602;
   reg _406603_406603 ; 
   reg __406603_406603;
   reg _406604_406604 ; 
   reg __406604_406604;
   reg _406605_406605 ; 
   reg __406605_406605;
   reg _406606_406606 ; 
   reg __406606_406606;
   reg _406607_406607 ; 
   reg __406607_406607;
   reg _406608_406608 ; 
   reg __406608_406608;
   reg _406609_406609 ; 
   reg __406609_406609;
   reg _406610_406610 ; 
   reg __406610_406610;
   reg _406611_406611 ; 
   reg __406611_406611;
   reg _406612_406612 ; 
   reg __406612_406612;
   reg _406613_406613 ; 
   reg __406613_406613;
   reg _406614_406614 ; 
   reg __406614_406614;
   reg _406615_406615 ; 
   reg __406615_406615;
   reg _406616_406616 ; 
   reg __406616_406616;
   reg _406617_406617 ; 
   reg __406617_406617;
   reg _406618_406618 ; 
   reg __406618_406618;
   reg _406619_406619 ; 
   reg __406619_406619;
   reg _406620_406620 ; 
   reg __406620_406620;
   reg _406621_406621 ; 
   reg __406621_406621;
   reg _406622_406622 ; 
   reg __406622_406622;
   reg _406623_406623 ; 
   reg __406623_406623;
   reg _406624_406624 ; 
   reg __406624_406624;
   reg _406625_406625 ; 
   reg __406625_406625;
   reg _406626_406626 ; 
   reg __406626_406626;
   reg _406627_406627 ; 
   reg __406627_406627;
   reg _406628_406628 ; 
   reg __406628_406628;
   reg _406629_406629 ; 
   reg __406629_406629;
   reg _406630_406630 ; 
   reg __406630_406630;
   reg _406631_406631 ; 
   reg __406631_406631;
   reg _406632_406632 ; 
   reg __406632_406632;
   reg _406633_406633 ; 
   reg __406633_406633;
   reg _406634_406634 ; 
   reg __406634_406634;
   reg _406635_406635 ; 
   reg __406635_406635;
   reg _406636_406636 ; 
   reg __406636_406636;
   reg _406637_406637 ; 
   reg __406637_406637;
   reg _406638_406638 ; 
   reg __406638_406638;
   reg _406639_406639 ; 
   reg __406639_406639;
   reg _406640_406640 ; 
   reg __406640_406640;
   reg _406641_406641 ; 
   reg __406641_406641;
   reg _406642_406642 ; 
   reg __406642_406642;
   reg _406643_406643 ; 
   reg __406643_406643;
   reg _406644_406644 ; 
   reg __406644_406644;
   reg _406645_406645 ; 
   reg __406645_406645;
   reg _406646_406646 ; 
   reg __406646_406646;
   reg _406647_406647 ; 
   reg __406647_406647;
   reg _406648_406648 ; 
   reg __406648_406648;
   reg _406649_406649 ; 
   reg __406649_406649;
   reg _406650_406650 ; 
   reg __406650_406650;
   reg _406651_406651 ; 
   reg __406651_406651;
   reg _406652_406652 ; 
   reg __406652_406652;
   reg _406653_406653 ; 
   reg __406653_406653;
   reg _406654_406654 ; 
   reg __406654_406654;
   reg _406655_406655 ; 
   reg __406655_406655;
   reg _406656_406656 ; 
   reg __406656_406656;
   reg _406657_406657 ; 
   reg __406657_406657;
   reg _406658_406658 ; 
   reg __406658_406658;
   reg _406659_406659 ; 
   reg __406659_406659;
   reg _406660_406660 ; 
   reg __406660_406660;
   reg _406661_406661 ; 
   reg __406661_406661;
   reg _406662_406662 ; 
   reg __406662_406662;
   reg _406663_406663 ; 
   reg __406663_406663;
   reg _406664_406664 ; 
   reg __406664_406664;
   reg _406665_406665 ; 
   reg __406665_406665;
   reg _406666_406666 ; 
   reg __406666_406666;
   reg _406667_406667 ; 
   reg __406667_406667;
   reg _406668_406668 ; 
   reg __406668_406668;
   reg _406669_406669 ; 
   reg __406669_406669;
   reg _406670_406670 ; 
   reg __406670_406670;
   reg _406671_406671 ; 
   reg __406671_406671;
   reg _406672_406672 ; 
   reg __406672_406672;
   reg _406673_406673 ; 
   reg __406673_406673;
   reg _406674_406674 ; 
   reg __406674_406674;
   reg _406675_406675 ; 
   reg __406675_406675;
   reg _406676_406676 ; 
   reg __406676_406676;
   reg _406677_406677 ; 
   reg __406677_406677;
   reg _406678_406678 ; 
   reg __406678_406678;
   reg _406679_406679 ; 
   reg __406679_406679;
   reg _406680_406680 ; 
   reg __406680_406680;
   reg _406681_406681 ; 
   reg __406681_406681;
   reg _406682_406682 ; 
   reg __406682_406682;
   reg _406683_406683 ; 
   reg __406683_406683;
   reg _406684_406684 ; 
   reg __406684_406684;
   reg _406685_406685 ; 
   reg __406685_406685;
   reg _406686_406686 ; 
   reg __406686_406686;
   reg _406687_406687 ; 
   reg __406687_406687;
   reg _406688_406688 ; 
   reg __406688_406688;
   reg _406689_406689 ; 
   reg __406689_406689;
   reg _406690_406690 ; 
   reg __406690_406690;
   reg _406691_406691 ; 
   reg __406691_406691;
   reg _406692_406692 ; 
   reg __406692_406692;
   reg _406693_406693 ; 
   reg __406693_406693;
   reg _406694_406694 ; 
   reg __406694_406694;
   reg _406695_406695 ; 
   reg __406695_406695;
   reg _406696_406696 ; 
   reg __406696_406696;
   reg _406697_406697 ; 
   reg __406697_406697;
   reg _406698_406698 ; 
   reg __406698_406698;
   reg _406699_406699 ; 
   reg __406699_406699;
   reg _406700_406700 ; 
   reg __406700_406700;
   reg _406701_406701 ; 
   reg __406701_406701;
   reg _406702_406702 ; 
   reg __406702_406702;
   reg _406703_406703 ; 
   reg __406703_406703;
   reg _406704_406704 ; 
   reg __406704_406704;
   reg _406705_406705 ; 
   reg __406705_406705;
   reg _406706_406706 ; 
   reg __406706_406706;
   reg _406707_406707 ; 
   reg __406707_406707;
   reg _406708_406708 ; 
   reg __406708_406708;
   reg _406709_406709 ; 
   reg __406709_406709;
   reg _406710_406710 ; 
   reg __406710_406710;
   reg _406711_406711 ; 
   reg __406711_406711;
   reg _406712_406712 ; 
   reg __406712_406712;
   reg _406713_406713 ; 
   reg __406713_406713;
   reg _406714_406714 ; 
   reg __406714_406714;
   reg _406715_406715 ; 
   reg __406715_406715;
   reg _406716_406716 ; 
   reg __406716_406716;
   reg _406717_406717 ; 
   reg __406717_406717;
   reg _406718_406718 ; 
   reg __406718_406718;
   reg _406719_406719 ; 
   reg __406719_406719;
   reg _406720_406720 ; 
   reg __406720_406720;
   reg _406721_406721 ; 
   reg __406721_406721;
   reg _406722_406722 ; 
   reg __406722_406722;
   reg _406723_406723 ; 
   reg __406723_406723;
   reg _406724_406724 ; 
   reg __406724_406724;
   reg _406725_406725 ; 
   reg __406725_406725;
   reg _406726_406726 ; 
   reg __406726_406726;
   reg _406727_406727 ; 
   reg __406727_406727;
   reg _406728_406728 ; 
   reg __406728_406728;
   reg _406729_406729 ; 
   reg __406729_406729;
   reg _406730_406730 ; 
   reg __406730_406730;
   reg _406731_406731 ; 
   reg __406731_406731;
   reg _406732_406732 ; 
   reg __406732_406732;
   reg _406733_406733 ; 
   reg __406733_406733;
   reg _406734_406734 ; 
   reg __406734_406734;
   reg _406735_406735 ; 
   reg __406735_406735;
   reg _406736_406736 ; 
   reg __406736_406736;
   reg _406737_406737 ; 
   reg __406737_406737;
   reg _406738_406738 ; 
   reg __406738_406738;
   reg _406739_406739 ; 
   reg __406739_406739;
   reg _406740_406740 ; 
   reg __406740_406740;
   reg _406741_406741 ; 
   reg __406741_406741;
   reg _406742_406742 ; 
   reg __406742_406742;
   reg _406743_406743 ; 
   reg __406743_406743;
   reg _406744_406744 ; 
   reg __406744_406744;
   reg _406745_406745 ; 
   reg __406745_406745;
   reg _406746_406746 ; 
   reg __406746_406746;
   reg _406747_406747 ; 
   reg __406747_406747;
   reg _406748_406748 ; 
   reg __406748_406748;
   reg _406749_406749 ; 
   reg __406749_406749;
   reg _406750_406750 ; 
   reg __406750_406750;
   reg _406751_406751 ; 
   reg __406751_406751;
   reg _406752_406752 ; 
   reg __406752_406752;
   reg _406753_406753 ; 
   reg __406753_406753;
   reg _406754_406754 ; 
   reg __406754_406754;
   reg _406755_406755 ; 
   reg __406755_406755;
   reg _406756_406756 ; 
   reg __406756_406756;
   reg _406757_406757 ; 
   reg __406757_406757;
   reg _406758_406758 ; 
   reg __406758_406758;
   reg _406759_406759 ; 
   reg __406759_406759;
   reg _406760_406760 ; 
   reg __406760_406760;
   reg _406761_406761 ; 
   reg __406761_406761;
   reg _406762_406762 ; 
   reg __406762_406762;
   reg _406763_406763 ; 
   reg __406763_406763;
   reg _406764_406764 ; 
   reg __406764_406764;
   reg _406765_406765 ; 
   reg __406765_406765;
   reg _406766_406766 ; 
   reg __406766_406766;
   reg _406767_406767 ; 
   reg __406767_406767;
   reg _406768_406768 ; 
   reg __406768_406768;
   reg _406769_406769 ; 
   reg __406769_406769;
   reg _406770_406770 ; 
   reg __406770_406770;
   reg _406771_406771 ; 
   reg __406771_406771;
   reg _406772_406772 ; 
   reg __406772_406772;
   reg _406773_406773 ; 
   reg __406773_406773;
   reg _406774_406774 ; 
   reg __406774_406774;
   reg _406775_406775 ; 
   reg __406775_406775;
   reg _406776_406776 ; 
   reg __406776_406776;
   reg _406777_406777 ; 
   reg __406777_406777;
   reg _406778_406778 ; 
   reg __406778_406778;
   reg _406779_406779 ; 
   reg __406779_406779;
   reg _406780_406780 ; 
   reg __406780_406780;
   reg _406781_406781 ; 
   reg __406781_406781;
   reg _406782_406782 ; 
   reg __406782_406782;
   reg _406783_406783 ; 
   reg __406783_406783;
   reg _406784_406784 ; 
   reg __406784_406784;
   reg _406785_406785 ; 
   reg __406785_406785;
   reg _406786_406786 ; 
   reg __406786_406786;
   reg _406787_406787 ; 
   reg __406787_406787;
   reg _406788_406788 ; 
   reg __406788_406788;
   reg _406789_406789 ; 
   reg __406789_406789;
   reg _406790_406790 ; 
   reg __406790_406790;
   reg _406791_406791 ; 
   reg __406791_406791;
   reg _406792_406792 ; 
   reg __406792_406792;
   reg _406793_406793 ; 
   reg __406793_406793;
   reg _406794_406794 ; 
   reg __406794_406794;
   reg _406795_406795 ; 
   reg __406795_406795;
   reg _406796_406796 ; 
   reg __406796_406796;
   reg _406797_406797 ; 
   reg __406797_406797;
   reg _406798_406798 ; 
   reg __406798_406798;
   reg _406799_406799 ; 
   reg __406799_406799;
   reg _406800_406800 ; 
   reg __406800_406800;
   reg _406801_406801 ; 
   reg __406801_406801;
   reg _406802_406802 ; 
   reg __406802_406802;
   reg _406803_406803 ; 
   reg __406803_406803;
   reg _406804_406804 ; 
   reg __406804_406804;
   reg _406805_406805 ; 
   reg __406805_406805;
   reg _406806_406806 ; 
   reg __406806_406806;
   reg _406807_406807 ; 
   reg __406807_406807;
   reg _406808_406808 ; 
   reg __406808_406808;
   reg _406809_406809 ; 
   reg __406809_406809;
   reg _406810_406810 ; 
   reg __406810_406810;
   reg _406811_406811 ; 
   reg __406811_406811;
   reg _406812_406812 ; 
   reg __406812_406812;
   reg _406813_406813 ; 
   reg __406813_406813;
   reg _406814_406814 ; 
   reg __406814_406814;
   reg _406815_406815 ; 
   reg __406815_406815;
   reg _406816_406816 ; 
   reg __406816_406816;
   reg _406817_406817 ; 
   reg __406817_406817;
   reg _406818_406818 ; 
   reg __406818_406818;
   reg _406819_406819 ; 
   reg __406819_406819;
   reg _406820_406820 ; 
   reg __406820_406820;
   reg _406821_406821 ; 
   reg __406821_406821;
   reg _406822_406822 ; 
   reg __406822_406822;
   reg _406823_406823 ; 
   reg __406823_406823;
   reg _406824_406824 ; 
   reg __406824_406824;
   reg _406825_406825 ; 
   reg __406825_406825;
   reg _406826_406826 ; 
   reg __406826_406826;
   reg _406827_406827 ; 
   reg __406827_406827;
   reg _406828_406828 ; 
   reg __406828_406828;
   reg _406829_406829 ; 
   reg __406829_406829;
   reg _406830_406830 ; 
   reg __406830_406830;
   reg _406831_406831 ; 
   reg __406831_406831;
   reg _406832_406832 ; 
   reg __406832_406832;
   reg _406833_406833 ; 
   reg __406833_406833;
   reg _406834_406834 ; 
   reg __406834_406834;
   reg _406835_406835 ; 
   reg __406835_406835;
   reg _406836_406836 ; 
   reg __406836_406836;
   reg _406837_406837 ; 
   reg __406837_406837;
   reg _406838_406838 ; 
   reg __406838_406838;
   reg _406839_406839 ; 
   reg __406839_406839;
   reg _406840_406840 ; 
   reg __406840_406840;
   reg _406841_406841 ; 
   reg __406841_406841;
   reg _406842_406842 ; 
   reg __406842_406842;
   reg _406843_406843 ; 
   reg __406843_406843;
   reg _406844_406844 ; 
   reg __406844_406844;
   reg _406845_406845 ; 
   reg __406845_406845;
   reg _406846_406846 ; 
   reg __406846_406846;
   reg _406847_406847 ; 
   reg __406847_406847;
   reg _406848_406848 ; 
   reg __406848_406848;
   reg _406849_406849 ; 
   reg __406849_406849;
   reg _406850_406850 ; 
   reg __406850_406850;
   reg _406851_406851 ; 
   reg __406851_406851;
   reg _406852_406852 ; 
   reg __406852_406852;
   reg _406853_406853 ; 
   reg __406853_406853;
   reg _406854_406854 ; 
   reg __406854_406854;
   reg _406855_406855 ; 
   reg __406855_406855;
   reg _406856_406856 ; 
   reg __406856_406856;
   reg _406857_406857 ; 
   reg __406857_406857;
   reg _406858_406858 ; 
   reg __406858_406858;
   reg _406859_406859 ; 
   reg __406859_406859;
   reg _406860_406860 ; 
   reg __406860_406860;
   reg _406861_406861 ; 
   reg __406861_406861;
   reg _406862_406862 ; 
   reg __406862_406862;
   reg _406863_406863 ; 
   reg __406863_406863;
   reg _406864_406864 ; 
   reg __406864_406864;
   reg _406865_406865 ; 
   reg __406865_406865;
   reg _406866_406866 ; 
   reg __406866_406866;
   reg _406867_406867 ; 
   reg __406867_406867;
   reg _406868_406868 ; 
   reg __406868_406868;
   reg _406869_406869 ; 
   reg __406869_406869;
   reg _406870_406870 ; 
   reg __406870_406870;
   reg _406871_406871 ; 
   reg __406871_406871;
   reg _406872_406872 ; 
   reg __406872_406872;
   reg _406873_406873 ; 
   reg __406873_406873;
   reg _406874_406874 ; 
   reg __406874_406874;
   reg _406875_406875 ; 
   reg __406875_406875;
   reg _406876_406876 ; 
   reg __406876_406876;
   reg _406877_406877 ; 
   reg __406877_406877;
   reg _406878_406878 ; 
   reg __406878_406878;
   reg _406879_406879 ; 
   reg __406879_406879;
   reg _406880_406880 ; 
   reg __406880_406880;
   reg _406881_406881 ; 
   reg __406881_406881;
   reg _406882_406882 ; 
   reg __406882_406882;
   reg _406883_406883 ; 
   reg __406883_406883;
   reg _406884_406884 ; 
   reg __406884_406884;
   reg _406885_406885 ; 
   reg __406885_406885;
   reg _406886_406886 ; 
   reg __406886_406886;
   reg _406887_406887 ; 
   reg __406887_406887;
   reg _406888_406888 ; 
   reg __406888_406888;
   reg _406889_406889 ; 
   reg __406889_406889;
   reg _406890_406890 ; 
   reg __406890_406890;
   reg _406891_406891 ; 
   reg __406891_406891;
   reg _406892_406892 ; 
   reg __406892_406892;
   reg _406893_406893 ; 
   reg __406893_406893;
   reg _406894_406894 ; 
   reg __406894_406894;
   reg _406895_406895 ; 
   reg __406895_406895;
   reg _406896_406896 ; 
   reg __406896_406896;
   reg _406897_406897 ; 
   reg __406897_406897;
   reg _406898_406898 ; 
   reg __406898_406898;
   reg _406899_406899 ; 
   reg __406899_406899;
   reg _406900_406900 ; 
   reg __406900_406900;
   reg _406901_406901 ; 
   reg __406901_406901;
   reg _406902_406902 ; 
   reg __406902_406902;
   reg _406903_406903 ; 
   reg __406903_406903;
   reg _406904_406904 ; 
   reg __406904_406904;
   reg _406905_406905 ; 
   reg __406905_406905;
   reg _406906_406906 ; 
   reg __406906_406906;
   reg _406907_406907 ; 
   reg __406907_406907;
   reg _406908_406908 ; 
   reg __406908_406908;
   reg _406909_406909 ; 
   reg __406909_406909;
   reg _406910_406910 ; 
   reg __406910_406910;
   reg _406911_406911 ; 
   reg __406911_406911;
   reg _406912_406912 ; 
   reg __406912_406912;
   reg _406913_406913 ; 
   reg __406913_406913;
   reg _406914_406914 ; 
   reg __406914_406914;
   reg _406915_406915 ; 
   reg __406915_406915;
   reg _406916_406916 ; 
   reg __406916_406916;
   reg _406917_406917 ; 
   reg __406917_406917;
   reg _406918_406918 ; 
   reg __406918_406918;
   reg _406919_406919 ; 
   reg __406919_406919;
   reg _406920_406920 ; 
   reg __406920_406920;
   reg _406921_406921 ; 
   reg __406921_406921;
   reg _406922_406922 ; 
   reg __406922_406922;
   reg _406923_406923 ; 
   reg __406923_406923;
   reg _406924_406924 ; 
   reg __406924_406924;
   reg _406925_406925 ; 
   reg __406925_406925;
   reg _406926_406926 ; 
   reg __406926_406926;
   reg _406927_406927 ; 
   reg __406927_406927;
   reg _406928_406928 ; 
   reg __406928_406928;
   reg _406929_406929 ; 
   reg __406929_406929;
   reg _406930_406930 ; 
   reg __406930_406930;
   reg _406931_406931 ; 
   reg __406931_406931;
   reg _406932_406932 ; 
   reg __406932_406932;
   reg _406933_406933 ; 
   reg __406933_406933;
   reg _406934_406934 ; 
   reg __406934_406934;
   reg _406935_406935 ; 
   reg __406935_406935;
   reg _406936_406936 ; 
   reg __406936_406936;
   reg _406937_406937 ; 
   reg __406937_406937;
   reg _406938_406938 ; 
   reg __406938_406938;
   reg _406939_406939 ; 
   reg __406939_406939;
   reg _406940_406940 ; 
   reg __406940_406940;
   reg _406941_406941 ; 
   reg __406941_406941;
   reg _406942_406942 ; 
   reg __406942_406942;
   reg _406943_406943 ; 
   reg __406943_406943;
   reg _406944_406944 ; 
   reg __406944_406944;
   reg _406945_406945 ; 
   reg __406945_406945;
   reg _406946_406946 ; 
   reg __406946_406946;
   reg _406947_406947 ; 
   reg __406947_406947;
   reg _406948_406948 ; 
   reg __406948_406948;
   reg _406949_406949 ; 
   reg __406949_406949;
   reg _406950_406950 ; 
   reg __406950_406950;
   reg _406951_406951 ; 
   reg __406951_406951;
   reg _406952_406952 ; 
   reg __406952_406952;
   reg _406953_406953 ; 
   reg __406953_406953;
   reg _406954_406954 ; 
   reg __406954_406954;
   reg _406955_406955 ; 
   reg __406955_406955;
   reg _406956_406956 ; 
   reg __406956_406956;
   reg _406957_406957 ; 
   reg __406957_406957;
   reg _406958_406958 ; 
   reg __406958_406958;
   reg _406959_406959 ; 
   reg __406959_406959;
   reg _406960_406960 ; 
   reg __406960_406960;
   reg _406961_406961 ; 
   reg __406961_406961;
   reg _406962_406962 ; 
   reg __406962_406962;
   reg _406963_406963 ; 
   reg __406963_406963;
   reg _406964_406964 ; 
   reg __406964_406964;
   reg _406965_406965 ; 
   reg __406965_406965;
   reg _406966_406966 ; 
   reg __406966_406966;
   reg _406967_406967 ; 
   reg __406967_406967;
   reg _406968_406968 ; 
   reg __406968_406968;
   reg _406969_406969 ; 
   reg __406969_406969;
   reg _406970_406970 ; 
   reg __406970_406970;
   reg _406971_406971 ; 
   reg __406971_406971;
   reg _406972_406972 ; 
   reg __406972_406972;
   reg _406973_406973 ; 
   reg __406973_406973;
   reg _406974_406974 ; 
   reg __406974_406974;
   reg _406975_406975 ; 
   reg __406975_406975;
   reg _406976_406976 ; 
   reg __406976_406976;
   reg _406977_406977 ; 
   reg __406977_406977;
   reg _406978_406978 ; 
   reg __406978_406978;
   reg _406979_406979 ; 
   reg __406979_406979;
   reg _406980_406980 ; 
   reg __406980_406980;
   reg _406981_406981 ; 
   reg __406981_406981;
   reg _406982_406982 ; 
   reg __406982_406982;
   reg _406983_406983 ; 
   reg __406983_406983;
   reg _406984_406984 ; 
   reg __406984_406984;
   reg _406985_406985 ; 
   reg __406985_406985;
   reg _406986_406986 ; 
   reg __406986_406986;
   reg _406987_406987 ; 
   reg __406987_406987;
   reg _406988_406988 ; 
   reg __406988_406988;
   reg _406989_406989 ; 
   reg __406989_406989;
   reg _406990_406990 ; 
   reg __406990_406990;
   reg _406991_406991 ; 
   reg __406991_406991;
   reg _406992_406992 ; 
   reg __406992_406992;
   reg _406993_406993 ; 
   reg __406993_406993;
   reg _406994_406994 ; 
   reg __406994_406994;
   reg _406995_406995 ; 
   reg __406995_406995;
   reg _406996_406996 ; 
   reg __406996_406996;
   reg _406997_406997 ; 
   reg __406997_406997;
   reg _406998_406998 ; 
   reg __406998_406998;
   reg _406999_406999 ; 
   reg __406999_406999;
   reg _407000_407000 ; 
   reg __407000_407000;
   reg _407001_407001 ; 
   reg __407001_407001;
   reg _407002_407002 ; 
   reg __407002_407002;
   reg _407003_407003 ; 
   reg __407003_407003;
   reg _407004_407004 ; 
   reg __407004_407004;
   reg _407005_407005 ; 
   reg __407005_407005;
   reg _407006_407006 ; 
   reg __407006_407006;
   reg _407007_407007 ; 
   reg __407007_407007;
   reg _407008_407008 ; 
   reg __407008_407008;
   reg _407009_407009 ; 
   reg __407009_407009;
   reg _407010_407010 ; 
   reg __407010_407010;
   reg _407011_407011 ; 
   reg __407011_407011;
   reg _407012_407012 ; 
   reg __407012_407012;
   reg _407013_407013 ; 
   reg __407013_407013;
   reg _407014_407014 ; 
   reg __407014_407014;
   reg _407015_407015 ; 
   reg __407015_407015;
   reg _407016_407016 ; 
   reg __407016_407016;
   reg _407017_407017 ; 
   reg __407017_407017;
   reg _407018_407018 ; 
   reg __407018_407018;
   reg _407019_407019 ; 
   reg __407019_407019;
   reg _407020_407020 ; 
   reg __407020_407020;
   reg _407021_407021 ; 
   reg __407021_407021;
   reg _407022_407022 ; 
   reg __407022_407022;
   reg _407023_407023 ; 
   reg __407023_407023;
   reg _407024_407024 ; 
   reg __407024_407024;
   reg _407025_407025 ; 
   reg __407025_407025;
   reg _407026_407026 ; 
   reg __407026_407026;
   reg _407027_407027 ; 
   reg __407027_407027;
   reg _407028_407028 ; 
   reg __407028_407028;
   reg _407029_407029 ; 
   reg __407029_407029;
   reg _407030_407030 ; 
   reg __407030_407030;
   reg _407031_407031 ; 
   reg __407031_407031;
   reg _407032_407032 ; 
   reg __407032_407032;
   reg _407033_407033 ; 
   reg __407033_407033;
   reg _407034_407034 ; 
   reg __407034_407034;
   reg _407035_407035 ; 
   reg __407035_407035;
   reg _407036_407036 ; 
   reg __407036_407036;
   reg _407037_407037 ; 
   reg __407037_407037;
   reg _407038_407038 ; 
   reg __407038_407038;
   reg _407039_407039 ; 
   reg __407039_407039;
   reg _407040_407040 ; 
   reg __407040_407040;
   reg _407041_407041 ; 
   reg __407041_407041;
   reg _407042_407042 ; 
   reg __407042_407042;
   reg _407043_407043 ; 
   reg __407043_407043;
   reg _407044_407044 ; 
   reg __407044_407044;
   reg _407045_407045 ; 
   reg __407045_407045;
   reg _407046_407046 ; 
   reg __407046_407046;
   reg _407047_407047 ; 
   reg __407047_407047;
   reg _407048_407048 ; 
   reg __407048_407048;
   reg _407049_407049 ; 
   reg __407049_407049;
   reg _407050_407050 ; 
   reg __407050_407050;
   reg _407051_407051 ; 
   reg __407051_407051;
   reg _407052_407052 ; 
   reg __407052_407052;
   reg _407053_407053 ; 
   reg __407053_407053;
   reg _407054_407054 ; 
   reg __407054_407054;
   reg _407055_407055 ; 
   reg __407055_407055;
   reg _407056_407056 ; 
   reg __407056_407056;
   reg _407057_407057 ; 
   reg __407057_407057;
   reg _407058_407058 ; 
   reg __407058_407058;
   reg _407059_407059 ; 
   reg __407059_407059;
   reg _407060_407060 ; 
   reg __407060_407060;
   reg _407061_407061 ; 
   reg __407061_407061;
   reg _407062_407062 ; 
   reg __407062_407062;
   reg _407063_407063 ; 
   reg __407063_407063;
   reg _407064_407064 ; 
   reg __407064_407064;
   reg _407065_407065 ; 
   reg __407065_407065;
   reg _407066_407066 ; 
   reg __407066_407066;
   reg _407067_407067 ; 
   reg __407067_407067;
   reg _407068_407068 ; 
   reg __407068_407068;
   reg _407069_407069 ; 
   reg __407069_407069;
   reg _407070_407070 ; 
   reg __407070_407070;
   reg _407071_407071 ; 
   reg __407071_407071;
   reg _407072_407072 ; 
   reg __407072_407072;
   reg _407073_407073 ; 
   reg __407073_407073;
   reg _407074_407074 ; 
   reg __407074_407074;
   reg _407075_407075 ; 
   reg __407075_407075;
   reg _407076_407076 ; 
   reg __407076_407076;
   reg _407077_407077 ; 
   reg __407077_407077;
   reg _407078_407078 ; 
   reg __407078_407078;
   reg _407079_407079 ; 
   reg __407079_407079;
   reg _407080_407080 ; 
   reg __407080_407080;
   reg _407081_407081 ; 
   reg __407081_407081;
   reg _407082_407082 ; 
   reg __407082_407082;
   reg _407083_407083 ; 
   reg __407083_407083;
   reg _407084_407084 ; 
   reg __407084_407084;
   reg _407085_407085 ; 
   reg __407085_407085;
   reg _407086_407086 ; 
   reg __407086_407086;
   reg _407087_407087 ; 
   reg __407087_407087;
   reg _407088_407088 ; 
   reg __407088_407088;
   reg _407089_407089 ; 
   reg __407089_407089;
   reg _407090_407090 ; 
   reg __407090_407090;
   reg _407091_407091 ; 
   reg __407091_407091;
   reg _407092_407092 ; 
   reg __407092_407092;
   reg _407093_407093 ; 
   reg __407093_407093;
   reg _407094_407094 ; 
   reg __407094_407094;
   reg _407095_407095 ; 
   reg __407095_407095;
   reg _407096_407096 ; 
   reg __407096_407096;
   reg _407097_407097 ; 
   reg __407097_407097;
   reg _407098_407098 ; 
   reg __407098_407098;
   reg _407099_407099 ; 
   reg __407099_407099;
   reg _407100_407100 ; 
   reg __407100_407100;
   reg _407101_407101 ; 
   reg __407101_407101;
   reg _407102_407102 ; 
   reg __407102_407102;
   reg _407103_407103 ; 
   reg __407103_407103;
   reg _407104_407104 ; 
   reg __407104_407104;
   reg _407105_407105 ; 
   reg __407105_407105;
   reg _407106_407106 ; 
   reg __407106_407106;
   reg _407107_407107 ; 
   reg __407107_407107;
   reg _407108_407108 ; 
   reg __407108_407108;
   reg _407109_407109 ; 
   reg __407109_407109;
   reg _407110_407110 ; 
   reg __407110_407110;
   reg _407111_407111 ; 
   reg __407111_407111;
   reg _407112_407112 ; 
   reg __407112_407112;
   reg _407113_407113 ; 
   reg __407113_407113;
   reg _407114_407114 ; 
   reg __407114_407114;
   reg _407115_407115 ; 
   reg __407115_407115;
   reg _407116_407116 ; 
   reg __407116_407116;
   reg _407117_407117 ; 
   reg __407117_407117;
   reg _407118_407118 ; 
   reg __407118_407118;
   reg _407119_407119 ; 
   reg __407119_407119;
   reg _407120_407120 ; 
   reg __407120_407120;
   reg _407121_407121 ; 
   reg __407121_407121;
   reg _407122_407122 ; 
   reg __407122_407122;
   reg _407123_407123 ; 
   reg __407123_407123;
   reg _407124_407124 ; 
   reg __407124_407124;
   reg _407125_407125 ; 
   reg __407125_407125;
   reg _407126_407126 ; 
   reg __407126_407126;
   reg _407127_407127 ; 
   reg __407127_407127;
   reg _407128_407128 ; 
   reg __407128_407128;
   reg _407129_407129 ; 
   reg __407129_407129;
   reg _407130_407130 ; 
   reg __407130_407130;
   reg _407131_407131 ; 
   reg __407131_407131;
   reg _407132_407132 ; 
   reg __407132_407132;
   reg _407133_407133 ; 
   reg __407133_407133;
   reg _407134_407134 ; 
   reg __407134_407134;
   reg _407135_407135 ; 
   reg __407135_407135;
   reg _407136_407136 ; 
   reg __407136_407136;
   reg _407137_407137 ; 
   reg __407137_407137;
   reg _407138_407138 ; 
   reg __407138_407138;
   reg _407139_407139 ; 
   reg __407139_407139;
   reg _407140_407140 ; 
   reg __407140_407140;
   reg _407141_407141 ; 
   reg __407141_407141;
   reg _407142_407142 ; 
   reg __407142_407142;
   reg _407143_407143 ; 
   reg __407143_407143;
   reg _407144_407144 ; 
   reg __407144_407144;
   reg _407145_407145 ; 
   reg __407145_407145;
   reg _407146_407146 ; 
   reg __407146_407146;
   reg _407147_407147 ; 
   reg __407147_407147;
   reg _407148_407148 ; 
   reg __407148_407148;
   reg _407149_407149 ; 
   reg __407149_407149;
   reg _407150_407150 ; 
   reg __407150_407150;
   reg _407151_407151 ; 
   reg __407151_407151;
   reg _407152_407152 ; 
   reg __407152_407152;
   reg _407153_407153 ; 
   reg __407153_407153;
   reg _407154_407154 ; 
   reg __407154_407154;
   reg _407155_407155 ; 
   reg __407155_407155;
   reg _407156_407156 ; 
   reg __407156_407156;
   reg _407157_407157 ; 
   reg __407157_407157;
   reg _407158_407158 ; 
   reg __407158_407158;
   reg _407159_407159 ; 
   reg __407159_407159;
   reg _407160_407160 ; 
   reg __407160_407160;
   reg _407161_407161 ; 
   reg __407161_407161;
   reg _407162_407162 ; 
   reg __407162_407162;
   reg _407163_407163 ; 
   reg __407163_407163;
   reg _407164_407164 ; 
   reg __407164_407164;
   reg _407165_407165 ; 
   reg __407165_407165;
   reg _407166_407166 ; 
   reg __407166_407166;
   reg _407167_407167 ; 
   reg __407167_407167;
   reg _407168_407168 ; 
   reg __407168_407168;
   reg _407169_407169 ; 
   reg __407169_407169;
   reg _407170_407170 ; 
   reg __407170_407170;
   reg _407171_407171 ; 
   reg __407171_407171;
   reg _407172_407172 ; 
   reg __407172_407172;
   reg _407173_407173 ; 
   reg __407173_407173;
   reg _407174_407174 ; 
   reg __407174_407174;
   reg _407175_407175 ; 
   reg __407175_407175;
   reg _407176_407176 ; 
   reg __407176_407176;
   reg _407177_407177 ; 
   reg __407177_407177;
   reg _407178_407178 ; 
   reg __407178_407178;
   reg _407179_407179 ; 
   reg __407179_407179;
   reg _407180_407180 ; 
   reg __407180_407180;
   reg _407181_407181 ; 
   reg __407181_407181;
   reg _407182_407182 ; 
   reg __407182_407182;
   reg _407183_407183 ; 
   reg __407183_407183;
   reg _407184_407184 ; 
   reg __407184_407184;
   reg _407185_407185 ; 
   reg __407185_407185;
   reg _407186_407186 ; 
   reg __407186_407186;
   reg _407187_407187 ; 
   reg __407187_407187;
   reg _407188_407188 ; 
   reg __407188_407188;
   reg _407189_407189 ; 
   reg __407189_407189;
   reg _407190_407190 ; 
   reg __407190_407190;
   reg _407191_407191 ; 
   reg __407191_407191;
   reg _407192_407192 ; 
   reg __407192_407192;
   reg _407193_407193 ; 
   reg __407193_407193;
   reg _407194_407194 ; 
   reg __407194_407194;
   reg _407195_407195 ; 
   reg __407195_407195;
   reg _407196_407196 ; 
   reg __407196_407196;
   reg _407197_407197 ; 
   reg __407197_407197;
   reg _407198_407198 ; 
   reg __407198_407198;
   reg _407199_407199 ; 
   reg __407199_407199;
   reg _407200_407200 ; 
   reg __407200_407200;
   reg _407201_407201 ; 
   reg __407201_407201;
   reg _407202_407202 ; 
   reg __407202_407202;
   reg _407203_407203 ; 
   reg __407203_407203;
   reg _407204_407204 ; 
   reg __407204_407204;
   reg _407205_407205 ; 
   reg __407205_407205;
   reg _407206_407206 ; 
   reg __407206_407206;
   reg _407207_407207 ; 
   reg __407207_407207;
   reg _407208_407208 ; 
   reg __407208_407208;
   reg _407209_407209 ; 
   reg __407209_407209;
   reg _407210_407210 ; 
   reg __407210_407210;
   reg _407211_407211 ; 
   reg __407211_407211;
   reg _407212_407212 ; 
   reg __407212_407212;
   reg _407213_407213 ; 
   reg __407213_407213;
   reg _407214_407214 ; 
   reg __407214_407214;
   reg _407215_407215 ; 
   reg __407215_407215;
   reg _407216_407216 ; 
   reg __407216_407216;
   reg _407217_407217 ; 
   reg __407217_407217;
   reg _407218_407218 ; 
   reg __407218_407218;
   reg _407219_407219 ; 
   reg __407219_407219;
   reg _407220_407220 ; 
   reg __407220_407220;
   reg _407221_407221 ; 
   reg __407221_407221;
   reg _407222_407222 ; 
   reg __407222_407222;
   reg _407223_407223 ; 
   reg __407223_407223;
   reg _407224_407224 ; 
   reg __407224_407224;
   reg _407225_407225 ; 
   reg __407225_407225;
   reg _407226_407226 ; 
   reg __407226_407226;
   reg _407227_407227 ; 
   reg __407227_407227;
   reg _407228_407228 ; 
   reg __407228_407228;
   reg _407229_407229 ; 
   reg __407229_407229;
   reg _407230_407230 ; 
   reg __407230_407230;
   reg _407231_407231 ; 
   reg __407231_407231;
   reg _407232_407232 ; 
   reg __407232_407232;
   reg _407233_407233 ; 
   reg __407233_407233;
   reg _407234_407234 ; 
   reg __407234_407234;
   reg _407235_407235 ; 
   reg __407235_407235;
   reg _407236_407236 ; 
   reg __407236_407236;
   reg _407237_407237 ; 
   reg __407237_407237;
   reg _407238_407238 ; 
   reg __407238_407238;
   reg _407239_407239 ; 
   reg __407239_407239;
   reg _407240_407240 ; 
   reg __407240_407240;
   reg _407241_407241 ; 
   reg __407241_407241;
   reg _407242_407242 ; 
   reg __407242_407242;
   reg _407243_407243 ; 
   reg __407243_407243;
   reg _407244_407244 ; 
   reg __407244_407244;
   reg _407245_407245 ; 
   reg __407245_407245;
   reg _407246_407246 ; 
   reg __407246_407246;
   reg _407247_407247 ; 
   reg __407247_407247;
   reg _407248_407248 ; 
   reg __407248_407248;
   reg _407249_407249 ; 
   reg __407249_407249;
   reg _407250_407250 ; 
   reg __407250_407250;
   reg _407251_407251 ; 
   reg __407251_407251;
   reg _407252_407252 ; 
   reg __407252_407252;
   reg _407253_407253 ; 
   reg __407253_407253;
   reg _407254_407254 ; 
   reg __407254_407254;
   reg _407255_407255 ; 
   reg __407255_407255;
   reg _407256_407256 ; 
   reg __407256_407256;
   reg _407257_407257 ; 
   reg __407257_407257;
   reg _407258_407258 ; 
   reg __407258_407258;
   reg _407259_407259 ; 
   reg __407259_407259;
   reg _407260_407260 ; 
   reg __407260_407260;
   reg _407261_407261 ; 
   reg __407261_407261;
   reg _407262_407262 ; 
   reg __407262_407262;
   reg _407263_407263 ; 
   reg __407263_407263;
   reg _407264_407264 ; 
   reg __407264_407264;
   reg _407265_407265 ; 
   reg __407265_407265;
   reg _407266_407266 ; 
   reg __407266_407266;
   reg _407267_407267 ; 
   reg __407267_407267;
   reg _407268_407268 ; 
   reg __407268_407268;
   reg _407269_407269 ; 
   reg __407269_407269;
   reg _407270_407270 ; 
   reg __407270_407270;
   reg _407271_407271 ; 
   reg __407271_407271;
   reg _407272_407272 ; 
   reg __407272_407272;
   reg _407273_407273 ; 
   reg __407273_407273;
   reg _407274_407274 ; 
   reg __407274_407274;
   reg _407275_407275 ; 
   reg __407275_407275;
   reg _407276_407276 ; 
   reg __407276_407276;
   reg _407277_407277 ; 
   reg __407277_407277;
   reg _407278_407278 ; 
   reg __407278_407278;
   reg _407279_407279 ; 
   reg __407279_407279;
   reg _407280_407280 ; 
   reg __407280_407280;
   reg _407281_407281 ; 
   reg __407281_407281;
   reg _407282_407282 ; 
   reg __407282_407282;
   reg _407283_407283 ; 
   reg __407283_407283;
   reg _407284_407284 ; 
   reg __407284_407284;
   reg _407285_407285 ; 
   reg __407285_407285;
   reg _407286_407286 ; 
   reg __407286_407286;
   reg _407287_407287 ; 
   reg __407287_407287;
   reg _407288_407288 ; 
   reg __407288_407288;
   reg _407289_407289 ; 
   reg __407289_407289;
   reg _407290_407290 ; 
   reg __407290_407290;
   reg _407291_407291 ; 
   reg __407291_407291;
   reg _407292_407292 ; 
   reg __407292_407292;
   reg _407293_407293 ; 
   reg __407293_407293;
   reg _407294_407294 ; 
   reg __407294_407294;
   reg _407295_407295 ; 
   reg __407295_407295;
   reg _407296_407296 ; 
   reg __407296_407296;
   reg _407297_407297 ; 
   reg __407297_407297;
   reg _407298_407298 ; 
   reg __407298_407298;
   reg _407299_407299 ; 
   reg __407299_407299;
   reg _407300_407300 ; 
   reg __407300_407300;
   reg _407301_407301 ; 
   reg __407301_407301;
   reg _407302_407302 ; 
   reg __407302_407302;
   reg _407303_407303 ; 
   reg __407303_407303;
   reg _407304_407304 ; 
   reg __407304_407304;
   reg _407305_407305 ; 
   reg __407305_407305;
   reg _407306_407306 ; 
   reg __407306_407306;
   reg _407307_407307 ; 
   reg __407307_407307;
   reg _407308_407308 ; 
   reg __407308_407308;
   reg _407309_407309 ; 
   reg __407309_407309;
   reg _407310_407310 ; 
   reg __407310_407310;
   reg _407311_407311 ; 
   reg __407311_407311;
   reg _407312_407312 ; 
   reg __407312_407312;
   reg _407313_407313 ; 
   reg __407313_407313;
   reg _407314_407314 ; 
   reg __407314_407314;
   reg _407315_407315 ; 
   reg __407315_407315;
   reg _407316_407316 ; 
   reg __407316_407316;
   reg _407317_407317 ; 
   reg __407317_407317;
   reg _407318_407318 ; 
   reg __407318_407318;
   reg _407319_407319 ; 
   reg __407319_407319;
   reg _407320_407320 ; 
   reg __407320_407320;
   reg _407321_407321 ; 
   reg __407321_407321;
   reg _407322_407322 ; 
   reg __407322_407322;
   reg _407323_407323 ; 
   reg __407323_407323;
   reg _407324_407324 ; 
   reg __407324_407324;
   reg _407325_407325 ; 
   reg __407325_407325;
   reg _407326_407326 ; 
   reg __407326_407326;
   reg _407327_407327 ; 
   reg __407327_407327;
   reg _407328_407328 ; 
   reg __407328_407328;
   reg _407329_407329 ; 
   reg __407329_407329;
   reg _407330_407330 ; 
   reg __407330_407330;
   reg _407331_407331 ; 
   reg __407331_407331;
   reg _407332_407332 ; 
   reg __407332_407332;
   reg _407333_407333 ; 
   reg __407333_407333;
   reg _407334_407334 ; 
   reg __407334_407334;
   reg _407335_407335 ; 
   reg __407335_407335;
   reg _407336_407336 ; 
   reg __407336_407336;
   reg _407337_407337 ; 
   reg __407337_407337;
   reg _407338_407338 ; 
   reg __407338_407338;
   reg _407339_407339 ; 
   reg __407339_407339;
   reg _407340_407340 ; 
   reg __407340_407340;
   reg _407341_407341 ; 
   reg __407341_407341;
   reg _407342_407342 ; 
   reg __407342_407342;
   reg _407343_407343 ; 
   reg __407343_407343;
   reg _407344_407344 ; 
   reg __407344_407344;
   reg _407345_407345 ; 
   reg __407345_407345;
   reg _407346_407346 ; 
   reg __407346_407346;
   reg _407347_407347 ; 
   reg __407347_407347;
   reg _407348_407348 ; 
   reg __407348_407348;
   reg _407349_407349 ; 
   reg __407349_407349;
   reg _407350_407350 ; 
   reg __407350_407350;
   reg _407351_407351 ; 
   reg __407351_407351;
   reg _407352_407352 ; 
   reg __407352_407352;
   reg _407353_407353 ; 
   reg __407353_407353;
   reg _407354_407354 ; 
   reg __407354_407354;
   reg _407355_407355 ; 
   reg __407355_407355;
   reg _407356_407356 ; 
   reg __407356_407356;
   reg _407357_407357 ; 
   reg __407357_407357;
   reg _407358_407358 ; 
   reg __407358_407358;
   reg _407359_407359 ; 
   reg __407359_407359;
   reg _407360_407360 ; 
   reg __407360_407360;
   reg _407361_407361 ; 
   reg __407361_407361;
   reg _407362_407362 ; 
   reg __407362_407362;
   reg _407363_407363 ; 
   reg __407363_407363;
   reg _407364_407364 ; 
   reg __407364_407364;
   reg _407365_407365 ; 
   reg __407365_407365;
   reg _407366_407366 ; 
   reg __407366_407366;
   reg _407367_407367 ; 
   reg __407367_407367;
   reg _407368_407368 ; 
   reg __407368_407368;
   reg _407369_407369 ; 
   reg __407369_407369;
   reg _407370_407370 ; 
   reg __407370_407370;
   reg _407371_407371 ; 
   reg __407371_407371;
   reg _407372_407372 ; 
   reg __407372_407372;
   reg _407373_407373 ; 
   reg __407373_407373;
   reg _407374_407374 ; 
   reg __407374_407374;
   reg _407375_407375 ; 
   reg __407375_407375;
   reg _407376_407376 ; 
   reg __407376_407376;
   reg _407377_407377 ; 
   reg __407377_407377;
   reg _407378_407378 ; 
   reg __407378_407378;
   reg _407379_407379 ; 
   reg __407379_407379;
   reg _407380_407380 ; 
   reg __407380_407380;
   reg _407381_407381 ; 
   reg __407381_407381;
   reg _407382_407382 ; 
   reg __407382_407382;
   reg _407383_407383 ; 
   reg __407383_407383;
   reg _407384_407384 ; 
   reg __407384_407384;
   reg _407385_407385 ; 
   reg __407385_407385;
   reg _407386_407386 ; 
   reg __407386_407386;
   reg _407387_407387 ; 
   reg __407387_407387;
   reg _407388_407388 ; 
   reg __407388_407388;
   reg _407389_407389 ; 
   reg __407389_407389;
   reg _407390_407390 ; 
   reg __407390_407390;
   reg _407391_407391 ; 
   reg __407391_407391;
   reg _407392_407392 ; 
   reg __407392_407392;
   reg _407393_407393 ; 
   reg __407393_407393;
   reg _407394_407394 ; 
   reg __407394_407394;
   reg _407395_407395 ; 
   reg __407395_407395;
   reg _407396_407396 ; 
   reg __407396_407396;
   reg _407397_407397 ; 
   reg __407397_407397;
   reg _407398_407398 ; 
   reg __407398_407398;
   reg _407399_407399 ; 
   reg __407399_407399;
   reg _407400_407400 ; 
   reg __407400_407400;
   reg _407401_407401 ; 
   reg __407401_407401;
   reg _407402_407402 ; 
   reg __407402_407402;
   reg _407403_407403 ; 
   reg __407403_407403;
   reg _407404_407404 ; 
   reg __407404_407404;
   reg _407405_407405 ; 
   reg __407405_407405;
   reg _407406_407406 ; 
   reg __407406_407406;
   reg _407407_407407 ; 
   reg __407407_407407;
   reg _407408_407408 ; 
   reg __407408_407408;
   reg _407409_407409 ; 
   reg __407409_407409;
   reg _407410_407410 ; 
   reg __407410_407410;
   reg _407411_407411 ; 
   reg __407411_407411;
   reg _407412_407412 ; 
   reg __407412_407412;
   reg _407413_407413 ; 
   reg __407413_407413;
   reg _407414_407414 ; 
   reg __407414_407414;
   reg _407415_407415 ; 
   reg __407415_407415;
   reg _407416_407416 ; 
   reg __407416_407416;
   reg _407417_407417 ; 
   reg __407417_407417;
   reg _407418_407418 ; 
   reg __407418_407418;
   reg _407419_407419 ; 
   reg __407419_407419;
   reg _407420_407420 ; 
   reg __407420_407420;
   reg _407421_407421 ; 
   reg __407421_407421;
   reg _407422_407422 ; 
   reg __407422_407422;
   reg _407423_407423 ; 
   reg __407423_407423;
   reg _407424_407424 ; 
   reg __407424_407424;
   reg _407425_407425 ; 
   reg __407425_407425;
   reg _407426_407426 ; 
   reg __407426_407426;
   reg _407427_407427 ; 
   reg __407427_407427;
   reg _407428_407428 ; 
   reg __407428_407428;
   reg _407429_407429 ; 
   reg __407429_407429;
   reg _407430_407430 ; 
   reg __407430_407430;
   reg _407431_407431 ; 
   reg __407431_407431;
   reg _407432_407432 ; 
   reg __407432_407432;
   reg _407433_407433 ; 
   reg __407433_407433;
   reg _407434_407434 ; 
   reg __407434_407434;
   reg _407435_407435 ; 
   reg __407435_407435;
   reg _407436_407436 ; 
   reg __407436_407436;
   reg _407437_407437 ; 
   reg __407437_407437;
   reg _407438_407438 ; 
   reg __407438_407438;
   reg _407439_407439 ; 
   reg __407439_407439;
   reg _407440_407440 ; 
   reg __407440_407440;
   reg _407441_407441 ; 
   reg __407441_407441;
   reg _407442_407442 ; 
   reg __407442_407442;
   reg _407443_407443 ; 
   reg __407443_407443;
   reg _407444_407444 ; 
   reg __407444_407444;
   reg _407445_407445 ; 
   reg __407445_407445;
   reg _407446_407446 ; 
   reg __407446_407446;
   reg _407447_407447 ; 
   reg __407447_407447;
   reg _407448_407448 ; 
   reg __407448_407448;
   reg _407449_407449 ; 
   reg __407449_407449;
   reg _407450_407450 ; 
   reg __407450_407450;
   reg _407451_407451 ; 
   reg __407451_407451;
   reg _407452_407452 ; 
   reg __407452_407452;
   reg _407453_407453 ; 
   reg __407453_407453;
   reg _407454_407454 ; 
   reg __407454_407454;
   reg _407455_407455 ; 
   reg __407455_407455;
   reg _407456_407456 ; 
   reg __407456_407456;
   reg _407457_407457 ; 
   reg __407457_407457;
   reg _407458_407458 ; 
   reg __407458_407458;
   reg _407459_407459 ; 
   reg __407459_407459;
   reg _407460_407460 ; 
   reg __407460_407460;
   reg _407461_407461 ; 
   reg __407461_407461;
   reg _407462_407462 ; 
   reg __407462_407462;
   reg _407463_407463 ; 
   reg __407463_407463;
   reg _407464_407464 ; 
   reg __407464_407464;
   reg _407465_407465 ; 
   reg __407465_407465;
   reg _407466_407466 ; 
   reg __407466_407466;
   reg _407467_407467 ; 
   reg __407467_407467;
   reg _407468_407468 ; 
   reg __407468_407468;
   reg _407469_407469 ; 
   reg __407469_407469;
   reg _407470_407470 ; 
   reg __407470_407470;
   reg _407471_407471 ; 
   reg __407471_407471;
   reg _407472_407472 ; 
   reg __407472_407472;
   reg _407473_407473 ; 
   reg __407473_407473;
   reg _407474_407474 ; 
   reg __407474_407474;
   reg _407475_407475 ; 
   reg __407475_407475;
   reg _407476_407476 ; 
   reg __407476_407476;
   reg _407477_407477 ; 
   reg __407477_407477;
   reg _407478_407478 ; 
   reg __407478_407478;
   reg _407479_407479 ; 
   reg __407479_407479;
   reg _407480_407480 ; 
   reg __407480_407480;
   reg _407481_407481 ; 
   reg __407481_407481;
   reg _407482_407482 ; 
   reg __407482_407482;
   reg _407483_407483 ; 
   reg __407483_407483;
   reg _407484_407484 ; 
   reg __407484_407484;
   reg _407485_407485 ; 
   reg __407485_407485;
   reg _407486_407486 ; 
   reg __407486_407486;
   reg _407487_407487 ; 
   reg __407487_407487;
   reg _407488_407488 ; 
   reg __407488_407488;
   reg _407489_407489 ; 
   reg __407489_407489;
   reg _407490_407490 ; 
   reg __407490_407490;
   reg _407491_407491 ; 
   reg __407491_407491;
   reg _407492_407492 ; 
   reg __407492_407492;
   reg _407493_407493 ; 
   reg __407493_407493;
   reg _407494_407494 ; 
   reg __407494_407494;
   reg _407495_407495 ; 
   reg __407495_407495;
   reg _407496_407496 ; 
   reg __407496_407496;
   reg _407497_407497 ; 
   reg __407497_407497;
   reg _407498_407498 ; 
   reg __407498_407498;
   reg _407499_407499 ; 
   reg __407499_407499;
   reg _407500_407500 ; 
   reg __407500_407500;
   reg _407501_407501 ; 
   reg __407501_407501;
   reg _407502_407502 ; 
   reg __407502_407502;
   reg _407503_407503 ; 
   reg __407503_407503;
   reg _407504_407504 ; 
   reg __407504_407504;
   reg _407505_407505 ; 
   reg __407505_407505;
   reg _407506_407506 ; 
   reg __407506_407506;
   reg _407507_407507 ; 
   reg __407507_407507;
   reg _407508_407508 ; 
   reg __407508_407508;
   reg _407509_407509 ; 
   reg __407509_407509;
   reg _407510_407510 ; 
   reg __407510_407510;
   reg _407511_407511 ; 
   reg __407511_407511;
   reg _407512_407512 ; 
   reg __407512_407512;
   reg _407513_407513 ; 
   reg __407513_407513;
   reg _407514_407514 ; 
   reg __407514_407514;
   reg _407515_407515 ; 
   reg __407515_407515;
   reg _407516_407516 ; 
   reg __407516_407516;
   reg _407517_407517 ; 
   reg __407517_407517;
   reg _407518_407518 ; 
   reg __407518_407518;
   reg _407519_407519 ; 
   reg __407519_407519;
   reg _407520_407520 ; 
   reg __407520_407520;
   reg _407521_407521 ; 
   reg __407521_407521;
   reg _407522_407522 ; 
   reg __407522_407522;
   reg _407523_407523 ; 
   reg __407523_407523;
   reg _407524_407524 ; 
   reg __407524_407524;
   reg _407525_407525 ; 
   reg __407525_407525;
   reg _407526_407526 ; 
   reg __407526_407526;
   reg _407527_407527 ; 
   reg __407527_407527;
   reg _407528_407528 ; 
   reg __407528_407528;
   reg _407529_407529 ; 
   reg __407529_407529;
   reg _407530_407530 ; 
   reg __407530_407530;
   reg _407531_407531 ; 
   reg __407531_407531;
   reg _407532_407532 ; 
   reg __407532_407532;
   reg _407533_407533 ; 
   reg __407533_407533;
   reg _407534_407534 ; 
   reg __407534_407534;
   reg _407535_407535 ; 
   reg __407535_407535;
   reg _407536_407536 ; 
   reg __407536_407536;
   reg _407537_407537 ; 
   reg __407537_407537;
   reg _407538_407538 ; 
   reg __407538_407538;
   reg _407539_407539 ; 
   reg __407539_407539;
   reg _407540_407540 ; 
   reg __407540_407540;
   reg _407541_407541 ; 
   reg __407541_407541;
   reg _407542_407542 ; 
   reg __407542_407542;
   reg _407543_407543 ; 
   reg __407543_407543;
   reg _407544_407544 ; 
   reg __407544_407544;
   reg _407545_407545 ; 
   reg __407545_407545;
   reg _407546_407546 ; 
   reg __407546_407546;
   reg _407547_407547 ; 
   reg __407547_407547;
   reg _407548_407548 ; 
   reg __407548_407548;
   reg _407549_407549 ; 
   reg __407549_407549;
   reg _407550_407550 ; 
   reg __407550_407550;
   reg _407551_407551 ; 
   reg __407551_407551;
   reg _407552_407552 ; 
   reg __407552_407552;
   reg _407553_407553 ; 
   reg __407553_407553;
   reg _407554_407554 ; 
   reg __407554_407554;
   reg _407555_407555 ; 
   reg __407555_407555;
   reg _407556_407556 ; 
   reg __407556_407556;
   reg _407557_407557 ; 
   reg __407557_407557;
   reg _407558_407558 ; 
   reg __407558_407558;
   reg _407559_407559 ; 
   reg __407559_407559;
   reg _407560_407560 ; 
   reg __407560_407560;
   reg _407561_407561 ; 
   reg __407561_407561;
   reg _407562_407562 ; 
   reg __407562_407562;
   reg _407563_407563 ; 
   reg __407563_407563;
   reg _407564_407564 ; 
   reg __407564_407564;
   reg _407565_407565 ; 
   reg __407565_407565;
   reg _407566_407566 ; 
   reg __407566_407566;
   reg _407567_407567 ; 
   reg __407567_407567;
   reg _407568_407568 ; 
   reg __407568_407568;
   reg _407569_407569 ; 
   reg __407569_407569;
   reg _407570_407570 ; 
   reg __407570_407570;
   reg _407571_407571 ; 
   reg __407571_407571;
   reg _407572_407572 ; 
   reg __407572_407572;
   reg _407573_407573 ; 
   reg __407573_407573;
   reg _407574_407574 ; 
   reg __407574_407574;
   reg _407575_407575 ; 
   reg __407575_407575;
   reg _407576_407576 ; 
   reg __407576_407576;
   reg _407577_407577 ; 
   reg __407577_407577;
   reg _407578_407578 ; 
   reg __407578_407578;
   reg _407579_407579 ; 
   reg __407579_407579;
   reg _407580_407580 ; 
   reg __407580_407580;
   reg _407581_407581 ; 
   reg __407581_407581;
   reg _407582_407582 ; 
   reg __407582_407582;
   reg _407583_407583 ; 
   reg __407583_407583;
   reg _407584_407584 ; 
   reg __407584_407584;
   reg _407585_407585 ; 
   reg __407585_407585;
   reg _407586_407586 ; 
   reg __407586_407586;
   reg _407587_407587 ; 
   reg __407587_407587;
   reg _407588_407588 ; 
   reg __407588_407588;
   reg _407589_407589 ; 
   reg __407589_407589;
   reg _407590_407590 ; 
   reg __407590_407590;
   reg _407591_407591 ; 
   reg __407591_407591;
   reg _407592_407592 ; 
   reg __407592_407592;
   reg _407593_407593 ; 
   reg __407593_407593;
   reg _407594_407594 ; 
   reg __407594_407594;
   reg _407595_407595 ; 
   reg __407595_407595;
   reg _407596_407596 ; 
   reg __407596_407596;
   reg _407597_407597 ; 
   reg __407597_407597;
   reg _407598_407598 ; 
   reg __407598_407598;
   reg _407599_407599 ; 
   reg __407599_407599;
   reg _407600_407600 ; 
   reg __407600_407600;
   reg _407601_407601 ; 
   reg __407601_407601;
   reg _407602_407602 ; 
   reg __407602_407602;
   reg _407603_407603 ; 
   reg __407603_407603;
   reg _407604_407604 ; 
   reg __407604_407604;
   reg _407605_407605 ; 
   reg __407605_407605;
   reg _407606_407606 ; 
   reg __407606_407606;
   reg _407607_407607 ; 
   reg __407607_407607;
   reg _407608_407608 ; 
   reg __407608_407608;
   reg _407609_407609 ; 
   reg __407609_407609;
   reg _407610_407610 ; 
   reg __407610_407610;
   reg _407611_407611 ; 
   reg __407611_407611;
   reg _407612_407612 ; 
   reg __407612_407612;
   reg _407613_407613 ; 
   reg __407613_407613;
   reg _407614_407614 ; 
   reg __407614_407614;
   reg _407615_407615 ; 
   reg __407615_407615;
   reg _407616_407616 ; 
   reg __407616_407616;
   reg _407617_407617 ; 
   reg __407617_407617;
   reg _407618_407618 ; 
   reg __407618_407618;
   reg _407619_407619 ; 
   reg __407619_407619;
   reg _407620_407620 ; 
   reg __407620_407620;
   reg _407621_407621 ; 
   reg __407621_407621;
   reg _407622_407622 ; 
   reg __407622_407622;
   reg _407623_407623 ; 
   reg __407623_407623;
   reg _407624_407624 ; 
   reg __407624_407624;
   reg _407625_407625 ; 
   reg __407625_407625;
   reg _407626_407626 ; 
   reg __407626_407626;
   reg _407627_407627 ; 
   reg __407627_407627;
   reg _407628_407628 ; 
   reg __407628_407628;
   reg _407629_407629 ; 
   reg __407629_407629;
   reg _407630_407630 ; 
   reg __407630_407630;
   reg _407631_407631 ; 
   reg __407631_407631;
   reg _407632_407632 ; 
   reg __407632_407632;
   reg _407633_407633 ; 
   reg __407633_407633;
   reg _407634_407634 ; 
   reg __407634_407634;
   reg _407635_407635 ; 
   reg __407635_407635;
   reg _407636_407636 ; 
   reg __407636_407636;
   reg _407637_407637 ; 
   reg __407637_407637;
   reg _407638_407638 ; 
   reg __407638_407638;
   reg _407639_407639 ; 
   reg __407639_407639;
   reg _407640_407640 ; 
   reg __407640_407640;
   reg _407641_407641 ; 
   reg __407641_407641;
   reg _407642_407642 ; 
   reg __407642_407642;
   reg _407643_407643 ; 
   reg __407643_407643;
   reg _407644_407644 ; 
   reg __407644_407644;
   reg _407645_407645 ; 
   reg __407645_407645;
   reg _407646_407646 ; 
   reg __407646_407646;
   reg _407647_407647 ; 
   reg __407647_407647;
   reg _407648_407648 ; 
   reg __407648_407648;
   reg _407649_407649 ; 
   reg __407649_407649;
   reg _407650_407650 ; 
   reg __407650_407650;
   reg _407651_407651 ; 
   reg __407651_407651;
   reg _407652_407652 ; 
   reg __407652_407652;
   reg _407653_407653 ; 
   reg __407653_407653;
   reg _407654_407654 ; 
   reg __407654_407654;
   reg _407655_407655 ; 
   reg __407655_407655;
   reg _407656_407656 ; 
   reg __407656_407656;
   reg _407657_407657 ; 
   reg __407657_407657;
   reg _407658_407658 ; 
   reg __407658_407658;
   reg _407659_407659 ; 
   reg __407659_407659;
   reg _407660_407660 ; 
   reg __407660_407660;
   reg _407661_407661 ; 
   reg __407661_407661;
   reg _407662_407662 ; 
   reg __407662_407662;
   reg _407663_407663 ; 
   reg __407663_407663;
   reg _407664_407664 ; 
   reg __407664_407664;
   reg _407665_407665 ; 
   reg __407665_407665;
   reg _407666_407666 ; 
   reg __407666_407666;
   reg _407667_407667 ; 
   reg __407667_407667;
   reg _407668_407668 ; 
   reg __407668_407668;
   reg _407669_407669 ; 
   reg __407669_407669;
   reg _407670_407670 ; 
   reg __407670_407670;
   reg _407671_407671 ; 
   reg __407671_407671;
   reg _407672_407672 ; 
   reg __407672_407672;
   reg _407673_407673 ; 
   reg __407673_407673;
   reg _407674_407674 ; 
   reg __407674_407674;
   reg _407675_407675 ; 
   reg __407675_407675;
   reg _407676_407676 ; 
   reg __407676_407676;
   reg _407677_407677 ; 
   reg __407677_407677;
   reg _407678_407678 ; 
   reg __407678_407678;
   reg _407679_407679 ; 
   reg __407679_407679;
   reg _407680_407680 ; 
   reg __407680_407680;
   reg _407681_407681 ; 
   reg __407681_407681;
   reg _407682_407682 ; 
   reg __407682_407682;
   reg _407683_407683 ; 
   reg __407683_407683;
   reg _407684_407684 ; 
   reg __407684_407684;
   reg _407685_407685 ; 
   reg __407685_407685;
   reg _407686_407686 ; 
   reg __407686_407686;
   reg _407687_407687 ; 
   reg __407687_407687;
   reg _407688_407688 ; 
   reg __407688_407688;
   reg _407689_407689 ; 
   reg __407689_407689;
   reg _407690_407690 ; 
   reg __407690_407690;
   reg _407691_407691 ; 
   reg __407691_407691;
   reg _407692_407692 ; 
   reg __407692_407692;
   reg _407693_407693 ; 
   reg __407693_407693;
   reg _407694_407694 ; 
   reg __407694_407694;
   reg _407695_407695 ; 
   reg __407695_407695;
   reg _407696_407696 ; 
   reg __407696_407696;
   reg _407697_407697 ; 
   reg __407697_407697;
   reg _407698_407698 ; 
   reg __407698_407698;
   reg _407699_407699 ; 
   reg __407699_407699;
   reg _407700_407700 ; 
   reg __407700_407700;
   reg _407701_407701 ; 
   reg __407701_407701;
   reg _407702_407702 ; 
   reg __407702_407702;
   reg _407703_407703 ; 
   reg __407703_407703;
   reg _407704_407704 ; 
   reg __407704_407704;
   reg _407705_407705 ; 
   reg __407705_407705;
   reg _407706_407706 ; 
   reg __407706_407706;
   reg _407707_407707 ; 
   reg __407707_407707;
   reg _407708_407708 ; 
   reg __407708_407708;
   reg _407709_407709 ; 
   reg __407709_407709;
   reg _407710_407710 ; 
   reg __407710_407710;
   reg _407711_407711 ; 
   reg __407711_407711;
   reg _407712_407712 ; 
   reg __407712_407712;
   reg _407713_407713 ; 
   reg __407713_407713;
   reg _407714_407714 ; 
   reg __407714_407714;
   reg _407715_407715 ; 
   reg __407715_407715;
   reg _407716_407716 ; 
   reg __407716_407716;
   reg _407717_407717 ; 
   reg __407717_407717;
   reg _407718_407718 ; 
   reg __407718_407718;
   reg _407719_407719 ; 
   reg __407719_407719;
   reg _407720_407720 ; 
   reg __407720_407720;
   reg _407721_407721 ; 
   reg __407721_407721;
   reg _407722_407722 ; 
   reg __407722_407722;
   reg _407723_407723 ; 
   reg __407723_407723;
   reg _407724_407724 ; 
   reg __407724_407724;
   reg _407725_407725 ; 
   reg __407725_407725;
   reg _407726_407726 ; 
   reg __407726_407726;
   reg _407727_407727 ; 
   reg __407727_407727;
   reg _407728_407728 ; 
   reg __407728_407728;
   reg _407729_407729 ; 
   reg __407729_407729;
   reg _407730_407730 ; 
   reg __407730_407730;
   reg _407731_407731 ; 
   reg __407731_407731;
   reg _407732_407732 ; 
   reg __407732_407732;
   reg _407733_407733 ; 
   reg __407733_407733;
   reg _407734_407734 ; 
   reg __407734_407734;
   reg _407735_407735 ; 
   reg __407735_407735;
   reg _407736_407736 ; 
   reg __407736_407736;
   reg _407737_407737 ; 
   reg __407737_407737;
   reg _407738_407738 ; 
   reg __407738_407738;
   reg _407739_407739 ; 
   reg __407739_407739;
   reg _407740_407740 ; 
   reg __407740_407740;
   reg _407741_407741 ; 
   reg __407741_407741;
   reg _407742_407742 ; 
   reg __407742_407742;
   reg _407743_407743 ; 
   reg __407743_407743;
   reg _407744_407744 ; 
   reg __407744_407744;
   reg _407745_407745 ; 
   reg __407745_407745;
   reg _407746_407746 ; 
   reg __407746_407746;
   reg _407747_407747 ; 
   reg __407747_407747;
   reg _407748_407748 ; 
   reg __407748_407748;
   reg _407749_407749 ; 
   reg __407749_407749;
   reg _407750_407750 ; 
   reg __407750_407750;
   reg _407751_407751 ; 
   reg __407751_407751;
   reg _407752_407752 ; 
   reg __407752_407752;
   reg _407753_407753 ; 
   reg __407753_407753;
   reg _407754_407754 ; 
   reg __407754_407754;
   reg _407755_407755 ; 
   reg __407755_407755;
   reg _407756_407756 ; 
   reg __407756_407756;
   reg _407757_407757 ; 
   reg __407757_407757;
   reg _407758_407758 ; 
   reg __407758_407758;
   reg _407759_407759 ; 
   reg __407759_407759;
   reg _407760_407760 ; 
   reg __407760_407760;
   reg _407761_407761 ; 
   reg __407761_407761;
   reg _407762_407762 ; 
   reg __407762_407762;
   reg _407763_407763 ; 
   reg __407763_407763;
   reg _407764_407764 ; 
   reg __407764_407764;
   reg _407765_407765 ; 
   reg __407765_407765;
   reg _407766_407766 ; 
   reg __407766_407766;
   reg _407767_407767 ; 
   reg __407767_407767;
   reg _407768_407768 ; 
   reg __407768_407768;
   reg _407769_407769 ; 
   reg __407769_407769;
   reg _407770_407770 ; 
   reg __407770_407770;
   reg _407771_407771 ; 
   reg __407771_407771;
   reg _407772_407772 ; 
   reg __407772_407772;
   reg _407773_407773 ; 
   reg __407773_407773;
   reg _407774_407774 ; 
   reg __407774_407774;
   reg _407775_407775 ; 
   reg __407775_407775;
   reg _407776_407776 ; 
   reg __407776_407776;
   reg _407777_407777 ; 
   reg __407777_407777;
   reg _407778_407778 ; 
   reg __407778_407778;
   reg _407779_407779 ; 
   reg __407779_407779;
   reg _407780_407780 ; 
   reg __407780_407780;
   reg _407781_407781 ; 
   reg __407781_407781;
   reg _407782_407782 ; 
   reg __407782_407782;
   reg _407783_407783 ; 
   reg __407783_407783;
   reg _407784_407784 ; 
   reg __407784_407784;
   reg _407785_407785 ; 
   reg __407785_407785;
   reg _407786_407786 ; 
   reg __407786_407786;
   reg _407787_407787 ; 
   reg __407787_407787;
   reg _407788_407788 ; 
   reg __407788_407788;
   reg _407789_407789 ; 
   reg __407789_407789;
   reg _407790_407790 ; 
   reg __407790_407790;
   reg _407791_407791 ; 
   reg __407791_407791;
   reg _407792_407792 ; 
   reg __407792_407792;
   reg _407793_407793 ; 
   reg __407793_407793;
   reg _407794_407794 ; 
   reg __407794_407794;
   reg _407795_407795 ; 
   reg __407795_407795;
   reg _407796_407796 ; 
   reg __407796_407796;
   reg _407797_407797 ; 
   reg __407797_407797;
   reg _407798_407798 ; 
   reg __407798_407798;
   reg _407799_407799 ; 
   reg __407799_407799;
   reg _407800_407800 ; 
   reg __407800_407800;
   reg _407801_407801 ; 
   reg __407801_407801;
   reg _407802_407802 ; 
   reg __407802_407802;
   reg _407803_407803 ; 
   reg __407803_407803;
   reg _407804_407804 ; 
   reg __407804_407804;
   reg _407805_407805 ; 
   reg __407805_407805;
   reg _407806_407806 ; 
   reg __407806_407806;
   reg _407807_407807 ; 
   reg __407807_407807;
   reg _407808_407808 ; 
   reg __407808_407808;
   reg _407809_407809 ; 
   reg __407809_407809;
   reg _407810_407810 ; 
   reg __407810_407810;
   reg _407811_407811 ; 
   reg __407811_407811;
   reg _407812_407812 ; 
   reg __407812_407812;
   reg _407813_407813 ; 
   reg __407813_407813;
   reg _407814_407814 ; 
   reg __407814_407814;
   reg _407815_407815 ; 
   reg __407815_407815;
   reg _407816_407816 ; 
   reg __407816_407816;
   reg _407817_407817 ; 
   reg __407817_407817;
   reg _407818_407818 ; 
   reg __407818_407818;
   reg _407819_407819 ; 
   reg __407819_407819;
   reg _407820_407820 ; 
   reg __407820_407820;
   reg _407821_407821 ; 
   reg __407821_407821;
   reg _407822_407822 ; 
   reg __407822_407822;
   reg _407823_407823 ; 
   reg __407823_407823;
   reg _407824_407824 ; 
   reg __407824_407824;
   reg _407825_407825 ; 
   reg __407825_407825;
   reg _407826_407826 ; 
   reg __407826_407826;
   reg _407827_407827 ; 
   reg __407827_407827;
   reg _407828_407828 ; 
   reg __407828_407828;
   reg _407829_407829 ; 
   reg __407829_407829;
   reg _407830_407830 ; 
   reg __407830_407830;
   reg _407831_407831 ; 
   reg __407831_407831;
   reg _407832_407832 ; 
   reg __407832_407832;
   reg _407833_407833 ; 
   reg __407833_407833;
   reg _407834_407834 ; 
   reg __407834_407834;
   reg _407835_407835 ; 
   reg __407835_407835;
   reg _407836_407836 ; 
   reg __407836_407836;
   reg _407837_407837 ; 
   reg __407837_407837;
   reg _407838_407838 ; 
   reg __407838_407838;
   reg _407839_407839 ; 
   reg __407839_407839;
   reg _407840_407840 ; 
   reg __407840_407840;
   reg _407841_407841 ; 
   reg __407841_407841;
   reg _407842_407842 ; 
   reg __407842_407842;
   reg _407843_407843 ; 
   reg __407843_407843;
   reg _407844_407844 ; 
   reg __407844_407844;
   reg _407845_407845 ; 
   reg __407845_407845;
   reg _407846_407846 ; 
   reg __407846_407846;
   reg _407847_407847 ; 
   reg __407847_407847;
   reg _407848_407848 ; 
   reg __407848_407848;
   reg _407849_407849 ; 
   reg __407849_407849;
   reg _407850_407850 ; 
   reg __407850_407850;
   reg _407851_407851 ; 
   reg __407851_407851;
   reg _407852_407852 ; 
   reg __407852_407852;
   reg _407853_407853 ; 
   reg __407853_407853;
   reg _407854_407854 ; 
   reg __407854_407854;
   reg _407855_407855 ; 
   reg __407855_407855;
   reg _407856_407856 ; 
   reg __407856_407856;
   reg _407857_407857 ; 
   reg __407857_407857;
   reg _407858_407858 ; 
   reg __407858_407858;
   reg _407859_407859 ; 
   reg __407859_407859;
   reg _407860_407860 ; 
   reg __407860_407860;
   reg _407861_407861 ; 
   reg __407861_407861;
   reg _407862_407862 ; 
   reg __407862_407862;
   reg _407863_407863 ; 
   reg __407863_407863;
   reg _407864_407864 ; 
   reg __407864_407864;
   reg _407865_407865 ; 
   reg __407865_407865;
   reg _407866_407866 ; 
   reg __407866_407866;
   reg _407867_407867 ; 
   reg __407867_407867;
   reg _407868_407868 ; 
   reg __407868_407868;
   reg _407869_407869 ; 
   reg __407869_407869;
   reg _407870_407870 ; 
   reg __407870_407870;
   reg _407871_407871 ; 
   reg __407871_407871;
   reg _407872_407872 ; 
   reg __407872_407872;
   reg _407873_407873 ; 
   reg __407873_407873;
   reg _407874_407874 ; 
   reg __407874_407874;
   reg _407875_407875 ; 
   reg __407875_407875;
   reg _407876_407876 ; 
   reg __407876_407876;
   reg _407877_407877 ; 
   reg __407877_407877;
   reg _407878_407878 ; 
   reg __407878_407878;
   reg _407879_407879 ; 
   reg __407879_407879;
   reg _407880_407880 ; 
   reg __407880_407880;
   reg _407881_407881 ; 
   reg __407881_407881;
   reg _407882_407882 ; 
   reg __407882_407882;
   reg _407883_407883 ; 
   reg __407883_407883;
   reg _407884_407884 ; 
   reg __407884_407884;
   reg _407885_407885 ; 
   reg __407885_407885;
   reg _407886_407886 ; 
   reg __407886_407886;
   reg _407887_407887 ; 
   reg __407887_407887;
   reg _407888_407888 ; 
   reg __407888_407888;
   reg _407889_407889 ; 
   reg __407889_407889;
   reg _407890_407890 ; 
   reg __407890_407890;
   reg _407891_407891 ; 
   reg __407891_407891;
   reg _407892_407892 ; 
   reg __407892_407892;
   reg _407893_407893 ; 
   reg __407893_407893;
   reg _407894_407894 ; 
   reg __407894_407894;
   reg _407895_407895 ; 
   reg __407895_407895;
   reg _407896_407896 ; 
   reg __407896_407896;
   reg _407897_407897 ; 
   reg __407897_407897;
   reg _407898_407898 ; 
   reg __407898_407898;
   reg _407899_407899 ; 
   reg __407899_407899;
   reg _407900_407900 ; 
   reg __407900_407900;
   reg _407901_407901 ; 
   reg __407901_407901;
   reg _407902_407902 ; 
   reg __407902_407902;
   reg _407903_407903 ; 
   reg __407903_407903;
   reg _407904_407904 ; 
   reg __407904_407904;
   reg _407905_407905 ; 
   reg __407905_407905;
   reg _407906_407906 ; 
   reg __407906_407906;
   reg _407907_407907 ; 
   reg __407907_407907;
   reg _407908_407908 ; 
   reg __407908_407908;
   reg _407909_407909 ; 
   reg __407909_407909;
   reg _407910_407910 ; 
   reg __407910_407910;
   reg _407911_407911 ; 
   reg __407911_407911;
   reg _407912_407912 ; 
   reg __407912_407912;
   reg _407913_407913 ; 
   reg __407913_407913;
   reg _407914_407914 ; 
   reg __407914_407914;
   reg _407915_407915 ; 
   reg __407915_407915;
   reg _407916_407916 ; 
   reg __407916_407916;
   reg _407917_407917 ; 
   reg __407917_407917;
   reg _407918_407918 ; 
   reg __407918_407918;
   reg _407919_407919 ; 
   reg __407919_407919;
   reg _407920_407920 ; 
   reg __407920_407920;
   reg _407921_407921 ; 
   reg __407921_407921;
   reg _407922_407922 ; 
   reg __407922_407922;
   reg _407923_407923 ; 
   reg __407923_407923;
   reg _407924_407924 ; 
   reg __407924_407924;
   reg _407925_407925 ; 
   reg __407925_407925;
   reg _407926_407926 ; 
   reg __407926_407926;
   reg _407927_407927 ; 
   reg __407927_407927;
   reg _407928_407928 ; 
   reg __407928_407928;
   reg _407929_407929 ; 
   reg __407929_407929;
   reg _407930_407930 ; 
   reg __407930_407930;
   reg _407931_407931 ; 
   reg __407931_407931;
   reg _407932_407932 ; 
   reg __407932_407932;
   reg _407933_407933 ; 
   reg __407933_407933;
   reg _407934_407934 ; 
   reg __407934_407934;
   reg _407935_407935 ; 
   reg __407935_407935;
   reg _407936_407936 ; 
   reg __407936_407936;
   reg _407937_407937 ; 
   reg __407937_407937;
   reg _407938_407938 ; 
   reg __407938_407938;
   reg _407939_407939 ; 
   reg __407939_407939;
   reg _407940_407940 ; 
   reg __407940_407940;
   reg _407941_407941 ; 
   reg __407941_407941;
   reg _407942_407942 ; 
   reg __407942_407942;
   reg _407943_407943 ; 
   reg __407943_407943;
   reg _407944_407944 ; 
   reg __407944_407944;
   reg _407945_407945 ; 
   reg __407945_407945;
   reg _407946_407946 ; 
   reg __407946_407946;
   reg _407947_407947 ; 
   reg __407947_407947;
   reg _407948_407948 ; 
   reg __407948_407948;
   reg _407949_407949 ; 
   reg __407949_407949;
   reg _407950_407950 ; 
   reg __407950_407950;
   reg _407951_407951 ; 
   reg __407951_407951;
   reg _407952_407952 ; 
   reg __407952_407952;
   reg _407953_407953 ; 
   reg __407953_407953;
   reg _407954_407954 ; 
   reg __407954_407954;
   reg _407955_407955 ; 
   reg __407955_407955;
   reg _407956_407956 ; 
   reg __407956_407956;
   reg _407957_407957 ; 
   reg __407957_407957;
   reg _407958_407958 ; 
   reg __407958_407958;
   reg _407959_407959 ; 
   reg __407959_407959;
   reg _407960_407960 ; 
   reg __407960_407960;
   reg _407961_407961 ; 
   reg __407961_407961;
   reg _407962_407962 ; 
   reg __407962_407962;
   reg _407963_407963 ; 
   reg __407963_407963;
   reg _407964_407964 ; 
   reg __407964_407964;
   reg _407965_407965 ; 
   reg __407965_407965;
   reg _407966_407966 ; 
   reg __407966_407966;
   reg _407967_407967 ; 
   reg __407967_407967;
   reg _407968_407968 ; 
   reg __407968_407968;
   reg _407969_407969 ; 
   reg __407969_407969;
   reg _407970_407970 ; 
   reg __407970_407970;
   reg _407971_407971 ; 
   reg __407971_407971;
   reg _407972_407972 ; 
   reg __407972_407972;
   reg _407973_407973 ; 
   reg __407973_407973;
   reg _407974_407974 ; 
   reg __407974_407974;
   reg _407975_407975 ; 
   reg __407975_407975;
   reg _407976_407976 ; 
   reg __407976_407976;
   reg _407977_407977 ; 
   reg __407977_407977;
   reg _407978_407978 ; 
   reg __407978_407978;
   reg _407979_407979 ; 
   reg __407979_407979;
   reg _407980_407980 ; 
   reg __407980_407980;
   reg _407981_407981 ; 
   reg __407981_407981;
   reg _407982_407982 ; 
   reg __407982_407982;
   reg _407983_407983 ; 
   reg __407983_407983;
   reg _407984_407984 ; 
   reg __407984_407984;
   reg _407985_407985 ; 
   reg __407985_407985;
   reg _407986_407986 ; 
   reg __407986_407986;
   reg _407987_407987 ; 
   reg __407987_407987;
   reg _407988_407988 ; 
   reg __407988_407988;
   reg _407989_407989 ; 
   reg __407989_407989;
   reg _407990_407990 ; 
   reg __407990_407990;
   reg _407991_407991 ; 
   reg __407991_407991;
   reg _407992_407992 ; 
   reg __407992_407992;
   reg _407993_407993 ; 
   reg __407993_407993;
   reg _407994_407994 ; 
   reg __407994_407994;
   reg _407995_407995 ; 
   reg __407995_407995;
   reg _407996_407996 ; 
   reg __407996_407996;
   reg _407997_407997 ; 
   reg __407997_407997;
   reg _407998_407998 ; 
   reg __407998_407998;
   reg _407999_407999 ; 
   reg __407999_407999;
   reg _408000_408000 ; 
   reg __408000_408000;
   reg _408001_408001 ; 
   reg __408001_408001;
   reg _408002_408002 ; 
   reg __408002_408002;
   reg _408003_408003 ; 
   reg __408003_408003;
   reg _408004_408004 ; 
   reg __408004_408004;
   reg _408005_408005 ; 
   reg __408005_408005;
   reg _408006_408006 ; 
   reg __408006_408006;
   reg _408007_408007 ; 
   reg __408007_408007;
   reg _408008_408008 ; 
   reg __408008_408008;
   reg _408009_408009 ; 
   reg __408009_408009;
   reg _408010_408010 ; 
   reg __408010_408010;
   reg _408011_408011 ; 
   reg __408011_408011;
   reg _408012_408012 ; 
   reg __408012_408012;
   reg _408013_408013 ; 
   reg __408013_408013;
   reg _408014_408014 ; 
   reg __408014_408014;
   reg _408015_408015 ; 
   reg __408015_408015;
   reg _408016_408016 ; 
   reg __408016_408016;
   reg _408017_408017 ; 
   reg __408017_408017;
   reg _408018_408018 ; 
   reg __408018_408018;
   reg _408019_408019 ; 
   reg __408019_408019;
   reg _408020_408020 ; 
   reg __408020_408020;
   reg _408021_408021 ; 
   reg __408021_408021;
   reg _408022_408022 ; 
   reg __408022_408022;
   reg _408023_408023 ; 
   reg __408023_408023;
   reg _408024_408024 ; 
   reg __408024_408024;
   reg _408025_408025 ; 
   reg __408025_408025;
   reg _408026_408026 ; 
   reg __408026_408026;
   reg _408027_408027 ; 
   reg __408027_408027;
   reg _408028_408028 ; 
   reg __408028_408028;
   reg _408029_408029 ; 
   reg __408029_408029;
   reg _408030_408030 ; 
   reg __408030_408030;
   reg _408031_408031 ; 
   reg __408031_408031;
   reg _408032_408032 ; 
   reg __408032_408032;
   reg _408033_408033 ; 
   reg __408033_408033;
   reg _408034_408034 ; 
   reg __408034_408034;
   reg _408035_408035 ; 
   reg __408035_408035;
   reg _408036_408036 ; 
   reg __408036_408036;
   reg _408037_408037 ; 
   reg __408037_408037;
   reg _408038_408038 ; 
   reg __408038_408038;
   reg _408039_408039 ; 
   reg __408039_408039;
   reg _408040_408040 ; 
   reg __408040_408040;
   reg _408041_408041 ; 
   reg __408041_408041;
   reg _408042_408042 ; 
   reg __408042_408042;
   reg _408043_408043 ; 
   reg __408043_408043;
   reg _408044_408044 ; 
   reg __408044_408044;
   reg _408045_408045 ; 
   reg __408045_408045;
   reg _408046_408046 ; 
   reg __408046_408046;
   reg _408047_408047 ; 
   reg __408047_408047;
   reg _408048_408048 ; 
   reg __408048_408048;
   reg _408049_408049 ; 
   reg __408049_408049;
   reg _408050_408050 ; 
   reg __408050_408050;
   reg _408051_408051 ; 
   reg __408051_408051;
   reg _408052_408052 ; 
   reg __408052_408052;
   reg _408053_408053 ; 
   reg __408053_408053;
   reg _408054_408054 ; 
   reg __408054_408054;
   reg _408055_408055 ; 
   reg __408055_408055;
   reg _408056_408056 ; 
   reg __408056_408056;
   reg _408057_408057 ; 
   reg __408057_408057;
   reg _408058_408058 ; 
   reg __408058_408058;
   reg _408059_408059 ; 
   reg __408059_408059;
   reg _408060_408060 ; 
   reg __408060_408060;
   reg _408061_408061 ; 
   reg __408061_408061;
   reg _408062_408062 ; 
   reg __408062_408062;
   reg _408063_408063 ; 
   reg __408063_408063;
   reg _408064_408064 ; 
   reg __408064_408064;
   reg _408065_408065 ; 
   reg __408065_408065;
   reg _408066_408066 ; 
   reg __408066_408066;
   reg _408067_408067 ; 
   reg __408067_408067;
   reg _408068_408068 ; 
   reg __408068_408068;
   reg _408069_408069 ; 
   reg __408069_408069;
   reg _408070_408070 ; 
   reg __408070_408070;
   reg _408071_408071 ; 
   reg __408071_408071;
   reg _408072_408072 ; 
   reg __408072_408072;
   reg _408073_408073 ; 
   reg __408073_408073;
   reg _408074_408074 ; 
   reg __408074_408074;
   reg _408075_408075 ; 
   reg __408075_408075;
   reg _408076_408076 ; 
   reg __408076_408076;
   reg _408077_408077 ; 
   reg __408077_408077;
   reg _408078_408078 ; 
   reg __408078_408078;
   reg _408079_408079 ; 
   reg __408079_408079;
   reg _408080_408080 ; 
   reg __408080_408080;
   reg _408081_408081 ; 
   reg __408081_408081;
   reg _408082_408082 ; 
   reg __408082_408082;
   reg _408083_408083 ; 
   reg __408083_408083;
   reg _408084_408084 ; 
   reg __408084_408084;
   reg _408085_408085 ; 
   reg __408085_408085;
   reg _408086_408086 ; 
   reg __408086_408086;
   reg _408087_408087 ; 
   reg __408087_408087;
   reg _408088_408088 ; 
   reg __408088_408088;
   reg _408089_408089 ; 
   reg __408089_408089;
   reg _408090_408090 ; 
   reg __408090_408090;
   reg _408091_408091 ; 
   reg __408091_408091;
   reg _408092_408092 ; 
   reg __408092_408092;
   reg _408093_408093 ; 
   reg __408093_408093;
   reg _408094_408094 ; 
   reg __408094_408094;
   reg _408095_408095 ; 
   reg __408095_408095;
   reg _408096_408096 ; 
   reg __408096_408096;
   reg _408097_408097 ; 
   reg __408097_408097;
   reg _408098_408098 ; 
   reg __408098_408098;
   reg _408099_408099 ; 
   reg __408099_408099;
   reg _408100_408100 ; 
   reg __408100_408100;
   reg _408101_408101 ; 
   reg __408101_408101;
   reg _408102_408102 ; 
   reg __408102_408102;
   reg _408103_408103 ; 
   reg __408103_408103;
   reg _408104_408104 ; 
   reg __408104_408104;
   reg _408105_408105 ; 
   reg __408105_408105;
   reg _408106_408106 ; 
   reg __408106_408106;
   reg _408107_408107 ; 
   reg __408107_408107;
   reg _408108_408108 ; 
   reg __408108_408108;
   reg _408109_408109 ; 
   reg __408109_408109;
   reg _408110_408110 ; 
   reg __408110_408110;
   reg _408111_408111 ; 
   reg __408111_408111;
   reg _408112_408112 ; 
   reg __408112_408112;
   reg _408113_408113 ; 
   reg __408113_408113;
   reg _408114_408114 ; 
   reg __408114_408114;
   reg _408115_408115 ; 
   reg __408115_408115;
   reg _408116_408116 ; 
   reg __408116_408116;
   reg _408117_408117 ; 
   reg __408117_408117;
   reg _408118_408118 ; 
   reg __408118_408118;
   reg _408119_408119 ; 
   reg __408119_408119;
   reg _408120_408120 ; 
   reg __408120_408120;
   reg _408121_408121 ; 
   reg __408121_408121;
   reg _408122_408122 ; 
   reg __408122_408122;
   reg _408123_408123 ; 
   reg __408123_408123;
   reg _408124_408124 ; 
   reg __408124_408124;
   reg _408125_408125 ; 
   reg __408125_408125;
   reg _408126_408126 ; 
   reg __408126_408126;
   reg _408127_408127 ; 
   reg __408127_408127;
   reg _408128_408128 ; 
   reg __408128_408128;
   reg _408129_408129 ; 
   reg __408129_408129;
   reg _408130_408130 ; 
   reg __408130_408130;
   reg _408131_408131 ; 
   reg __408131_408131;
   reg _408132_408132 ; 
   reg __408132_408132;
   reg _408133_408133 ; 
   reg __408133_408133;
   reg _408134_408134 ; 
   reg __408134_408134;
   reg _408135_408135 ; 
   reg __408135_408135;
   reg _408136_408136 ; 
   reg __408136_408136;
   reg _408137_408137 ; 
   reg __408137_408137;
   reg _408138_408138 ; 
   reg __408138_408138;
   reg _408139_408139 ; 
   reg __408139_408139;
   reg _408140_408140 ; 
   reg __408140_408140;
   reg _408141_408141 ; 
   reg __408141_408141;
   reg _408142_408142 ; 
   reg __408142_408142;
   reg _408143_408143 ; 
   reg __408143_408143;
   reg _408144_408144 ; 
   reg __408144_408144;
   reg _408145_408145 ; 
   reg __408145_408145;
   reg _408146_408146 ; 
   reg __408146_408146;
   reg _408147_408147 ; 
   reg __408147_408147;
   reg _408148_408148 ; 
   reg __408148_408148;
   reg _408149_408149 ; 
   reg __408149_408149;
   reg _408150_408150 ; 
   reg __408150_408150;
   reg _408151_408151 ; 
   reg __408151_408151;
   reg _408152_408152 ; 
   reg __408152_408152;
   reg _408153_408153 ; 
   reg __408153_408153;
   reg _408154_408154 ; 
   reg __408154_408154;
   reg _408155_408155 ; 
   reg __408155_408155;
   reg _408156_408156 ; 
   reg __408156_408156;
   reg _408157_408157 ; 
   reg __408157_408157;
   reg _408158_408158 ; 
   reg __408158_408158;
   reg _408159_408159 ; 
   reg __408159_408159;
   reg _408160_408160 ; 
   reg __408160_408160;
   reg _408161_408161 ; 
   reg __408161_408161;
   reg _408162_408162 ; 
   reg __408162_408162;
   reg _408163_408163 ; 
   reg __408163_408163;
   reg _408164_408164 ; 
   reg __408164_408164;
   reg _408165_408165 ; 
   reg __408165_408165;
   reg _408166_408166 ; 
   reg __408166_408166;
   reg _408167_408167 ; 
   reg __408167_408167;
   reg _408168_408168 ; 
   reg __408168_408168;
   reg _408169_408169 ; 
   reg __408169_408169;
   reg _408170_408170 ; 
   reg __408170_408170;
   reg _408171_408171 ; 
   reg __408171_408171;
   reg _408172_408172 ; 
   reg __408172_408172;
   reg _408173_408173 ; 
   reg __408173_408173;
   reg _408174_408174 ; 
   reg __408174_408174;
   reg _408175_408175 ; 
   reg __408175_408175;
   reg _408176_408176 ; 
   reg __408176_408176;
   reg _408177_408177 ; 
   reg __408177_408177;
   reg _408178_408178 ; 
   reg __408178_408178;
   reg _408179_408179 ; 
   reg __408179_408179;
   reg _408180_408180 ; 
   reg __408180_408180;
   reg _408181_408181 ; 
   reg __408181_408181;
   reg _408182_408182 ; 
   reg __408182_408182;
   reg _408183_408183 ; 
   reg __408183_408183;
   reg _408184_408184 ; 
   reg __408184_408184;
   reg _408185_408185 ; 
   reg __408185_408185;
   reg _408186_408186 ; 
   reg __408186_408186;
   reg _408187_408187 ; 
   reg __408187_408187;
   reg _408188_408188 ; 
   reg __408188_408188;
   reg _408189_408189 ; 
   reg __408189_408189;
   reg _408190_408190 ; 
   reg __408190_408190;
   reg _408191_408191 ; 
   reg __408191_408191;
   reg _408192_408192 ; 
   reg __408192_408192;
   reg _408193_408193 ; 
   reg __408193_408193;
   reg _408194_408194 ; 
   reg __408194_408194;
   reg _408195_408195 ; 
   reg __408195_408195;
   reg _408196_408196 ; 
   reg __408196_408196;
   reg _408197_408197 ; 
   reg __408197_408197;
   reg _408198_408198 ; 
   reg __408198_408198;
   reg _408199_408199 ; 
   reg __408199_408199;
   reg _408200_408200 ; 
   reg __408200_408200;
   reg _408201_408201 ; 
   reg __408201_408201;
   reg _408202_408202 ; 
   reg __408202_408202;
   reg _408203_408203 ; 
   reg __408203_408203;
   reg _408204_408204 ; 
   reg __408204_408204;
   reg _408205_408205 ; 
   reg __408205_408205;
   reg _408206_408206 ; 
   reg __408206_408206;
   reg _408207_408207 ; 
   reg __408207_408207;
   reg _408208_408208 ; 
   reg __408208_408208;
   reg _408209_408209 ; 
   reg __408209_408209;
   reg _408210_408210 ; 
   reg __408210_408210;
   reg _408211_408211 ; 
   reg __408211_408211;
   reg _408212_408212 ; 
   reg __408212_408212;
   reg _408213_408213 ; 
   reg __408213_408213;
   reg _408214_408214 ; 
   reg __408214_408214;
   reg _408215_408215 ; 
   reg __408215_408215;
   reg _408216_408216 ; 
   reg __408216_408216;
   reg _408217_408217 ; 
   reg __408217_408217;
   reg _408218_408218 ; 
   reg __408218_408218;
   reg _408219_408219 ; 
   reg __408219_408219;
   reg _408220_408220 ; 
   reg __408220_408220;
   reg _408221_408221 ; 
   reg __408221_408221;
   reg _408222_408222 ; 
   reg __408222_408222;
   reg _408223_408223 ; 
   reg __408223_408223;
   reg _408224_408224 ; 
   reg __408224_408224;
   reg _408225_408225 ; 
   reg __408225_408225;
   reg _408226_408226 ; 
   reg __408226_408226;
   reg _408227_408227 ; 
   reg __408227_408227;
   reg _408228_408228 ; 
   reg __408228_408228;
   reg _408229_408229 ; 
   reg __408229_408229;
   reg _408230_408230 ; 
   reg __408230_408230;
   reg _408231_408231 ; 
   reg __408231_408231;
   reg _408232_408232 ; 
   reg __408232_408232;
   reg _408233_408233 ; 
   reg __408233_408233;
   reg _408234_408234 ; 
   reg __408234_408234;
   reg _408235_408235 ; 
   reg __408235_408235;
   reg _408236_408236 ; 
   reg __408236_408236;
   reg _408237_408237 ; 
   reg __408237_408237;
   reg _408238_408238 ; 
   reg __408238_408238;
   reg _408239_408239 ; 
   reg __408239_408239;
   reg _408240_408240 ; 
   reg __408240_408240;
   reg _408241_408241 ; 
   reg __408241_408241;
   reg _408242_408242 ; 
   reg __408242_408242;
   reg _408243_408243 ; 
   reg __408243_408243;
   reg _408244_408244 ; 
   reg __408244_408244;
   reg _408245_408245 ; 
   reg __408245_408245;
   reg _408246_408246 ; 
   reg __408246_408246;
   reg _408247_408247 ; 
   reg __408247_408247;
   reg _408248_408248 ; 
   reg __408248_408248;
   reg _408249_408249 ; 
   reg __408249_408249;
   reg _408250_408250 ; 
   reg __408250_408250;
   reg _408251_408251 ; 
   reg __408251_408251;
   reg _408252_408252 ; 
   reg __408252_408252;
   reg _408253_408253 ; 
   reg __408253_408253;
   reg _408254_408254 ; 
   reg __408254_408254;
   reg _408255_408255 ; 
   reg __408255_408255;
   reg _408256_408256 ; 
   reg __408256_408256;
   reg _408257_408257 ; 
   reg __408257_408257;
   reg _408258_408258 ; 
   reg __408258_408258;
   reg _408259_408259 ; 
   reg __408259_408259;
   reg _408260_408260 ; 
   reg __408260_408260;
   reg _408261_408261 ; 
   reg __408261_408261;
   reg _408262_408262 ; 
   reg __408262_408262;
   reg _408263_408263 ; 
   reg __408263_408263;
   reg _408264_408264 ; 
   reg __408264_408264;
   reg _408265_408265 ; 
   reg __408265_408265;
   reg _408266_408266 ; 
   reg __408266_408266;
   reg _408267_408267 ; 
   reg __408267_408267;
   reg _408268_408268 ; 
   reg __408268_408268;
   reg _408269_408269 ; 
   reg __408269_408269;
   reg _408270_408270 ; 
   reg __408270_408270;
   reg _408271_408271 ; 
   reg __408271_408271;
   reg _408272_408272 ; 
   reg __408272_408272;
   reg _408273_408273 ; 
   reg __408273_408273;
   reg _408274_408274 ; 
   reg __408274_408274;
   reg _408275_408275 ; 
   reg __408275_408275;
   reg _408276_408276 ; 
   reg __408276_408276;
   reg _408277_408277 ; 
   reg __408277_408277;
   reg _408278_408278 ; 
   reg __408278_408278;
   reg _408279_408279 ; 
   reg __408279_408279;
   reg _408280_408280 ; 
   reg __408280_408280;
   reg _408281_408281 ; 
   reg __408281_408281;
   reg _408282_408282 ; 
   reg __408282_408282;
   reg _408283_408283 ; 
   reg __408283_408283;
   reg _408284_408284 ; 
   reg __408284_408284;
   reg _408285_408285 ; 
   reg __408285_408285;
   reg _408286_408286 ; 
   reg __408286_408286;
   reg _408287_408287 ; 
   reg __408287_408287;
   reg _408288_408288 ; 
   reg __408288_408288;
   reg _408289_408289 ; 
   reg __408289_408289;
   reg _408290_408290 ; 
   reg __408290_408290;
   reg _408291_408291 ; 
   reg __408291_408291;
   reg _408292_408292 ; 
   reg __408292_408292;
   reg _408293_408293 ; 
   reg __408293_408293;
   reg _408294_408294 ; 
   reg __408294_408294;
   reg _408295_408295 ; 
   reg __408295_408295;
   reg _408296_408296 ; 
   reg __408296_408296;
   reg _408297_408297 ; 
   reg __408297_408297;
   reg _408298_408298 ; 
   reg __408298_408298;
   reg _408299_408299 ; 
   reg __408299_408299;
   reg _408300_408300 ; 
   reg __408300_408300;
   reg _408301_408301 ; 
   reg __408301_408301;
   reg _408302_408302 ; 
   reg __408302_408302;
   reg _408303_408303 ; 
   reg __408303_408303;
   reg _408304_408304 ; 
   reg __408304_408304;
   reg _408305_408305 ; 
   reg __408305_408305;
   reg _408306_408306 ; 
   reg __408306_408306;
   reg _408307_408307 ; 
   reg __408307_408307;
   reg _408308_408308 ; 
   reg __408308_408308;
   reg _408309_408309 ; 
   reg __408309_408309;
   reg _408310_408310 ; 
   reg __408310_408310;
   reg _408311_408311 ; 
   reg __408311_408311;
   reg _408312_408312 ; 
   reg __408312_408312;
   reg _408313_408313 ; 
   reg __408313_408313;
   reg _408314_408314 ; 
   reg __408314_408314;
   reg _408315_408315 ; 
   reg __408315_408315;
   reg _408316_408316 ; 
   reg __408316_408316;
   reg _408317_408317 ; 
   reg __408317_408317;
   reg _408318_408318 ; 
   reg __408318_408318;
   reg _408319_408319 ; 
   reg __408319_408319;
   reg _408320_408320 ; 
   reg __408320_408320;
   reg _408321_408321 ; 
   reg __408321_408321;
   reg _408322_408322 ; 
   reg __408322_408322;
   reg _408323_408323 ; 
   reg __408323_408323;
   reg _408324_408324 ; 
   reg __408324_408324;
   reg _408325_408325 ; 
   reg __408325_408325;
   reg _408326_408326 ; 
   reg __408326_408326;
   reg _408327_408327 ; 
   reg __408327_408327;
   reg _408328_408328 ; 
   reg __408328_408328;
   reg _408329_408329 ; 
   reg __408329_408329;
   reg _408330_408330 ; 
   reg __408330_408330;
   reg _408331_408331 ; 
   reg __408331_408331;
   reg _408332_408332 ; 
   reg __408332_408332;
   reg _408333_408333 ; 
   reg __408333_408333;
   reg _408334_408334 ; 
   reg __408334_408334;
   reg _408335_408335 ; 
   reg __408335_408335;
   reg _408336_408336 ; 
   reg __408336_408336;
   reg _408337_408337 ; 
   reg __408337_408337;
   reg _408338_408338 ; 
   reg __408338_408338;
   reg _408339_408339 ; 
   reg __408339_408339;
   reg _408340_408340 ; 
   reg __408340_408340;
   reg _408341_408341 ; 
   reg __408341_408341;
   reg _408342_408342 ; 
   reg __408342_408342;
   reg _408343_408343 ; 
   reg __408343_408343;
   reg _408344_408344 ; 
   reg __408344_408344;
   reg _408345_408345 ; 
   reg __408345_408345;
   reg _408346_408346 ; 
   reg __408346_408346;
   reg _408347_408347 ; 
   reg __408347_408347;
   reg _408348_408348 ; 
   reg __408348_408348;
   reg _408349_408349 ; 
   reg __408349_408349;
   reg _408350_408350 ; 
   reg __408350_408350;
   reg _408351_408351 ; 
   reg __408351_408351;
   reg _408352_408352 ; 
   reg __408352_408352;
   reg _408353_408353 ; 
   reg __408353_408353;
   reg _408354_408354 ; 
   reg __408354_408354;
   reg _408355_408355 ; 
   reg __408355_408355;
   reg _408356_408356 ; 
   reg __408356_408356;
   reg _408357_408357 ; 
   reg __408357_408357;
   reg _408358_408358 ; 
   reg __408358_408358;
   reg _408359_408359 ; 
   reg __408359_408359;
   reg _408360_408360 ; 
   reg __408360_408360;
   reg _408361_408361 ; 
   reg __408361_408361;
   reg _408362_408362 ; 
   reg __408362_408362;
   reg _408363_408363 ; 
   reg __408363_408363;
   reg _408364_408364 ; 
   reg __408364_408364;
   reg _408365_408365 ; 
   reg __408365_408365;
   reg _408366_408366 ; 
   reg __408366_408366;
   reg _408367_408367 ; 
   reg __408367_408367;
   reg _408368_408368 ; 
   reg __408368_408368;
   reg _408369_408369 ; 
   reg __408369_408369;
   reg _408370_408370 ; 
   reg __408370_408370;
   reg _408371_408371 ; 
   reg __408371_408371;
   reg _408372_408372 ; 
   reg __408372_408372;
   reg _408373_408373 ; 
   reg __408373_408373;
   reg _408374_408374 ; 
   reg __408374_408374;
   reg _408375_408375 ; 
   reg __408375_408375;
   reg _408376_408376 ; 
   reg __408376_408376;
   reg _408377_408377 ; 
   reg __408377_408377;
   reg _408378_408378 ; 
   reg __408378_408378;
   reg _408379_408379 ; 
   reg __408379_408379;
   reg _408380_408380 ; 
   reg __408380_408380;
   reg _408381_408381 ; 
   reg __408381_408381;
   reg _408382_408382 ; 
   reg __408382_408382;
   reg _408383_408383 ; 
   reg __408383_408383;
   reg _408384_408384 ; 
   reg __408384_408384;
   reg _408385_408385 ; 
   reg __408385_408385;
   reg _408386_408386 ; 
   reg __408386_408386;
   reg _408387_408387 ; 
   reg __408387_408387;
   reg _408388_408388 ; 
   reg __408388_408388;
   reg _408389_408389 ; 
   reg __408389_408389;
   reg _408390_408390 ; 
   reg __408390_408390;
   reg _408391_408391 ; 
   reg __408391_408391;
   reg _408392_408392 ; 
   reg __408392_408392;
   reg _408393_408393 ; 
   reg __408393_408393;
   reg _408394_408394 ; 
   reg __408394_408394;
   reg _408395_408395 ; 
   reg __408395_408395;
   reg _408396_408396 ; 
   reg __408396_408396;
   reg _408397_408397 ; 
   reg __408397_408397;
   reg _408398_408398 ; 
   reg __408398_408398;
   reg _408399_408399 ; 
   reg __408399_408399;
   reg _408400_408400 ; 
   reg __408400_408400;
   reg _408401_408401 ; 
   reg __408401_408401;
   reg _408402_408402 ; 
   reg __408402_408402;
   reg _408403_408403 ; 
   reg __408403_408403;
   reg _408404_408404 ; 
   reg __408404_408404;
   reg _408405_408405 ; 
   reg __408405_408405;
   reg _408406_408406 ; 
   reg __408406_408406;
   reg _408407_408407 ; 
   reg __408407_408407;
   reg _408408_408408 ; 
   reg __408408_408408;
   reg _408409_408409 ; 
   reg __408409_408409;
   reg _408410_408410 ; 
   reg __408410_408410;
   reg _408411_408411 ; 
   reg __408411_408411;
   reg _408412_408412 ; 
   reg __408412_408412;
   reg _408413_408413 ; 
   reg __408413_408413;
   reg _408414_408414 ; 
   reg __408414_408414;
   reg _408415_408415 ; 
   reg __408415_408415;
   reg _408416_408416 ; 
   reg __408416_408416;
   reg _408417_408417 ; 
   reg __408417_408417;
   reg _408418_408418 ; 
   reg __408418_408418;
   reg _408419_408419 ; 
   reg __408419_408419;
   reg _408420_408420 ; 
   reg __408420_408420;
   reg _408421_408421 ; 
   reg __408421_408421;
   reg _408422_408422 ; 
   reg __408422_408422;
   reg _408423_408423 ; 
   reg __408423_408423;
   reg _408424_408424 ; 
   reg __408424_408424;
   reg _408425_408425 ; 
   reg __408425_408425;
   reg _408426_408426 ; 
   reg __408426_408426;
   reg _408427_408427 ; 
   reg __408427_408427;
   reg _408428_408428 ; 
   reg __408428_408428;
   reg _408429_408429 ; 
   reg __408429_408429;
   reg _408430_408430 ; 
   reg __408430_408430;
   reg _408431_408431 ; 
   reg __408431_408431;
   reg _408432_408432 ; 
   reg __408432_408432;
   reg _408433_408433 ; 
   reg __408433_408433;
   reg _408434_408434 ; 
   reg __408434_408434;
   reg _408435_408435 ; 
   reg __408435_408435;
   reg _408436_408436 ; 
   reg __408436_408436;
   reg _408437_408437 ; 
   reg __408437_408437;
   reg _408438_408438 ; 
   reg __408438_408438;
   reg _408439_408439 ; 
   reg __408439_408439;
   reg _408440_408440 ; 
   reg __408440_408440;
   reg _408441_408441 ; 
   reg __408441_408441;
   reg _408442_408442 ; 
   reg __408442_408442;
   reg _408443_408443 ; 
   reg __408443_408443;
   reg _408444_408444 ; 
   reg __408444_408444;
   reg _408445_408445 ; 
   reg __408445_408445;
   reg _408446_408446 ; 
   reg __408446_408446;
   reg _408447_408447 ; 
   reg __408447_408447;
   reg _408448_408448 ; 
   reg __408448_408448;
   reg _408449_408449 ; 
   reg __408449_408449;
   reg _408450_408450 ; 
   reg __408450_408450;
   reg _408451_408451 ; 
   reg __408451_408451;
   reg _408452_408452 ; 
   reg __408452_408452;
   reg _408453_408453 ; 
   reg __408453_408453;
   reg _408454_408454 ; 
   reg __408454_408454;
   reg _408455_408455 ; 
   reg __408455_408455;
   reg _408456_408456 ; 
   reg __408456_408456;
   reg _408457_408457 ; 
   reg __408457_408457;
   reg _408458_408458 ; 
   reg __408458_408458;
   reg _408459_408459 ; 
   reg __408459_408459;
   reg _408460_408460 ; 
   reg __408460_408460;
   reg _408461_408461 ; 
   reg __408461_408461;
   reg _408462_408462 ; 
   reg __408462_408462;
   reg _408463_408463 ; 
   reg __408463_408463;
   reg _408464_408464 ; 
   reg __408464_408464;
   reg _408465_408465 ; 
   reg __408465_408465;
   reg _408466_408466 ; 
   reg __408466_408466;
   reg _408467_408467 ; 
   reg __408467_408467;
   reg _408468_408468 ; 
   reg __408468_408468;
   reg _408469_408469 ; 
   reg __408469_408469;
   reg _408470_408470 ; 
   reg __408470_408470;
   reg _408471_408471 ; 
   reg __408471_408471;
   reg _408472_408472 ; 
   reg __408472_408472;
   reg _408473_408473 ; 
   reg __408473_408473;
   reg _408474_408474 ; 
   reg __408474_408474;
   reg _408475_408475 ; 
   reg __408475_408475;
   reg _408476_408476 ; 
   reg __408476_408476;
   reg _408477_408477 ; 
   reg __408477_408477;
   reg _408478_408478 ; 
   reg __408478_408478;
   reg _408479_408479 ; 
   reg __408479_408479;
   reg _408480_408480 ; 
   reg __408480_408480;
   reg _408481_408481 ; 
   reg __408481_408481;
   reg _408482_408482 ; 
   reg __408482_408482;
   reg _408483_408483 ; 
   reg __408483_408483;
   reg _408484_408484 ; 
   reg __408484_408484;
   reg _408485_408485 ; 
   reg __408485_408485;
   reg _408486_408486 ; 
   reg __408486_408486;
   reg _408487_408487 ; 
   reg __408487_408487;
   reg _408488_408488 ; 
   reg __408488_408488;
   reg _408489_408489 ; 
   reg __408489_408489;
   reg _408490_408490 ; 
   reg __408490_408490;
   reg _408491_408491 ; 
   reg __408491_408491;
   reg _408492_408492 ; 
   reg __408492_408492;
   reg _408493_408493 ; 
   reg __408493_408493;
   reg _408494_408494 ; 
   reg __408494_408494;
   reg _408495_408495 ; 
   reg __408495_408495;
   reg _408496_408496 ; 
   reg __408496_408496;
   reg _408497_408497 ; 
   reg __408497_408497;
   reg _408498_408498 ; 
   reg __408498_408498;
   reg _408499_408499 ; 
   reg __408499_408499;
   reg _408500_408500 ; 
   reg __408500_408500;
   reg _408501_408501 ; 
   reg __408501_408501;
   reg _408502_408502 ; 
   reg __408502_408502;
   reg _408503_408503 ; 
   reg __408503_408503;
   reg _408504_408504 ; 
   reg __408504_408504;
   reg _408505_408505 ; 
   reg __408505_408505;
   reg _408506_408506 ; 
   reg __408506_408506;
   reg _408507_408507 ; 
   reg __408507_408507;
   reg _408508_408508 ; 
   reg __408508_408508;
   reg _408509_408509 ; 
   reg __408509_408509;
   reg _408510_408510 ; 
   reg __408510_408510;
   reg _408511_408511 ; 
   reg __408511_408511;
   reg _408512_408512 ; 
   reg __408512_408512;
   reg _408513_408513 ; 
   reg __408513_408513;
   reg _408514_408514 ; 
   reg __408514_408514;
   reg _408515_408515 ; 
   reg __408515_408515;
   reg _408516_408516 ; 
   reg __408516_408516;
   reg _408517_408517 ; 
   reg __408517_408517;
   reg _408518_408518 ; 
   reg __408518_408518;
   reg _408519_408519 ; 
   reg __408519_408519;
   reg _408520_408520 ; 
   reg __408520_408520;
   reg _408521_408521 ; 
   reg __408521_408521;
   reg _408522_408522 ; 
   reg __408522_408522;
   reg _408523_408523 ; 
   reg __408523_408523;
   reg _408524_408524 ; 
   reg __408524_408524;
   reg _408525_408525 ; 
   reg __408525_408525;
   reg _408526_408526 ; 
   reg __408526_408526;
   reg _408527_408527 ; 
   reg __408527_408527;
   reg _408528_408528 ; 
   reg __408528_408528;
   reg _408529_408529 ; 
   reg __408529_408529;
   reg _408530_408530 ; 
   reg __408530_408530;
   reg _408531_408531 ; 
   reg __408531_408531;
   reg _408532_408532 ; 
   reg __408532_408532;
   reg _408533_408533 ; 
   reg __408533_408533;
   reg _408534_408534 ; 
   reg __408534_408534;
   reg _408535_408535 ; 
   reg __408535_408535;
   reg _408536_408536 ; 
   reg __408536_408536;
   reg _408537_408537 ; 
   reg __408537_408537;
   reg _408538_408538 ; 
   reg __408538_408538;
   reg _408539_408539 ; 
   reg __408539_408539;
   reg _408540_408540 ; 
   reg __408540_408540;
   reg _408541_408541 ; 
   reg __408541_408541;
   reg _408542_408542 ; 
   reg __408542_408542;
   reg _408543_408543 ; 
   reg __408543_408543;
   reg _408544_408544 ; 
   reg __408544_408544;
   reg _408545_408545 ; 
   reg __408545_408545;
   reg _408546_408546 ; 
   reg __408546_408546;
   reg _408547_408547 ; 
   reg __408547_408547;
   reg _408548_408548 ; 
   reg __408548_408548;
   reg _408549_408549 ; 
   reg __408549_408549;
   reg _408550_408550 ; 
   reg __408550_408550;
   reg _408551_408551 ; 
   reg __408551_408551;
   reg _408552_408552 ; 
   reg __408552_408552;
   reg _408553_408553 ; 
   reg __408553_408553;
   reg _408554_408554 ; 
   reg __408554_408554;
   reg _408555_408555 ; 
   reg __408555_408555;
   reg _408556_408556 ; 
   reg __408556_408556;
   reg _408557_408557 ; 
   reg __408557_408557;
   reg _408558_408558 ; 
   reg __408558_408558;
   reg _408559_408559 ; 
   reg __408559_408559;
   reg _408560_408560 ; 
   reg __408560_408560;
   reg _408561_408561 ; 
   reg __408561_408561;
   reg _408562_408562 ; 
   reg __408562_408562;
   reg _408563_408563 ; 
   reg __408563_408563;
   reg _408564_408564 ; 
   reg __408564_408564;
   reg _408565_408565 ; 
   reg __408565_408565;
   reg _408566_408566 ; 
   reg __408566_408566;
   reg _408567_408567 ; 
   reg __408567_408567;
   reg _408568_408568 ; 
   reg __408568_408568;
   reg _408569_408569 ; 
   reg __408569_408569;
   reg _408570_408570 ; 
   reg __408570_408570;
   reg _408571_408571 ; 
   reg __408571_408571;
   reg _408572_408572 ; 
   reg __408572_408572;
   reg _408573_408573 ; 
   reg __408573_408573;
   reg _408574_408574 ; 
   reg __408574_408574;
   reg _408575_408575 ; 
   reg __408575_408575;
   reg _408576_408576 ; 
   reg __408576_408576;
   reg _408577_408577 ; 
   reg __408577_408577;
   reg _408578_408578 ; 
   reg __408578_408578;
   reg _408579_408579 ; 
   reg __408579_408579;
   reg _408580_408580 ; 
   reg __408580_408580;
   reg _408581_408581 ; 
   reg __408581_408581;
   reg _408582_408582 ; 
   reg __408582_408582;
   reg _408583_408583 ; 
   reg __408583_408583;
   reg _408584_408584 ; 
   reg __408584_408584;
   reg _408585_408585 ; 
   reg __408585_408585;
   reg _408586_408586 ; 
   reg __408586_408586;
   reg _408587_408587 ; 
   reg __408587_408587;
   reg _408588_408588 ; 
   reg __408588_408588;
   reg _408589_408589 ; 
   reg __408589_408589;
   reg _408590_408590 ; 
   reg __408590_408590;
   reg _408591_408591 ; 
   reg __408591_408591;
   reg _408592_408592 ; 
   reg __408592_408592;
   reg _408593_408593 ; 
   reg __408593_408593;
   reg _408594_408594 ; 
   reg __408594_408594;
   reg _408595_408595 ; 
   reg __408595_408595;
   reg _408596_408596 ; 
   reg __408596_408596;
   reg _408597_408597 ; 
   reg __408597_408597;
   reg _408598_408598 ; 
   reg __408598_408598;
   reg _408599_408599 ; 
   reg __408599_408599;
   reg _408600_408600 ; 
   reg __408600_408600;
   reg _408601_408601 ; 
   reg __408601_408601;
   reg _408602_408602 ; 
   reg __408602_408602;
   reg _408603_408603 ; 
   reg __408603_408603;
   reg _408604_408604 ; 
   reg __408604_408604;
   reg _408605_408605 ; 
   reg __408605_408605;
   reg _408606_408606 ; 
   reg __408606_408606;
   reg _408607_408607 ; 
   reg __408607_408607;
   reg _408608_408608 ; 
   reg __408608_408608;
   reg _408609_408609 ; 
   reg __408609_408609;
   reg _408610_408610 ; 
   reg __408610_408610;
   reg _408611_408611 ; 
   reg __408611_408611;
   reg _408612_408612 ; 
   reg __408612_408612;
   reg _408613_408613 ; 
   reg __408613_408613;
   reg _408614_408614 ; 
   reg __408614_408614;
   reg _408615_408615 ; 
   reg __408615_408615;
   reg _408616_408616 ; 
   reg __408616_408616;
   reg _408617_408617 ; 
   reg __408617_408617;
   reg _408618_408618 ; 
   reg __408618_408618;
   reg _408619_408619 ; 
   reg __408619_408619;
   reg _408620_408620 ; 
   reg __408620_408620;
   reg _408621_408621 ; 
   reg __408621_408621;
   reg _408622_408622 ; 
   reg __408622_408622;
   reg _408623_408623 ; 
   reg __408623_408623;
   reg _408624_408624 ; 
   reg __408624_408624;
   reg _408625_408625 ; 
   reg __408625_408625;
   reg _408626_408626 ; 
   reg __408626_408626;
   reg _408627_408627 ; 
   reg __408627_408627;
   reg _408628_408628 ; 
   reg __408628_408628;
   reg _408629_408629 ; 
   reg __408629_408629;
   reg _408630_408630 ; 
   reg __408630_408630;
   reg _408631_408631 ; 
   reg __408631_408631;
   reg _408632_408632 ; 
   reg __408632_408632;
   reg _408633_408633 ; 
   reg __408633_408633;
   reg _408634_408634 ; 
   reg __408634_408634;
   reg _408635_408635 ; 
   reg __408635_408635;
   reg _408636_408636 ; 
   reg __408636_408636;
   reg _408637_408637 ; 
   reg __408637_408637;
   reg _408638_408638 ; 
   reg __408638_408638;
   reg _408639_408639 ; 
   reg __408639_408639;
   reg _408640_408640 ; 
   reg __408640_408640;
   reg _408641_408641 ; 
   reg __408641_408641;
   reg _408642_408642 ; 
   reg __408642_408642;
   reg _408643_408643 ; 
   reg __408643_408643;
   reg _408644_408644 ; 
   reg __408644_408644;
   reg _408645_408645 ; 
   reg __408645_408645;
   reg _408646_408646 ; 
   reg __408646_408646;
   reg _408647_408647 ; 
   reg __408647_408647;
   reg _408648_408648 ; 
   reg __408648_408648;
   reg _408649_408649 ; 
   reg __408649_408649;
   reg _408650_408650 ; 
   reg __408650_408650;
   reg _408651_408651 ; 
   reg __408651_408651;
   reg _408652_408652 ; 
   reg __408652_408652;
   reg _408653_408653 ; 
   reg __408653_408653;
   reg _408654_408654 ; 
   reg __408654_408654;
   reg _408655_408655 ; 
   reg __408655_408655;
   reg _408656_408656 ; 
   reg __408656_408656;
   reg _408657_408657 ; 
   reg __408657_408657;
   reg _408658_408658 ; 
   reg __408658_408658;
   reg _408659_408659 ; 
   reg __408659_408659;
   reg _408660_408660 ; 
   reg __408660_408660;
   reg _408661_408661 ; 
   reg __408661_408661;
   reg _408662_408662 ; 
   reg __408662_408662;
   reg _408663_408663 ; 
   reg __408663_408663;
   reg _408664_408664 ; 
   reg __408664_408664;
   reg _408665_408665 ; 
   reg __408665_408665;
   reg _408666_408666 ; 
   reg __408666_408666;
   reg _408667_408667 ; 
   reg __408667_408667;
   reg _408668_408668 ; 
   reg __408668_408668;
   reg _408669_408669 ; 
   reg __408669_408669;
   reg _408670_408670 ; 
   reg __408670_408670;
   reg _408671_408671 ; 
   reg __408671_408671;
   reg _408672_408672 ; 
   reg __408672_408672;
   reg _408673_408673 ; 
   reg __408673_408673;
   reg _408674_408674 ; 
   reg __408674_408674;
   reg _408675_408675 ; 
   reg __408675_408675;
   reg _408676_408676 ; 
   reg __408676_408676;
   reg _408677_408677 ; 
   reg __408677_408677;
   reg _408678_408678 ; 
   reg __408678_408678;
   reg _408679_408679 ; 
   reg __408679_408679;
   reg _408680_408680 ; 
   reg __408680_408680;
   reg _408681_408681 ; 
   reg __408681_408681;
   reg _408682_408682 ; 
   reg __408682_408682;
   reg _408683_408683 ; 
   reg __408683_408683;
   reg _408684_408684 ; 
   reg __408684_408684;
   reg _408685_408685 ; 
   reg __408685_408685;
   reg _408686_408686 ; 
   reg __408686_408686;
   reg _408687_408687 ; 
   reg __408687_408687;
   reg _408688_408688 ; 
   reg __408688_408688;
   reg _408689_408689 ; 
   reg __408689_408689;
   reg _408690_408690 ; 
   reg __408690_408690;
   reg _408691_408691 ; 
   reg __408691_408691;
   reg _408692_408692 ; 
   reg __408692_408692;
   reg _408693_408693 ; 
   reg __408693_408693;
   reg _408694_408694 ; 
   reg __408694_408694;
   reg _408695_408695 ; 
   reg __408695_408695;
   reg _408696_408696 ; 
   reg __408696_408696;
   reg _408697_408697 ; 
   reg __408697_408697;
   reg _408698_408698 ; 
   reg __408698_408698;
   reg _408699_408699 ; 
   reg __408699_408699;
   reg _408700_408700 ; 
   reg __408700_408700;
   reg _408701_408701 ; 
   reg __408701_408701;
   reg _408702_408702 ; 
   reg __408702_408702;
   reg _408703_408703 ; 
   reg __408703_408703;
   reg _408704_408704 ; 
   reg __408704_408704;
   reg _408705_408705 ; 
   reg __408705_408705;
   reg _408706_408706 ; 
   reg __408706_408706;
   reg _408707_408707 ; 
   reg __408707_408707;
   reg _408708_408708 ; 
   reg __408708_408708;
   reg _408709_408709 ; 
   reg __408709_408709;
   reg _408710_408710 ; 
   reg __408710_408710;
   reg _408711_408711 ; 
   reg __408711_408711;
   reg _408712_408712 ; 
   reg __408712_408712;
   reg _408713_408713 ; 
   reg __408713_408713;
   reg _408714_408714 ; 
   reg __408714_408714;
   reg _408715_408715 ; 
   reg __408715_408715;
   reg _408716_408716 ; 
   reg __408716_408716;
   reg _408717_408717 ; 
   reg __408717_408717;
   reg _408718_408718 ; 
   reg __408718_408718;
   reg _408719_408719 ; 
   reg __408719_408719;
   reg _408720_408720 ; 
   reg __408720_408720;
   reg _408721_408721 ; 
   reg __408721_408721;
   reg _408722_408722 ; 
   reg __408722_408722;
   reg _408723_408723 ; 
   reg __408723_408723;
   reg _408724_408724 ; 
   reg __408724_408724;
   reg _408725_408725 ; 
   reg __408725_408725;
   reg _408726_408726 ; 
   reg __408726_408726;
   reg _408727_408727 ; 
   reg __408727_408727;
   reg _408728_408728 ; 
   reg __408728_408728;
   reg _408729_408729 ; 
   reg __408729_408729;
   reg _408730_408730 ; 
   reg __408730_408730;
   reg _408731_408731 ; 
   reg __408731_408731;
   reg _408732_408732 ; 
   reg __408732_408732;
   reg _408733_408733 ; 
   reg __408733_408733;
   reg _408734_408734 ; 
   reg __408734_408734;
   reg _408735_408735 ; 
   reg __408735_408735;
   reg _408736_408736 ; 
   reg __408736_408736;
   reg _408737_408737 ; 
   reg __408737_408737;
   reg _408738_408738 ; 
   reg __408738_408738;
   reg _408739_408739 ; 
   reg __408739_408739;
   reg _408740_408740 ; 
   reg __408740_408740;
   reg _408741_408741 ; 
   reg __408741_408741;
   reg _408742_408742 ; 
   reg __408742_408742;
   reg _408743_408743 ; 
   reg __408743_408743;
   reg _408744_408744 ; 
   reg __408744_408744;
   reg _408745_408745 ; 
   reg __408745_408745;
   reg _408746_408746 ; 
   reg __408746_408746;
   reg _408747_408747 ; 
   reg __408747_408747;
   reg _408748_408748 ; 
   reg __408748_408748;
   reg _408749_408749 ; 
   reg __408749_408749;
   reg _408750_408750 ; 
   reg __408750_408750;
   reg _408751_408751 ; 
   reg __408751_408751;
   reg _408752_408752 ; 
   reg __408752_408752;
   reg _408753_408753 ; 
   reg __408753_408753;
   reg _408754_408754 ; 
   reg __408754_408754;
   reg _408755_408755 ; 
   reg __408755_408755;
   reg _408756_408756 ; 
   reg __408756_408756;
   reg _408757_408757 ; 
   reg __408757_408757;
   reg _408758_408758 ; 
   reg __408758_408758;
   reg _408759_408759 ; 
   reg __408759_408759;
   reg _408760_408760 ; 
   reg __408760_408760;
   reg _408761_408761 ; 
   reg __408761_408761;
   reg _408762_408762 ; 
   reg __408762_408762;
   reg _408763_408763 ; 
   reg __408763_408763;
   reg _408764_408764 ; 
   reg __408764_408764;
   reg _408765_408765 ; 
   reg __408765_408765;
   reg _408766_408766 ; 
   reg __408766_408766;
   reg _408767_408767 ; 
   reg __408767_408767;
   reg _408768_408768 ; 
   reg __408768_408768;
   reg _408769_408769 ; 
   reg __408769_408769;
   reg _408770_408770 ; 
   reg __408770_408770;
   reg _408771_408771 ; 
   reg __408771_408771;
   reg _408772_408772 ; 
   reg __408772_408772;
   reg _408773_408773 ; 
   reg __408773_408773;
   reg _408774_408774 ; 
   reg __408774_408774;
   reg _408775_408775 ; 
   reg __408775_408775;
   reg _408776_408776 ; 
   reg __408776_408776;
   reg _408777_408777 ; 
   reg __408777_408777;
   reg _408778_408778 ; 
   reg __408778_408778;
   reg _408779_408779 ; 
   reg __408779_408779;
   reg _408780_408780 ; 
   reg __408780_408780;
   reg _408781_408781 ; 
   reg __408781_408781;
   reg _408782_408782 ; 
   reg __408782_408782;
   reg _408783_408783 ; 
   reg __408783_408783;
   reg _408784_408784 ; 
   reg __408784_408784;
   reg _408785_408785 ; 
   reg __408785_408785;
   reg _408786_408786 ; 
   reg __408786_408786;
   reg _408787_408787 ; 
   reg __408787_408787;
   reg _408788_408788 ; 
   reg __408788_408788;
   reg _408789_408789 ; 
   reg __408789_408789;
   reg _408790_408790 ; 
   reg __408790_408790;
   reg _408791_408791 ; 
   reg __408791_408791;
   reg _408792_408792 ; 
   reg __408792_408792;
   reg _408793_408793 ; 
   reg __408793_408793;
   reg _408794_408794 ; 
   reg __408794_408794;
   reg _408795_408795 ; 
   reg __408795_408795;
   reg _408796_408796 ; 
   reg __408796_408796;
   reg _408797_408797 ; 
   reg __408797_408797;
   reg _408798_408798 ; 
   reg __408798_408798;
   reg _408799_408799 ; 
   reg __408799_408799;
   reg _408800_408800 ; 
   reg __408800_408800;
   reg _408801_408801 ; 
   reg __408801_408801;
   reg _408802_408802 ; 
   reg __408802_408802;
   reg _408803_408803 ; 
   reg __408803_408803;
   reg _408804_408804 ; 
   reg __408804_408804;
   reg _408805_408805 ; 
   reg __408805_408805;
   reg _408806_408806 ; 
   reg __408806_408806;
   reg _408807_408807 ; 
   reg __408807_408807;
   reg _408808_408808 ; 
   reg __408808_408808;
   reg _408809_408809 ; 
   reg __408809_408809;
   reg _408810_408810 ; 
   reg __408810_408810;
   reg _408811_408811 ; 
   reg __408811_408811;
   reg _408812_408812 ; 
   reg __408812_408812;
   reg _408813_408813 ; 
   reg __408813_408813;
   reg _408814_408814 ; 
   reg __408814_408814;
   reg _408815_408815 ; 
   reg __408815_408815;
   reg _408816_408816 ; 
   reg __408816_408816;
   reg _408817_408817 ; 
   reg __408817_408817;
   reg _408818_408818 ; 
   reg __408818_408818;
   reg _408819_408819 ; 
   reg __408819_408819;
   reg _408820_408820 ; 
   reg __408820_408820;
   reg _408821_408821 ; 
   reg __408821_408821;
   reg _408822_408822 ; 
   reg __408822_408822;
   reg _408823_408823 ; 
   reg __408823_408823;
   reg _408824_408824 ; 
   reg __408824_408824;
   reg _408825_408825 ; 
   reg __408825_408825;
   reg _408826_408826 ; 
   reg __408826_408826;
   reg _408827_408827 ; 
   reg __408827_408827;
   reg _408828_408828 ; 
   reg __408828_408828;
   reg _408829_408829 ; 
   reg __408829_408829;
   reg _408830_408830 ; 
   reg __408830_408830;
   reg _408831_408831 ; 
   reg __408831_408831;
   reg _408832_408832 ; 
   reg __408832_408832;
   reg _408833_408833 ; 
   reg __408833_408833;
   reg _408834_408834 ; 
   reg __408834_408834;
   reg _408835_408835 ; 
   reg __408835_408835;
   reg _408836_408836 ; 
   reg __408836_408836;
   reg _408837_408837 ; 
   reg __408837_408837;
   reg _408838_408838 ; 
   reg __408838_408838;
   reg _408839_408839 ; 
   reg __408839_408839;
   reg _408840_408840 ; 
   reg __408840_408840;
   reg _408841_408841 ; 
   reg __408841_408841;
   reg _408842_408842 ; 
   reg __408842_408842;
   reg _408843_408843 ; 
   reg __408843_408843;
   reg _408844_408844 ; 
   reg __408844_408844;
   reg _408845_408845 ; 
   reg __408845_408845;
   reg _408846_408846 ; 
   reg __408846_408846;
   reg _408847_408847 ; 
   reg __408847_408847;
   reg _408848_408848 ; 
   reg __408848_408848;
   reg _408849_408849 ; 
   reg __408849_408849;
   reg _408850_408850 ; 
   reg __408850_408850;
   reg _408851_408851 ; 
   reg __408851_408851;
   reg _408852_408852 ; 
   reg __408852_408852;
   reg _408853_408853 ; 
   reg __408853_408853;
   reg _408854_408854 ; 
   reg __408854_408854;
   reg _408855_408855 ; 
   reg __408855_408855;
   reg _408856_408856 ; 
   reg __408856_408856;
   reg _408857_408857 ; 
   reg __408857_408857;
   reg _408858_408858 ; 
   reg __408858_408858;
   reg _408859_408859 ; 
   reg __408859_408859;
   reg _408860_408860 ; 
   reg __408860_408860;
   reg _408861_408861 ; 
   reg __408861_408861;
   reg _408862_408862 ; 
   reg __408862_408862;
   reg _408863_408863 ; 
   reg __408863_408863;
   reg _408864_408864 ; 
   reg __408864_408864;
   reg _408865_408865 ; 
   reg __408865_408865;
   reg _408866_408866 ; 
   reg __408866_408866;
   reg _408867_408867 ; 
   reg __408867_408867;
   reg _408868_408868 ; 
   reg __408868_408868;
   reg _408869_408869 ; 
   reg __408869_408869;
   reg _408870_408870 ; 
   reg __408870_408870;
   reg _408871_408871 ; 
   reg __408871_408871;
   reg _408872_408872 ; 
   reg __408872_408872;
   reg _408873_408873 ; 
   reg __408873_408873;
   reg _408874_408874 ; 
   reg __408874_408874;
   reg _408875_408875 ; 
   reg __408875_408875;
   reg _408876_408876 ; 
   reg __408876_408876;
   reg _408877_408877 ; 
   reg __408877_408877;
   reg _408878_408878 ; 
   reg __408878_408878;
   reg _408879_408879 ; 
   reg __408879_408879;
   reg _408880_408880 ; 
   reg __408880_408880;
   reg _408881_408881 ; 
   reg __408881_408881;
   reg _408882_408882 ; 
   reg __408882_408882;
   reg _408883_408883 ; 
   reg __408883_408883;
   reg _408884_408884 ; 
   reg __408884_408884;
   reg _408885_408885 ; 
   reg __408885_408885;
   reg _408886_408886 ; 
   reg __408886_408886;
   reg _408887_408887 ; 
   reg __408887_408887;
   reg _408888_408888 ; 
   reg __408888_408888;
   reg _408889_408889 ; 
   reg __408889_408889;
   reg _408890_408890 ; 
   reg __408890_408890;
   reg _408891_408891 ; 
   reg __408891_408891;
   reg _408892_408892 ; 
   reg __408892_408892;
   reg _408893_408893 ; 
   reg __408893_408893;
   reg _408894_408894 ; 
   reg __408894_408894;
   reg _408895_408895 ; 
   reg __408895_408895;
   reg _408896_408896 ; 
   reg __408896_408896;
   reg _408897_408897 ; 
   reg __408897_408897;
   reg _408898_408898 ; 
   reg __408898_408898;
   reg _408899_408899 ; 
   reg __408899_408899;
   reg _408900_408900 ; 
   reg __408900_408900;
   reg _408901_408901 ; 
   reg __408901_408901;
   reg _408902_408902 ; 
   reg __408902_408902;
   reg _408903_408903 ; 
   reg __408903_408903;
   reg _408904_408904 ; 
   reg __408904_408904;
   reg _408905_408905 ; 
   reg __408905_408905;
   reg _408906_408906 ; 
   reg __408906_408906;
   reg _408907_408907 ; 
   reg __408907_408907;
   reg _408908_408908 ; 
   reg __408908_408908;
   reg _408909_408909 ; 
   reg __408909_408909;
   reg _408910_408910 ; 
   reg __408910_408910;
   reg _408911_408911 ; 
   reg __408911_408911;
   reg _408912_408912 ; 
   reg __408912_408912;
   reg _408913_408913 ; 
   reg __408913_408913;
   reg _408914_408914 ; 
   reg __408914_408914;
   reg _408915_408915 ; 
   reg __408915_408915;
   reg _408916_408916 ; 
   reg __408916_408916;
   reg _408917_408917 ; 
   reg __408917_408917;
   reg _408918_408918 ; 
   reg __408918_408918;
   reg _408919_408919 ; 
   reg __408919_408919;
   reg _408920_408920 ; 
   reg __408920_408920;
   reg _408921_408921 ; 
   reg __408921_408921;
   reg _408922_408922 ; 
   reg __408922_408922;
   reg _408923_408923 ; 
   reg __408923_408923;
   reg _408924_408924 ; 
   reg __408924_408924;
   reg _408925_408925 ; 
   reg __408925_408925;
   reg _408926_408926 ; 
   reg __408926_408926;
   reg _408927_408927 ; 
   reg __408927_408927;
   reg _408928_408928 ; 
   reg __408928_408928;
   reg _408929_408929 ; 
   reg __408929_408929;
   reg _408930_408930 ; 
   reg __408930_408930;
   reg _408931_408931 ; 
   reg __408931_408931;
   reg _408932_408932 ; 
   reg __408932_408932;
   reg _408933_408933 ; 
   reg __408933_408933;
   reg _408934_408934 ; 
   reg __408934_408934;
   reg _408935_408935 ; 
   reg __408935_408935;
   reg _408936_408936 ; 
   reg __408936_408936;
   reg _408937_408937 ; 
   reg __408937_408937;
   reg _408938_408938 ; 
   reg __408938_408938;
   reg _408939_408939 ; 
   reg __408939_408939;
   reg _408940_408940 ; 
   reg __408940_408940;
   reg _408941_408941 ; 
   reg __408941_408941;
   reg _408942_408942 ; 
   reg __408942_408942;
   reg _408943_408943 ; 
   reg __408943_408943;
   reg _408944_408944 ; 
   reg __408944_408944;
   reg _408945_408945 ; 
   reg __408945_408945;
   reg _408946_408946 ; 
   reg __408946_408946;
   reg _408947_408947 ; 
   reg __408947_408947;
   reg _408948_408948 ; 
   reg __408948_408948;
   reg _408949_408949 ; 
   reg __408949_408949;
   reg _408950_408950 ; 
   reg __408950_408950;
   reg _408951_408951 ; 
   reg __408951_408951;
   reg _408952_408952 ; 
   reg __408952_408952;
   reg _408953_408953 ; 
   reg __408953_408953;
   reg _408954_408954 ; 
   reg __408954_408954;
   reg _408955_408955 ; 
   reg __408955_408955;
   reg _408956_408956 ; 
   reg __408956_408956;
   reg _408957_408957 ; 
   reg __408957_408957;
   reg _408958_408958 ; 
   reg __408958_408958;
   reg _408959_408959 ; 
   reg __408959_408959;
   reg _408960_408960 ; 
   reg __408960_408960;
   reg _408961_408961 ; 
   reg __408961_408961;
   reg _408962_408962 ; 
   reg __408962_408962;
   reg _408963_408963 ; 
   reg __408963_408963;
   reg _408964_408964 ; 
   reg __408964_408964;
   reg _408965_408965 ; 
   reg __408965_408965;
   reg _408966_408966 ; 
   reg __408966_408966;
   reg _408967_408967 ; 
   reg __408967_408967;
   reg _408968_408968 ; 
   reg __408968_408968;
   reg _408969_408969 ; 
   reg __408969_408969;
   reg _408970_408970 ; 
   reg __408970_408970;
   reg _408971_408971 ; 
   reg __408971_408971;
   reg _408972_408972 ; 
   reg __408972_408972;
   reg _408973_408973 ; 
   reg __408973_408973;
   reg _408974_408974 ; 
   reg __408974_408974;
   reg _408975_408975 ; 
   reg __408975_408975;
   reg _408976_408976 ; 
   reg __408976_408976;
   reg _408977_408977 ; 
   reg __408977_408977;
   reg _408978_408978 ; 
   reg __408978_408978;
   reg _408979_408979 ; 
   reg __408979_408979;
   reg _408980_408980 ; 
   reg __408980_408980;
   reg _408981_408981 ; 
   reg __408981_408981;
   reg _408982_408982 ; 
   reg __408982_408982;
   reg _408983_408983 ; 
   reg __408983_408983;
   reg _408984_408984 ; 
   reg __408984_408984;
   reg _408985_408985 ; 
   reg __408985_408985;
   reg _408986_408986 ; 
   reg __408986_408986;
   reg _408987_408987 ; 
   reg __408987_408987;
   reg _408988_408988 ; 
   reg __408988_408988;
   reg _408989_408989 ; 
   reg __408989_408989;
   reg _408990_408990 ; 
   reg __408990_408990;
   reg _408991_408991 ; 
   reg __408991_408991;
   reg _408992_408992 ; 
   reg __408992_408992;
   reg _408993_408993 ; 
   reg __408993_408993;
   reg _408994_408994 ; 
   reg __408994_408994;
   reg _408995_408995 ; 
   reg __408995_408995;
   reg _408996_408996 ; 
   reg __408996_408996;
   reg _408997_408997 ; 
   reg __408997_408997;
   reg _408998_408998 ; 
   reg __408998_408998;
   reg _408999_408999 ; 
   reg __408999_408999;
   reg _409000_409000 ; 
   reg __409000_409000;
   reg _409001_409001 ; 
   reg __409001_409001;
   reg _409002_409002 ; 
   reg __409002_409002;
   reg _409003_409003 ; 
   reg __409003_409003;
   reg _409004_409004 ; 
   reg __409004_409004;
   reg _409005_409005 ; 
   reg __409005_409005;
   reg _409006_409006 ; 
   reg __409006_409006;
   reg _409007_409007 ; 
   reg __409007_409007;
   reg _409008_409008 ; 
   reg __409008_409008;
   reg _409009_409009 ; 
   reg __409009_409009;
   reg _409010_409010 ; 
   reg __409010_409010;
   reg _409011_409011 ; 
   reg __409011_409011;
   reg _409012_409012 ; 
   reg __409012_409012;
   reg _409013_409013 ; 
   reg __409013_409013;
   reg _409014_409014 ; 
   reg __409014_409014;
   reg _409015_409015 ; 
   reg __409015_409015;
   reg _409016_409016 ; 
   reg __409016_409016;
   reg _409017_409017 ; 
   reg __409017_409017;
   reg _409018_409018 ; 
   reg __409018_409018;
   reg _409019_409019 ; 
   reg __409019_409019;
   reg _409020_409020 ; 
   reg __409020_409020;
   reg _409021_409021 ; 
   reg __409021_409021;
   reg _409022_409022 ; 
   reg __409022_409022;
   reg _409023_409023 ; 
   reg __409023_409023;
   reg _409024_409024 ; 
   reg __409024_409024;
   reg _409025_409025 ; 
   reg __409025_409025;
   reg _409026_409026 ; 
   reg __409026_409026;
   reg _409027_409027 ; 
   reg __409027_409027;
   reg _409028_409028 ; 
   reg __409028_409028;
   reg _409029_409029 ; 
   reg __409029_409029;
   reg _409030_409030 ; 
   reg __409030_409030;
   reg _409031_409031 ; 
   reg __409031_409031;
   reg _409032_409032 ; 
   reg __409032_409032;
   reg _409033_409033 ; 
   reg __409033_409033;
   reg _409034_409034 ; 
   reg __409034_409034;
   reg _409035_409035 ; 
   reg __409035_409035;
   reg _409036_409036 ; 
   reg __409036_409036;
   reg _409037_409037 ; 
   reg __409037_409037;
   reg _409038_409038 ; 
   reg __409038_409038;
   reg _409039_409039 ; 
   reg __409039_409039;
   reg _409040_409040 ; 
   reg __409040_409040;
   reg _409041_409041 ; 
   reg __409041_409041;
   reg _409042_409042 ; 
   reg __409042_409042;
   reg _409043_409043 ; 
   reg __409043_409043;
   reg _409044_409044 ; 
   reg __409044_409044;
   reg _409045_409045 ; 
   reg __409045_409045;
   reg _409046_409046 ; 
   reg __409046_409046;
   reg _409047_409047 ; 
   reg __409047_409047;
   reg _409048_409048 ; 
   reg __409048_409048;
   reg _409049_409049 ; 
   reg __409049_409049;
   reg _409050_409050 ; 
   reg __409050_409050;
   reg _409051_409051 ; 
   reg __409051_409051;
   reg _409052_409052 ; 
   reg __409052_409052;
   reg _409053_409053 ; 
   reg __409053_409053;
   reg _409054_409054 ; 
   reg __409054_409054;
   reg _409055_409055 ; 
   reg __409055_409055;
   reg _409056_409056 ; 
   reg __409056_409056;
   reg _409057_409057 ; 
   reg __409057_409057;
   reg _409058_409058 ; 
   reg __409058_409058;
   reg _409059_409059 ; 
   reg __409059_409059;
   reg _409060_409060 ; 
   reg __409060_409060;
   reg _409061_409061 ; 
   reg __409061_409061;
   reg _409062_409062 ; 
   reg __409062_409062;
   reg _409063_409063 ; 
   reg __409063_409063;
   reg _409064_409064 ; 
   reg __409064_409064;
   reg _409065_409065 ; 
   reg __409065_409065;
   reg _409066_409066 ; 
   reg __409066_409066;
   reg _409067_409067 ; 
   reg __409067_409067;
   reg _409068_409068 ; 
   reg __409068_409068;
   reg _409069_409069 ; 
   reg __409069_409069;
   reg _409070_409070 ; 
   reg __409070_409070;
   reg _409071_409071 ; 
   reg __409071_409071;
   reg _409072_409072 ; 
   reg __409072_409072;
   reg _409073_409073 ; 
   reg __409073_409073;
   reg _409074_409074 ; 
   reg __409074_409074;
   reg _409075_409075 ; 
   reg __409075_409075;
   reg _409076_409076 ; 
   reg __409076_409076;
   reg _409077_409077 ; 
   reg __409077_409077;
   reg _409078_409078 ; 
   reg __409078_409078;
   reg _409079_409079 ; 
   reg __409079_409079;
   reg _409080_409080 ; 
   reg __409080_409080;
   reg _409081_409081 ; 
   reg __409081_409081;
   reg _409082_409082 ; 
   reg __409082_409082;
   reg _409083_409083 ; 
   reg __409083_409083;
   reg _409084_409084 ; 
   reg __409084_409084;
   reg _409085_409085 ; 
   reg __409085_409085;
   reg _409086_409086 ; 
   reg __409086_409086;
   reg _409087_409087 ; 
   reg __409087_409087;
   reg _409088_409088 ; 
   reg __409088_409088;
   reg _409089_409089 ; 
   reg __409089_409089;
   reg _409090_409090 ; 
   reg __409090_409090;
   reg _409091_409091 ; 
   reg __409091_409091;
   reg _409092_409092 ; 
   reg __409092_409092;
   reg _409093_409093 ; 
   reg __409093_409093;
   reg _409094_409094 ; 
   reg __409094_409094;
   reg _409095_409095 ; 
   reg __409095_409095;
   reg _409096_409096 ; 
   reg __409096_409096;
   reg _409097_409097 ; 
   reg __409097_409097;
   reg _409098_409098 ; 
   reg __409098_409098;
   reg _409099_409099 ; 
   reg __409099_409099;
   reg _409100_409100 ; 
   reg __409100_409100;
   reg _409101_409101 ; 
   reg __409101_409101;
   reg _409102_409102 ; 
   reg __409102_409102;
   reg _409103_409103 ; 
   reg __409103_409103;
   reg _409104_409104 ; 
   reg __409104_409104;
   reg _409105_409105 ; 
   reg __409105_409105;
   reg _409106_409106 ; 
   reg __409106_409106;
   reg _409107_409107 ; 
   reg __409107_409107;
   reg _409108_409108 ; 
   reg __409108_409108;
   reg _409109_409109 ; 
   reg __409109_409109;
   reg _409110_409110 ; 
   reg __409110_409110;
   reg _409111_409111 ; 
   reg __409111_409111;
   reg _409112_409112 ; 
   reg __409112_409112;
   reg _409113_409113 ; 
   reg __409113_409113;
   reg _409114_409114 ; 
   reg __409114_409114;
   reg _409115_409115 ; 
   reg __409115_409115;
   reg _409116_409116 ; 
   reg __409116_409116;
   reg _409117_409117 ; 
   reg __409117_409117;
   reg _409118_409118 ; 
   reg __409118_409118;
   reg _409119_409119 ; 
   reg __409119_409119;
   reg _409120_409120 ; 
   reg __409120_409120;
   reg _409121_409121 ; 
   reg __409121_409121;
   reg _409122_409122 ; 
   reg __409122_409122;
   reg _409123_409123 ; 
   reg __409123_409123;
   reg _409124_409124 ; 
   reg __409124_409124;
   reg _409125_409125 ; 
   reg __409125_409125;
   reg _409126_409126 ; 
   reg __409126_409126;
   reg _409127_409127 ; 
   reg __409127_409127;
   reg _409128_409128 ; 
   reg __409128_409128;
   reg _409129_409129 ; 
   reg __409129_409129;
   reg _409130_409130 ; 
   reg __409130_409130;
   reg _409131_409131 ; 
   reg __409131_409131;
   reg _409132_409132 ; 
   reg __409132_409132;
   reg _409133_409133 ; 
   reg __409133_409133;
   reg _409134_409134 ; 
   reg __409134_409134;
   reg _409135_409135 ; 
   reg __409135_409135;
   reg _409136_409136 ; 
   reg __409136_409136;
   reg _409137_409137 ; 
   reg __409137_409137;
   reg _409138_409138 ; 
   reg __409138_409138;
   reg _409139_409139 ; 
   reg __409139_409139;
   reg _409140_409140 ; 
   reg __409140_409140;
   reg _409141_409141 ; 
   reg __409141_409141;
   reg _409142_409142 ; 
   reg __409142_409142;
   reg _409143_409143 ; 
   reg __409143_409143;
   reg _409144_409144 ; 
   reg __409144_409144;
   reg _409145_409145 ; 
   reg __409145_409145;
   reg _409146_409146 ; 
   reg __409146_409146;
   reg _409147_409147 ; 
   reg __409147_409147;
   reg _409148_409148 ; 
   reg __409148_409148;
   reg _409149_409149 ; 
   reg __409149_409149;
   reg _409150_409150 ; 
   reg __409150_409150;
   reg _409151_409151 ; 
   reg __409151_409151;
   reg _409152_409152 ; 
   reg __409152_409152;
   reg _409153_409153 ; 
   reg __409153_409153;
   reg _409154_409154 ; 
   reg __409154_409154;
   reg _409155_409155 ; 
   reg __409155_409155;
   reg _409156_409156 ; 
   reg __409156_409156;
   reg _409157_409157 ; 
   reg __409157_409157;
   reg _409158_409158 ; 
   reg __409158_409158;
   reg _409159_409159 ; 
   reg __409159_409159;
   reg _409160_409160 ; 
   reg __409160_409160;
   reg _409161_409161 ; 
   reg __409161_409161;
   reg _409162_409162 ; 
   reg __409162_409162;
   reg _409163_409163 ; 
   reg __409163_409163;
   reg _409164_409164 ; 
   reg __409164_409164;
   reg _409165_409165 ; 
   reg __409165_409165;
   reg _409166_409166 ; 
   reg __409166_409166;
   reg _409167_409167 ; 
   reg __409167_409167;
   reg _409168_409168 ; 
   reg __409168_409168;
   reg _409169_409169 ; 
   reg __409169_409169;
   reg _409170_409170 ; 
   reg __409170_409170;
   reg _409171_409171 ; 
   reg __409171_409171;
   reg _409172_409172 ; 
   reg __409172_409172;
   reg _409173_409173 ; 
   reg __409173_409173;
   reg _409174_409174 ; 
   reg __409174_409174;
   reg _409175_409175 ; 
   reg __409175_409175;
   reg _409176_409176 ; 
   reg __409176_409176;
   reg _409177_409177 ; 
   reg __409177_409177;
   reg _409178_409178 ; 
   reg __409178_409178;
   reg _409179_409179 ; 
   reg __409179_409179;
   reg _409180_409180 ; 
   reg __409180_409180;
   reg _409181_409181 ; 
   reg __409181_409181;
   reg _409182_409182 ; 
   reg __409182_409182;
   reg _409183_409183 ; 
   reg __409183_409183;
   reg _409184_409184 ; 
   reg __409184_409184;
   reg _409185_409185 ; 
   reg __409185_409185;
   reg _409186_409186 ; 
   reg __409186_409186;
   reg _409187_409187 ; 
   reg __409187_409187;
   reg _409188_409188 ; 
   reg __409188_409188;
   reg _409189_409189 ; 
   reg __409189_409189;
   reg _409190_409190 ; 
   reg __409190_409190;
   reg _409191_409191 ; 
   reg __409191_409191;
   reg _409192_409192 ; 
   reg __409192_409192;
   reg _409193_409193 ; 
   reg __409193_409193;
   reg _409194_409194 ; 
   reg __409194_409194;
   reg _409195_409195 ; 
   reg __409195_409195;
   reg _409196_409196 ; 
   reg __409196_409196;
   reg _409197_409197 ; 
   reg __409197_409197;
   reg _409198_409198 ; 
   reg __409198_409198;
   reg _409199_409199 ; 
   reg __409199_409199;
   reg _409200_409200 ; 
   reg __409200_409200;
   reg _409201_409201 ; 
   reg __409201_409201;
   reg _409202_409202 ; 
   reg __409202_409202;
   reg _409203_409203 ; 
   reg __409203_409203;
   reg _409204_409204 ; 
   reg __409204_409204;
   reg _409205_409205 ; 
   reg __409205_409205;
   reg _409206_409206 ; 
   reg __409206_409206;
   reg _409207_409207 ; 
   reg __409207_409207;
   reg _409208_409208 ; 
   reg __409208_409208;
   reg _409209_409209 ; 
   reg __409209_409209;
   reg _409210_409210 ; 
   reg __409210_409210;
   reg _409211_409211 ; 
   reg __409211_409211;
   reg _409212_409212 ; 
   reg __409212_409212;
   reg _409213_409213 ; 
   reg __409213_409213;
   reg _409214_409214 ; 
   reg __409214_409214;
   reg _409215_409215 ; 
   reg __409215_409215;
   reg _409216_409216 ; 
   reg __409216_409216;
   reg _409217_409217 ; 
   reg __409217_409217;
   reg _409218_409218 ; 
   reg __409218_409218;
   reg _409219_409219 ; 
   reg __409219_409219;
   reg _409220_409220 ; 
   reg __409220_409220;
   reg _409221_409221 ; 
   reg __409221_409221;
   reg _409222_409222 ; 
   reg __409222_409222;
   reg _409223_409223 ; 
   reg __409223_409223;
   reg _409224_409224 ; 
   reg __409224_409224;
   reg _409225_409225 ; 
   reg __409225_409225;
   reg _409226_409226 ; 
   reg __409226_409226;
   reg _409227_409227 ; 
   reg __409227_409227;
   reg _409228_409228 ; 
   reg __409228_409228;
   reg _409229_409229 ; 
   reg __409229_409229;
   reg _409230_409230 ; 
   reg __409230_409230;
   reg _409231_409231 ; 
   reg __409231_409231;
   reg _409232_409232 ; 
   reg __409232_409232;
   reg _409233_409233 ; 
   reg __409233_409233;
   reg _409234_409234 ; 
   reg __409234_409234;
   reg _409235_409235 ; 
   reg __409235_409235;
   reg _409236_409236 ; 
   reg __409236_409236;
   reg _409237_409237 ; 
   reg __409237_409237;
   reg _409238_409238 ; 
   reg __409238_409238;
   reg _409239_409239 ; 
   reg __409239_409239;
   reg _409240_409240 ; 
   reg __409240_409240;
   reg _409241_409241 ; 
   reg __409241_409241;
   reg _409242_409242 ; 
   reg __409242_409242;
   reg _409243_409243 ; 
   reg __409243_409243;
   reg _409244_409244 ; 
   reg __409244_409244;
   reg _409245_409245 ; 
   reg __409245_409245;
   reg _409246_409246 ; 
   reg __409246_409246;
   reg _409247_409247 ; 
   reg __409247_409247;
   reg _409248_409248 ; 
   reg __409248_409248;
   reg _409249_409249 ; 
   reg __409249_409249;
   reg _409250_409250 ; 
   reg __409250_409250;
   reg _409251_409251 ; 
   reg __409251_409251;
   reg _409252_409252 ; 
   reg __409252_409252;
   reg _409253_409253 ; 
   reg __409253_409253;
   reg _409254_409254 ; 
   reg __409254_409254;
   reg _409255_409255 ; 
   reg __409255_409255;
   reg _409256_409256 ; 
   reg __409256_409256;
   reg _409257_409257 ; 
   reg __409257_409257;
   reg _409258_409258 ; 
   reg __409258_409258;
   reg _409259_409259 ; 
   reg __409259_409259;
   reg _409260_409260 ; 
   reg __409260_409260;
   reg _409261_409261 ; 
   reg __409261_409261;
   reg _409262_409262 ; 
   reg __409262_409262;
   reg _409263_409263 ; 
   reg __409263_409263;
   reg _409264_409264 ; 
   reg __409264_409264;
   reg _409265_409265 ; 
   reg __409265_409265;
   reg _409266_409266 ; 
   reg __409266_409266;
   reg _409267_409267 ; 
   reg __409267_409267;
   reg _409268_409268 ; 
   reg __409268_409268;
   reg _409269_409269 ; 
   reg __409269_409269;
   reg _409270_409270 ; 
   reg __409270_409270;
   reg _409271_409271 ; 
   reg __409271_409271;
   reg _409272_409272 ; 
   reg __409272_409272;
   reg _409273_409273 ; 
   reg __409273_409273;
   reg _409274_409274 ; 
   reg __409274_409274;
   reg _409275_409275 ; 
   reg __409275_409275;
   reg _409276_409276 ; 
   reg __409276_409276;
   reg _409277_409277 ; 
   reg __409277_409277;
   reg _409278_409278 ; 
   reg __409278_409278;
   reg _409279_409279 ; 
   reg __409279_409279;
   reg _409280_409280 ; 
   reg __409280_409280;
   reg _409281_409281 ; 
   reg __409281_409281;
   reg _409282_409282 ; 
   reg __409282_409282;
   reg _409283_409283 ; 
   reg __409283_409283;
   reg _409284_409284 ; 
   reg __409284_409284;
   reg _409285_409285 ; 
   reg __409285_409285;
   reg _409286_409286 ; 
   reg __409286_409286;
   reg _409287_409287 ; 
   reg __409287_409287;
   reg _409288_409288 ; 
   reg __409288_409288;
   reg _409289_409289 ; 
   reg __409289_409289;
   reg _409290_409290 ; 
   reg __409290_409290;
   reg _409291_409291 ; 
   reg __409291_409291;
   reg _409292_409292 ; 
   reg __409292_409292;
   reg _409293_409293 ; 
   reg __409293_409293;
   reg _409294_409294 ; 
   reg __409294_409294;
   reg _409295_409295 ; 
   reg __409295_409295;
   reg _409296_409296 ; 
   reg __409296_409296;
   reg _409297_409297 ; 
   reg __409297_409297;
   reg _409298_409298 ; 
   reg __409298_409298;
   reg _409299_409299 ; 
   reg __409299_409299;
   reg _409300_409300 ; 
   reg __409300_409300;
   reg _409301_409301 ; 
   reg __409301_409301;
   reg _409302_409302 ; 
   reg __409302_409302;
   reg _409303_409303 ; 
   reg __409303_409303;
   reg _409304_409304 ; 
   reg __409304_409304;
   reg _409305_409305 ; 
   reg __409305_409305;
   reg _409306_409306 ; 
   reg __409306_409306;
   reg _409307_409307 ; 
   reg __409307_409307;
   reg _409308_409308 ; 
   reg __409308_409308;
   reg _409309_409309 ; 
   reg __409309_409309;
   reg _409310_409310 ; 
   reg __409310_409310;
   reg _409311_409311 ; 
   reg __409311_409311;
   reg _409312_409312 ; 
   reg __409312_409312;
   reg _409313_409313 ; 
   reg __409313_409313;
   reg _409314_409314 ; 
   reg __409314_409314;
   reg _409315_409315 ; 
   reg __409315_409315;
   reg _409316_409316 ; 
   reg __409316_409316;
   reg _409317_409317 ; 
   reg __409317_409317;
   reg _409318_409318 ; 
   reg __409318_409318;
   reg _409319_409319 ; 
   reg __409319_409319;
   reg _409320_409320 ; 
   reg __409320_409320;
   reg _409321_409321 ; 
   reg __409321_409321;
   reg _409322_409322 ; 
   reg __409322_409322;
   reg _409323_409323 ; 
   reg __409323_409323;
   reg _409324_409324 ; 
   reg __409324_409324;
   reg _409325_409325 ; 
   reg __409325_409325;
   reg _409326_409326 ; 
   reg __409326_409326;
   reg _409327_409327 ; 
   reg __409327_409327;
   reg _409328_409328 ; 
   reg __409328_409328;
   reg _409329_409329 ; 
   reg __409329_409329;
   reg _409330_409330 ; 
   reg __409330_409330;
   reg _409331_409331 ; 
   reg __409331_409331;
   reg _409332_409332 ; 
   reg __409332_409332;
   reg _409333_409333 ; 
   reg __409333_409333;
   reg _409334_409334 ; 
   reg __409334_409334;
   reg _409335_409335 ; 
   reg __409335_409335;
   reg _409336_409336 ; 
   reg __409336_409336;
   reg _409337_409337 ; 
   reg __409337_409337;
   reg _409338_409338 ; 
   reg __409338_409338;
   reg _409339_409339 ; 
   reg __409339_409339;
   reg _409340_409340 ; 
   reg __409340_409340;
   reg _409341_409341 ; 
   reg __409341_409341;
   reg _409342_409342 ; 
   reg __409342_409342;
   reg _409343_409343 ; 
   reg __409343_409343;
   reg _409344_409344 ; 
   reg __409344_409344;
   reg _409345_409345 ; 
   reg __409345_409345;
   reg _409346_409346 ; 
   reg __409346_409346;
   reg _409347_409347 ; 
   reg __409347_409347;
   reg _409348_409348 ; 
   reg __409348_409348;
   reg _409349_409349 ; 
   reg __409349_409349;
   reg _409350_409350 ; 
   reg __409350_409350;
   reg _409351_409351 ; 
   reg __409351_409351;
   reg _409352_409352 ; 
   reg __409352_409352;
   reg _409353_409353 ; 
   reg __409353_409353;
   reg _409354_409354 ; 
   reg __409354_409354;
   reg _409355_409355 ; 
   reg __409355_409355;
   reg _409356_409356 ; 
   reg __409356_409356;
   reg _409357_409357 ; 
   reg __409357_409357;
   reg _409358_409358 ; 
   reg __409358_409358;
   reg _409359_409359 ; 
   reg __409359_409359;
   reg _409360_409360 ; 
   reg __409360_409360;
   reg _409361_409361 ; 
   reg __409361_409361;
   reg _409362_409362 ; 
   reg __409362_409362;
   reg _409363_409363 ; 
   reg __409363_409363;
   reg _409364_409364 ; 
   reg __409364_409364;
   reg _409365_409365 ; 
   reg __409365_409365;
   reg _409366_409366 ; 
   reg __409366_409366;
   reg _409367_409367 ; 
   reg __409367_409367;
   reg _409368_409368 ; 
   reg __409368_409368;
   reg _409369_409369 ; 
   reg __409369_409369;
   reg _409370_409370 ; 
   reg __409370_409370;
   reg _409371_409371 ; 
   reg __409371_409371;
   reg _409372_409372 ; 
   reg __409372_409372;
   reg _409373_409373 ; 
   reg __409373_409373;
   reg _409374_409374 ; 
   reg __409374_409374;
   reg _409375_409375 ; 
   reg __409375_409375;
   reg _409376_409376 ; 
   reg __409376_409376;
   reg _409377_409377 ; 
   reg __409377_409377;
   reg _409378_409378 ; 
   reg __409378_409378;
   reg _409379_409379 ; 
   reg __409379_409379;
   reg _409380_409380 ; 
   reg __409380_409380;
   reg _409381_409381 ; 
   reg __409381_409381;
   reg _409382_409382 ; 
   reg __409382_409382;
   reg _409383_409383 ; 
   reg __409383_409383;
   reg _409384_409384 ; 
   reg __409384_409384;
   reg _409385_409385 ; 
   reg __409385_409385;
   reg _409386_409386 ; 
   reg __409386_409386;
   reg _409387_409387 ; 
   reg __409387_409387;
   reg _409388_409388 ; 
   reg __409388_409388;
   reg _409389_409389 ; 
   reg __409389_409389;
   reg _409390_409390 ; 
   reg __409390_409390;
   reg _409391_409391 ; 
   reg __409391_409391;
   reg _409392_409392 ; 
   reg __409392_409392;
   reg _409393_409393 ; 
   reg __409393_409393;
   reg _409394_409394 ; 
   reg __409394_409394;
   reg _409395_409395 ; 
   reg __409395_409395;
   reg _409396_409396 ; 
   reg __409396_409396;
   reg _409397_409397 ; 
   reg __409397_409397;
   reg _409398_409398 ; 
   reg __409398_409398;
   reg _409399_409399 ; 
   reg __409399_409399;
   reg _409400_409400 ; 
   reg __409400_409400;
   reg _409401_409401 ; 
   reg __409401_409401;
   reg _409402_409402 ; 
   reg __409402_409402;
   reg _409403_409403 ; 
   reg __409403_409403;
   reg _409404_409404 ; 
   reg __409404_409404;
   reg _409405_409405 ; 
   reg __409405_409405;
   reg _409406_409406 ; 
   reg __409406_409406;
   reg _409407_409407 ; 
   reg __409407_409407;
   reg _409408_409408 ; 
   reg __409408_409408;
   reg _409409_409409 ; 
   reg __409409_409409;
   reg _409410_409410 ; 
   reg __409410_409410;
   reg _409411_409411 ; 
   reg __409411_409411;
   reg _409412_409412 ; 
   reg __409412_409412;
   reg _409413_409413 ; 
   reg __409413_409413;
   reg _409414_409414 ; 
   reg __409414_409414;
   reg _409415_409415 ; 
   reg __409415_409415;
   reg _409416_409416 ; 
   reg __409416_409416;
   reg _409417_409417 ; 
   reg __409417_409417;
   reg _409418_409418 ; 
   reg __409418_409418;
   reg _409419_409419 ; 
   reg __409419_409419;
   reg _409420_409420 ; 
   reg __409420_409420;
   reg _409421_409421 ; 
   reg __409421_409421;
   reg _409422_409422 ; 
   reg __409422_409422;
   reg _409423_409423 ; 
   reg __409423_409423;
   reg _409424_409424 ; 
   reg __409424_409424;
   reg _409425_409425 ; 
   reg __409425_409425;
   reg _409426_409426 ; 
   reg __409426_409426;
   reg _409427_409427 ; 
   reg __409427_409427;
   reg _409428_409428 ; 
   reg __409428_409428;
   reg _409429_409429 ; 
   reg __409429_409429;
   reg _409430_409430 ; 
   reg __409430_409430;
   reg _409431_409431 ; 
   reg __409431_409431;
   reg _409432_409432 ; 
   reg __409432_409432;
   reg _409433_409433 ; 
   reg __409433_409433;
   reg _409434_409434 ; 
   reg __409434_409434;
   reg _409435_409435 ; 
   reg __409435_409435;
   reg _409436_409436 ; 
   reg __409436_409436;
   reg _409437_409437 ; 
   reg __409437_409437;
   reg _409438_409438 ; 
   reg __409438_409438;
   reg _409439_409439 ; 
   reg __409439_409439;
   reg _409440_409440 ; 
   reg __409440_409440;
   reg _409441_409441 ; 
   reg __409441_409441;
   reg _409442_409442 ; 
   reg __409442_409442;
   reg _409443_409443 ; 
   reg __409443_409443;
   reg _409444_409444 ; 
   reg __409444_409444;
   reg _409445_409445 ; 
   reg __409445_409445;
   reg _409446_409446 ; 
   reg __409446_409446;
   reg _409447_409447 ; 
   reg __409447_409447;
   reg _409448_409448 ; 
   reg __409448_409448;
   reg _409449_409449 ; 
   reg __409449_409449;
   reg _409450_409450 ; 
   reg __409450_409450;
   reg _409451_409451 ; 
   reg __409451_409451;
   reg _409452_409452 ; 
   reg __409452_409452;
   reg _409453_409453 ; 
   reg __409453_409453;
   reg _409454_409454 ; 
   reg __409454_409454;
   reg _409455_409455 ; 
   reg __409455_409455;
   reg _409456_409456 ; 
   reg __409456_409456;
   reg _409457_409457 ; 
   reg __409457_409457;
   reg _409458_409458 ; 
   reg __409458_409458;
   reg _409459_409459 ; 
   reg __409459_409459;
   reg _409460_409460 ; 
   reg __409460_409460;
   reg _409461_409461 ; 
   reg __409461_409461;
   reg _409462_409462 ; 
   reg __409462_409462;
   reg _409463_409463 ; 
   reg __409463_409463;
   reg _409464_409464 ; 
   reg __409464_409464;
   reg _409465_409465 ; 
   reg __409465_409465;
   reg _409466_409466 ; 
   reg __409466_409466;
   reg _409467_409467 ; 
   reg __409467_409467;
   reg _409468_409468 ; 
   reg __409468_409468;
   reg _409469_409469 ; 
   reg __409469_409469;
   reg _409470_409470 ; 
   reg __409470_409470;
   reg _409471_409471 ; 
   reg __409471_409471;
   reg _409472_409472 ; 
   reg __409472_409472;
   reg _409473_409473 ; 
   reg __409473_409473;
   reg _409474_409474 ; 
   reg __409474_409474;
   reg _409475_409475 ; 
   reg __409475_409475;
   reg _409476_409476 ; 
   reg __409476_409476;
   reg _409477_409477 ; 
   reg __409477_409477;
   reg _409478_409478 ; 
   reg __409478_409478;
   reg _409479_409479 ; 
   reg __409479_409479;
   reg _409480_409480 ; 
   reg __409480_409480;
   reg _409481_409481 ; 
   reg __409481_409481;
   reg _409482_409482 ; 
   reg __409482_409482;
   reg _409483_409483 ; 
   reg __409483_409483;
   reg _409484_409484 ; 
   reg __409484_409484;
   reg _409485_409485 ; 
   reg __409485_409485;
   reg _409486_409486 ; 
   reg __409486_409486;
   reg _409487_409487 ; 
   reg __409487_409487;
   reg _409488_409488 ; 
   reg __409488_409488;
   reg _409489_409489 ; 
   reg __409489_409489;
   reg _409490_409490 ; 
   reg __409490_409490;
   reg _409491_409491 ; 
   reg __409491_409491;
   reg _409492_409492 ; 
   reg __409492_409492;
   reg _409493_409493 ; 
   reg __409493_409493;
   reg _409494_409494 ; 
   reg __409494_409494;
   reg _409495_409495 ; 
   reg __409495_409495;
   reg _409496_409496 ; 
   reg __409496_409496;
   reg _409497_409497 ; 
   reg __409497_409497;
   reg _409498_409498 ; 
   reg __409498_409498;
   reg _409499_409499 ; 
   reg __409499_409499;
   reg _409500_409500 ; 
   reg __409500_409500;
   reg _409501_409501 ; 
   reg __409501_409501;
   reg _409502_409502 ; 
   reg __409502_409502;
   reg _409503_409503 ; 
   reg __409503_409503;
   reg _409504_409504 ; 
   reg __409504_409504;
   reg _409505_409505 ; 
   reg __409505_409505;
   reg _409506_409506 ; 
   reg __409506_409506;
   reg _409507_409507 ; 
   reg __409507_409507;
   reg _409508_409508 ; 
   reg __409508_409508;
   reg _409509_409509 ; 
   reg __409509_409509;
   reg _409510_409510 ; 
   reg __409510_409510;
   reg _409511_409511 ; 
   reg __409511_409511;
   reg _409512_409512 ; 
   reg __409512_409512;
   reg _409513_409513 ; 
   reg __409513_409513;
   reg _409514_409514 ; 
   reg __409514_409514;
   reg _409515_409515 ; 
   reg __409515_409515;
   reg _409516_409516 ; 
   reg __409516_409516;
   reg _409517_409517 ; 
   reg __409517_409517;
   reg _409518_409518 ; 
   reg __409518_409518;
   reg _409519_409519 ; 
   reg __409519_409519;
   reg _409520_409520 ; 
   reg __409520_409520;
   reg _409521_409521 ; 
   reg __409521_409521;
   reg _409522_409522 ; 
   reg __409522_409522;
   reg _409523_409523 ; 
   reg __409523_409523;
   reg _409524_409524 ; 
   reg __409524_409524;
   reg _409525_409525 ; 
   reg __409525_409525;
   reg _409526_409526 ; 
   reg __409526_409526;
   reg _409527_409527 ; 
   reg __409527_409527;
   reg _409528_409528 ; 
   reg __409528_409528;
   reg _409529_409529 ; 
   reg __409529_409529;
   reg _409530_409530 ; 
   reg __409530_409530;
   reg _409531_409531 ; 
   reg __409531_409531;
   reg _409532_409532 ; 
   reg __409532_409532;
   reg _409533_409533 ; 
   reg __409533_409533;
   reg _409534_409534 ; 
   reg __409534_409534;
   reg _409535_409535 ; 
   reg __409535_409535;
   reg _409536_409536 ; 
   reg __409536_409536;
   reg _409537_409537 ; 
   reg __409537_409537;
   reg _409538_409538 ; 
   reg __409538_409538;
   reg _409539_409539 ; 
   reg __409539_409539;
   reg _409540_409540 ; 
   reg __409540_409540;
   reg _409541_409541 ; 
   reg __409541_409541;
   reg _409542_409542 ; 
   reg __409542_409542;
   reg _409543_409543 ; 
   reg __409543_409543;
   reg _409544_409544 ; 
   reg __409544_409544;
   reg _409545_409545 ; 
   reg __409545_409545;
   reg _409546_409546 ; 
   reg __409546_409546;
   reg _409547_409547 ; 
   reg __409547_409547;
   reg _409548_409548 ; 
   reg __409548_409548;
   reg _409549_409549 ; 
   reg __409549_409549;
   reg _409550_409550 ; 
   reg __409550_409550;
   reg _409551_409551 ; 
   reg __409551_409551;
   reg _409552_409552 ; 
   reg __409552_409552;
   reg _409553_409553 ; 
   reg __409553_409553;
   reg _409554_409554 ; 
   reg __409554_409554;
   reg _409555_409555 ; 
   reg __409555_409555;
   reg _409556_409556 ; 
   reg __409556_409556;
   reg _409557_409557 ; 
   reg __409557_409557;
   reg _409558_409558 ; 
   reg __409558_409558;
   reg _409559_409559 ; 
   reg __409559_409559;
   reg _409560_409560 ; 
   reg __409560_409560;
   reg _409561_409561 ; 
   reg __409561_409561;
   reg _409562_409562 ; 
   reg __409562_409562;
   reg _409563_409563 ; 
   reg __409563_409563;
   reg _409564_409564 ; 
   reg __409564_409564;
   reg _409565_409565 ; 
   reg __409565_409565;
   reg _409566_409566 ; 
   reg __409566_409566;
   reg _409567_409567 ; 
   reg __409567_409567;
   reg _409568_409568 ; 
   reg __409568_409568;
   reg _409569_409569 ; 
   reg __409569_409569;
   reg _409570_409570 ; 
   reg __409570_409570;
   reg _409571_409571 ; 
   reg __409571_409571;
   reg _409572_409572 ; 
   reg __409572_409572;
   reg _409573_409573 ; 
   reg __409573_409573;
   reg _409574_409574 ; 
   reg __409574_409574;
   reg _409575_409575 ; 
   reg __409575_409575;
   reg _409576_409576 ; 
   reg __409576_409576;
   reg _409577_409577 ; 
   reg __409577_409577;
   reg _409578_409578 ; 
   reg __409578_409578;
   reg _409579_409579 ; 
   reg __409579_409579;
   reg _409580_409580 ; 
   reg __409580_409580;
   reg _409581_409581 ; 
   reg __409581_409581;
   reg _409582_409582 ; 
   reg __409582_409582;
   reg _409583_409583 ; 
   reg __409583_409583;
   reg _409584_409584 ; 
   reg __409584_409584;
   reg _409585_409585 ; 
   reg __409585_409585;
   reg _409586_409586 ; 
   reg __409586_409586;
   reg _409587_409587 ; 
   reg __409587_409587;
   reg _409588_409588 ; 
   reg __409588_409588;
   reg _409589_409589 ; 
   reg __409589_409589;
   reg _409590_409590 ; 
   reg __409590_409590;
   reg _409591_409591 ; 
   reg __409591_409591;
   reg _409592_409592 ; 
   reg __409592_409592;
   reg _409593_409593 ; 
   reg __409593_409593;
   reg _409594_409594 ; 
   reg __409594_409594;
   reg _409595_409595 ; 
   reg __409595_409595;
   reg _409596_409596 ; 
   reg __409596_409596;
   reg _409597_409597 ; 
   reg __409597_409597;
   reg _409598_409598 ; 
   reg __409598_409598;
   reg _409599_409599 ; 
   reg __409599_409599;
   reg _409600_409600 ; 
   reg __409600_409600;
   reg _409601_409601 ; 
   reg __409601_409601;
   reg _409602_409602 ; 
   reg __409602_409602;
   reg _409603_409603 ; 
   reg __409603_409603;
   reg _409604_409604 ; 
   reg __409604_409604;
   reg _409605_409605 ; 
   reg __409605_409605;
   reg _409606_409606 ; 
   reg __409606_409606;
   reg _409607_409607 ; 
   reg __409607_409607;
   reg _409608_409608 ; 
   reg __409608_409608;
   reg _409609_409609 ; 
   reg __409609_409609;
   reg _409610_409610 ; 
   reg __409610_409610;
   reg _409611_409611 ; 
   reg __409611_409611;
   reg _409612_409612 ; 
   reg __409612_409612;
   reg _409613_409613 ; 
   reg __409613_409613;
   reg _409614_409614 ; 
   reg __409614_409614;
   reg _409615_409615 ; 
   reg __409615_409615;
   reg _409616_409616 ; 
   reg __409616_409616;
   reg _409617_409617 ; 
   reg __409617_409617;
   reg _409618_409618 ; 
   reg __409618_409618;
   reg _409619_409619 ; 
   reg __409619_409619;
   reg _409620_409620 ; 
   reg __409620_409620;
   reg _409621_409621 ; 
   reg __409621_409621;
   reg _409622_409622 ; 
   reg __409622_409622;
   reg _409623_409623 ; 
   reg __409623_409623;
   reg _409624_409624 ; 
   reg __409624_409624;
   reg _409625_409625 ; 
   reg __409625_409625;
   reg _409626_409626 ; 
   reg __409626_409626;
   reg _409627_409627 ; 
   reg __409627_409627;
   reg _409628_409628 ; 
   reg __409628_409628;
   reg _409629_409629 ; 
   reg __409629_409629;
   reg _409630_409630 ; 
   reg __409630_409630;
   reg _409631_409631 ; 
   reg __409631_409631;
   reg _409632_409632 ; 
   reg __409632_409632;
   reg _409633_409633 ; 
   reg __409633_409633;
   reg _409634_409634 ; 
   reg __409634_409634;
   reg _409635_409635 ; 
   reg __409635_409635;
   reg _409636_409636 ; 
   reg __409636_409636;
   reg _409637_409637 ; 
   reg __409637_409637;
   reg _409638_409638 ; 
   reg __409638_409638;
   reg _409639_409639 ; 
   reg __409639_409639;
   reg _409640_409640 ; 
   reg __409640_409640;
   reg _409641_409641 ; 
   reg __409641_409641;
   reg _409642_409642 ; 
   reg __409642_409642;
   reg _409643_409643 ; 
   reg __409643_409643;
   reg _409644_409644 ; 
   reg __409644_409644;
   reg _409645_409645 ; 
   reg __409645_409645;
   reg _409646_409646 ; 
   reg __409646_409646;
   reg _409647_409647 ; 
   reg __409647_409647;
   reg _409648_409648 ; 
   reg __409648_409648;
   reg _409649_409649 ; 
   reg __409649_409649;
   reg _409650_409650 ; 
   reg __409650_409650;
   reg _409651_409651 ; 
   reg __409651_409651;
   reg _409652_409652 ; 
   reg __409652_409652;
   reg _409653_409653 ; 
   reg __409653_409653;
   reg _409654_409654 ; 
   reg __409654_409654;
   reg _409655_409655 ; 
   reg __409655_409655;
   reg _409656_409656 ; 
   reg __409656_409656;
   reg _409657_409657 ; 
   reg __409657_409657;
   reg _409658_409658 ; 
   reg __409658_409658;
   reg _409659_409659 ; 
   reg __409659_409659;
   reg _409660_409660 ; 
   reg __409660_409660;
   reg _409661_409661 ; 
   reg __409661_409661;
   reg _409662_409662 ; 
   reg __409662_409662;
   reg _409663_409663 ; 
   reg __409663_409663;
   reg _409664_409664 ; 
   reg __409664_409664;
   reg _409665_409665 ; 
   reg __409665_409665;
   reg _409666_409666 ; 
   reg __409666_409666;
   reg _409667_409667 ; 
   reg __409667_409667;
   reg _409668_409668 ; 
   reg __409668_409668;
   reg _409669_409669 ; 
   reg __409669_409669;
   reg _409670_409670 ; 
   reg __409670_409670;
   reg _409671_409671 ; 
   reg __409671_409671;
   reg _409672_409672 ; 
   reg __409672_409672;
   reg _409673_409673 ; 
   reg __409673_409673;
   reg _409674_409674 ; 
   reg __409674_409674;
   reg _409675_409675 ; 
   reg __409675_409675;
   reg _409676_409676 ; 
   reg __409676_409676;
   reg _409677_409677 ; 
   reg __409677_409677;
   reg _409678_409678 ; 
   reg __409678_409678;
   reg _409679_409679 ; 
   reg __409679_409679;
   reg _409680_409680 ; 
   reg __409680_409680;
   reg _409681_409681 ; 
   reg __409681_409681;
   reg _409682_409682 ; 
   reg __409682_409682;
   reg _409683_409683 ; 
   reg __409683_409683;
   reg _409684_409684 ; 
   reg __409684_409684;
   reg _409685_409685 ; 
   reg __409685_409685;
   reg _409686_409686 ; 
   reg __409686_409686;
   reg _409687_409687 ; 
   reg __409687_409687;
   reg _409688_409688 ; 
   reg __409688_409688;
   reg _409689_409689 ; 
   reg __409689_409689;
   reg _409690_409690 ; 
   reg __409690_409690;
   reg _409691_409691 ; 
   reg __409691_409691;
   reg _409692_409692 ; 
   reg __409692_409692;
   reg _409693_409693 ; 
   reg __409693_409693;
   reg _409694_409694 ; 
   reg __409694_409694;
   reg _409695_409695 ; 
   reg __409695_409695;
   reg _409696_409696 ; 
   reg __409696_409696;
   reg _409697_409697 ; 
   reg __409697_409697;
   reg _409698_409698 ; 
   reg __409698_409698;
   reg _409699_409699 ; 
   reg __409699_409699;
   reg _409700_409700 ; 
   reg __409700_409700;
   reg _409701_409701 ; 
   reg __409701_409701;
   reg _409702_409702 ; 
   reg __409702_409702;
   reg _409703_409703 ; 
   reg __409703_409703;
   reg _409704_409704 ; 
   reg __409704_409704;
   reg _409705_409705 ; 
   reg __409705_409705;
   reg _409706_409706 ; 
   reg __409706_409706;
   reg _409707_409707 ; 
   reg __409707_409707;
   reg _409708_409708 ; 
   reg __409708_409708;
   reg _409709_409709 ; 
   reg __409709_409709;
   reg _409710_409710 ; 
   reg __409710_409710;
   reg _409711_409711 ; 
   reg __409711_409711;
   reg _409712_409712 ; 
   reg __409712_409712;
   reg _409713_409713 ; 
   reg __409713_409713;
   reg _409714_409714 ; 
   reg __409714_409714;
   reg _409715_409715 ; 
   reg __409715_409715;
   reg _409716_409716 ; 
   reg __409716_409716;
   reg _409717_409717 ; 
   reg __409717_409717;
   reg _409718_409718 ; 
   reg __409718_409718;
   reg _409719_409719 ; 
   reg __409719_409719;
   reg _409720_409720 ; 
   reg __409720_409720;
   reg _409721_409721 ; 
   reg __409721_409721;
   reg _409722_409722 ; 
   reg __409722_409722;
   reg _409723_409723 ; 
   reg __409723_409723;
   reg _409724_409724 ; 
   reg __409724_409724;
   reg _409725_409725 ; 
   reg __409725_409725;
   reg _409726_409726 ; 
   reg __409726_409726;
   reg _409727_409727 ; 
   reg __409727_409727;
   reg _409728_409728 ; 
   reg __409728_409728;
   reg _409729_409729 ; 
   reg __409729_409729;
   reg _409730_409730 ; 
   reg __409730_409730;
   reg _409731_409731 ; 
   reg __409731_409731;
   reg _409732_409732 ; 
   reg __409732_409732;
   reg _409733_409733 ; 
   reg __409733_409733;
   reg _409734_409734 ; 
   reg __409734_409734;
   reg _409735_409735 ; 
   reg __409735_409735;
   reg _409736_409736 ; 
   reg __409736_409736;
   reg _409737_409737 ; 
   reg __409737_409737;
   reg _409738_409738 ; 
   reg __409738_409738;
   reg _409739_409739 ; 
   reg __409739_409739;
   reg _409740_409740 ; 
   reg __409740_409740;
   reg _409741_409741 ; 
   reg __409741_409741;
   reg _409742_409742 ; 
   reg __409742_409742;
   reg _409743_409743 ; 
   reg __409743_409743;
   reg _409744_409744 ; 
   reg __409744_409744;
   reg _409745_409745 ; 
   reg __409745_409745;
   reg _409746_409746 ; 
   reg __409746_409746;
   reg _409747_409747 ; 
   reg __409747_409747;
   reg _409748_409748 ; 
   reg __409748_409748;
   reg _409749_409749 ; 
   reg __409749_409749;
   reg _409750_409750 ; 
   reg __409750_409750;
   reg _409751_409751 ; 
   reg __409751_409751;
   reg _409752_409752 ; 
   reg __409752_409752;
   reg _409753_409753 ; 
   reg __409753_409753;
   reg _409754_409754 ; 
   reg __409754_409754;
   reg _409755_409755 ; 
   reg __409755_409755;
   reg _409756_409756 ; 
   reg __409756_409756;
   reg _409757_409757 ; 
   reg __409757_409757;
   reg _409758_409758 ; 
   reg __409758_409758;
   reg _409759_409759 ; 
   reg __409759_409759;
   reg _409760_409760 ; 
   reg __409760_409760;
   reg _409761_409761 ; 
   reg __409761_409761;
   reg _409762_409762 ; 
   reg __409762_409762;
   reg _409763_409763 ; 
   reg __409763_409763;
   reg _409764_409764 ; 
   reg __409764_409764;
   reg _409765_409765 ; 
   reg __409765_409765;
   reg _409766_409766 ; 
   reg __409766_409766;
   reg _409767_409767 ; 
   reg __409767_409767;
   reg _409768_409768 ; 
   reg __409768_409768;
   reg _409769_409769 ; 
   reg __409769_409769;
   reg _409770_409770 ; 
   reg __409770_409770;
   reg _409771_409771 ; 
   reg __409771_409771;
   reg _409772_409772 ; 
   reg __409772_409772;
   reg _409773_409773 ; 
   reg __409773_409773;
   reg _409774_409774 ; 
   reg __409774_409774;
   reg _409775_409775 ; 
   reg __409775_409775;
   reg _409776_409776 ; 
   reg __409776_409776;
   reg _409777_409777 ; 
   reg __409777_409777;
   reg _409778_409778 ; 
   reg __409778_409778;
   reg _409779_409779 ; 
   reg __409779_409779;
   reg _409780_409780 ; 
   reg __409780_409780;
   reg _409781_409781 ; 
   reg __409781_409781;
   reg _409782_409782 ; 
   reg __409782_409782;
   reg _409783_409783 ; 
   reg __409783_409783;
   reg _409784_409784 ; 
   reg __409784_409784;
   reg _409785_409785 ; 
   reg __409785_409785;
   reg _409786_409786 ; 
   reg __409786_409786;
   reg _409787_409787 ; 
   reg __409787_409787;
   reg _409788_409788 ; 
   reg __409788_409788;
   reg _409789_409789 ; 
   reg __409789_409789;
   reg _409790_409790 ; 
   reg __409790_409790;
   reg _409791_409791 ; 
   reg __409791_409791;
   reg _409792_409792 ; 
   reg __409792_409792;
   reg _409793_409793 ; 
   reg __409793_409793;
   reg _409794_409794 ; 
   reg __409794_409794;
   reg _409795_409795 ; 
   reg __409795_409795;
   reg _409796_409796 ; 
   reg __409796_409796;
   reg _409797_409797 ; 
   reg __409797_409797;
   reg _409798_409798 ; 
   reg __409798_409798;
   reg _409799_409799 ; 
   reg __409799_409799;
   reg _409800_409800 ; 
   reg __409800_409800;
   reg _409801_409801 ; 
   reg __409801_409801;
   reg _409802_409802 ; 
   reg __409802_409802;
   reg _409803_409803 ; 
   reg __409803_409803;
   reg _409804_409804 ; 
   reg __409804_409804;
   reg _409805_409805 ; 
   reg __409805_409805;
   reg _409806_409806 ; 
   reg __409806_409806;
   reg _409807_409807 ; 
   reg __409807_409807;
   reg _409808_409808 ; 
   reg __409808_409808;
   reg _409809_409809 ; 
   reg __409809_409809;
   reg _409810_409810 ; 
   reg __409810_409810;
   reg _409811_409811 ; 
   reg __409811_409811;
   reg _409812_409812 ; 
   reg __409812_409812;
   reg _409813_409813 ; 
   reg __409813_409813;
   reg _409814_409814 ; 
   reg __409814_409814;
   reg _409815_409815 ; 
   reg __409815_409815;
   reg _409816_409816 ; 
   reg __409816_409816;
   reg _409817_409817 ; 
   reg __409817_409817;
   reg _409818_409818 ; 
   reg __409818_409818;
   reg _409819_409819 ; 
   reg __409819_409819;
   reg _409820_409820 ; 
   reg __409820_409820;
   reg _409821_409821 ; 
   reg __409821_409821;
   reg _409822_409822 ; 
   reg __409822_409822;
   reg _409823_409823 ; 
   reg __409823_409823;
   reg _409824_409824 ; 
   reg __409824_409824;
   reg _409825_409825 ; 
   reg __409825_409825;
   reg _409826_409826 ; 
   reg __409826_409826;
   reg _409827_409827 ; 
   reg __409827_409827;
   reg _409828_409828 ; 
   reg __409828_409828;
   reg _409829_409829 ; 
   reg __409829_409829;
   reg _409830_409830 ; 
   reg __409830_409830;
   reg _409831_409831 ; 
   reg __409831_409831;
   reg _409832_409832 ; 
   reg __409832_409832;
   reg _409833_409833 ; 
   reg __409833_409833;
   reg _409834_409834 ; 
   reg __409834_409834;
   reg _409835_409835 ; 
   reg __409835_409835;
   reg _409836_409836 ; 
   reg __409836_409836;
   reg _409837_409837 ; 
   reg __409837_409837;
   reg _409838_409838 ; 
   reg __409838_409838;
   reg _409839_409839 ; 
   reg __409839_409839;
   reg _409840_409840 ; 
   reg __409840_409840;
   reg _409841_409841 ; 
   reg __409841_409841;
   reg _409842_409842 ; 
   reg __409842_409842;
   reg _409843_409843 ; 
   reg __409843_409843;
   reg _409844_409844 ; 
   reg __409844_409844;
   reg _409845_409845 ; 
   reg __409845_409845;
   reg _409846_409846 ; 
   reg __409846_409846;
   reg _409847_409847 ; 
   reg __409847_409847;
   reg _409848_409848 ; 
   reg __409848_409848;
   reg _409849_409849 ; 
   reg __409849_409849;
   reg _409850_409850 ; 
   reg __409850_409850;
   reg _409851_409851 ; 
   reg __409851_409851;
   reg _409852_409852 ; 
   reg __409852_409852;
   reg _409853_409853 ; 
   reg __409853_409853;
   reg _409854_409854 ; 
   reg __409854_409854;
   reg _409855_409855 ; 
   reg __409855_409855;
   reg _409856_409856 ; 
   reg __409856_409856;
   reg _409857_409857 ; 
   reg __409857_409857;
   reg _409858_409858 ; 
   reg __409858_409858;
   reg _409859_409859 ; 
   reg __409859_409859;
   reg _409860_409860 ; 
   reg __409860_409860;
   reg _409861_409861 ; 
   reg __409861_409861;
   reg _409862_409862 ; 
   reg __409862_409862;
   reg _409863_409863 ; 
   reg __409863_409863;
   reg _409864_409864 ; 
   reg __409864_409864;
   reg _409865_409865 ; 
   reg __409865_409865;
   reg _409866_409866 ; 
   reg __409866_409866;
   reg _409867_409867 ; 
   reg __409867_409867;
   reg _409868_409868 ; 
   reg __409868_409868;
   reg _409869_409869 ; 
   reg __409869_409869;
   reg _409870_409870 ; 
   reg __409870_409870;
   reg _409871_409871 ; 
   reg __409871_409871;
   reg _409872_409872 ; 
   reg __409872_409872;
   reg _409873_409873 ; 
   reg __409873_409873;
   reg _409874_409874 ; 
   reg __409874_409874;
   reg _409875_409875 ; 
   reg __409875_409875;
   reg _409876_409876 ; 
   reg __409876_409876;
   reg _409877_409877 ; 
   reg __409877_409877;
   reg _409878_409878 ; 
   reg __409878_409878;
   reg _409879_409879 ; 
   reg __409879_409879;
   reg _409880_409880 ; 
   reg __409880_409880;
   reg _409881_409881 ; 
   reg __409881_409881;
   reg _409882_409882 ; 
   reg __409882_409882;
   reg _409883_409883 ; 
   reg __409883_409883;
   reg _409884_409884 ; 
   reg __409884_409884;
   reg _409885_409885 ; 
   reg __409885_409885;
   reg _409886_409886 ; 
   reg __409886_409886;
   reg _409887_409887 ; 
   reg __409887_409887;
   reg _409888_409888 ; 
   reg __409888_409888;
   reg _409889_409889 ; 
   reg __409889_409889;
   reg _409890_409890 ; 
   reg __409890_409890;
   reg _409891_409891 ; 
   reg __409891_409891;
   reg _409892_409892 ; 
   reg __409892_409892;
   reg _409893_409893 ; 
   reg __409893_409893;
   reg _409894_409894 ; 
   reg __409894_409894;
   reg _409895_409895 ; 
   reg __409895_409895;
   reg _409896_409896 ; 
   reg __409896_409896;
   reg _409897_409897 ; 
   reg __409897_409897;
   reg _409898_409898 ; 
   reg __409898_409898;
   reg _409899_409899 ; 
   reg __409899_409899;
   reg _409900_409900 ; 
   reg __409900_409900;
   reg _409901_409901 ; 
   reg __409901_409901;
   reg _409902_409902 ; 
   reg __409902_409902;
   reg _409903_409903 ; 
   reg __409903_409903;
   reg _409904_409904 ; 
   reg __409904_409904;
   reg _409905_409905 ; 
   reg __409905_409905;
   reg _409906_409906 ; 
   reg __409906_409906;
   reg _409907_409907 ; 
   reg __409907_409907;
   reg _409908_409908 ; 
   reg __409908_409908;
   reg _409909_409909 ; 
   reg __409909_409909;
   reg _409910_409910 ; 
   reg __409910_409910;
   reg _409911_409911 ; 
   reg __409911_409911;
   reg _409912_409912 ; 
   reg __409912_409912;
   reg _409913_409913 ; 
   reg __409913_409913;
   reg _409914_409914 ; 
   reg __409914_409914;
   reg _409915_409915 ; 
   reg __409915_409915;
   reg _409916_409916 ; 
   reg __409916_409916;
   reg _409917_409917 ; 
   reg __409917_409917;
   reg _409918_409918 ; 
   reg __409918_409918;
   reg _409919_409919 ; 
   reg __409919_409919;
   reg _409920_409920 ; 
   reg __409920_409920;
   reg _409921_409921 ; 
   reg __409921_409921;
   reg _409922_409922 ; 
   reg __409922_409922;
   reg _409923_409923 ; 
   reg __409923_409923;
   reg _409924_409924 ; 
   reg __409924_409924;
   reg _409925_409925 ; 
   reg __409925_409925;
   reg _409926_409926 ; 
   reg __409926_409926;
   reg _409927_409927 ; 
   reg __409927_409927;
   reg _409928_409928 ; 
   reg __409928_409928;
   reg _409929_409929 ; 
   reg __409929_409929;
   reg _409930_409930 ; 
   reg __409930_409930;
   reg _409931_409931 ; 
   reg __409931_409931;
   reg _409932_409932 ; 
   reg __409932_409932;
   reg _409933_409933 ; 
   reg __409933_409933;
   reg _409934_409934 ; 
   reg __409934_409934;
   reg _409935_409935 ; 
   reg __409935_409935;
   reg _409936_409936 ; 
   reg __409936_409936;
   reg _409937_409937 ; 
   reg __409937_409937;
   reg _409938_409938 ; 
   reg __409938_409938;
   reg _409939_409939 ; 
   reg __409939_409939;
   reg _409940_409940 ; 
   reg __409940_409940;
   reg _409941_409941 ; 
   reg __409941_409941;
   reg _409942_409942 ; 
   reg __409942_409942;
   reg _409943_409943 ; 
   reg __409943_409943;
   reg _409944_409944 ; 
   reg __409944_409944;
   reg _409945_409945 ; 
   reg __409945_409945;
   reg _409946_409946 ; 
   reg __409946_409946;
   reg _409947_409947 ; 
   reg __409947_409947;
   reg _409948_409948 ; 
   reg __409948_409948;
   reg _409949_409949 ; 
   reg __409949_409949;
   reg _409950_409950 ; 
   reg __409950_409950;
   reg _409951_409951 ; 
   reg __409951_409951;
   reg _409952_409952 ; 
   reg __409952_409952;
   reg _409953_409953 ; 
   reg __409953_409953;
   reg _409954_409954 ; 
   reg __409954_409954;
   reg _409955_409955 ; 
   reg __409955_409955;
   reg _409956_409956 ; 
   reg __409956_409956;
   reg _409957_409957 ; 
   reg __409957_409957;
   reg _409958_409958 ; 
   reg __409958_409958;
   reg _409959_409959 ; 
   reg __409959_409959;
   reg _409960_409960 ; 
   reg __409960_409960;
   reg _409961_409961 ; 
   reg __409961_409961;
   reg _409962_409962 ; 
   reg __409962_409962;
   reg _409963_409963 ; 
   reg __409963_409963;
   reg _409964_409964 ; 
   reg __409964_409964;
   reg _409965_409965 ; 
   reg __409965_409965;
   reg _409966_409966 ; 
   reg __409966_409966;
   reg _409967_409967 ; 
   reg __409967_409967;
   reg _409968_409968 ; 
   reg __409968_409968;
   reg _409969_409969 ; 
   reg __409969_409969;
   reg _409970_409970 ; 
   reg __409970_409970;
   reg _409971_409971 ; 
   reg __409971_409971;
   reg _409972_409972 ; 
   reg __409972_409972;
   reg _409973_409973 ; 
   reg __409973_409973;
   reg _409974_409974 ; 
   reg __409974_409974;
   reg _409975_409975 ; 
   reg __409975_409975;
   reg _409976_409976 ; 
   reg __409976_409976;
   reg _409977_409977 ; 
   reg __409977_409977;
   reg _409978_409978 ; 
   reg __409978_409978;
   reg _409979_409979 ; 
   reg __409979_409979;
   reg _409980_409980 ; 
   reg __409980_409980;
   reg _409981_409981 ; 
   reg __409981_409981;
   reg _409982_409982 ; 
   reg __409982_409982;
   reg _409983_409983 ; 
   reg __409983_409983;
   reg _409984_409984 ; 
   reg __409984_409984;
   reg _409985_409985 ; 
   reg __409985_409985;
   reg _409986_409986 ; 
   reg __409986_409986;
   reg _409987_409987 ; 
   reg __409987_409987;
   reg _409988_409988 ; 
   reg __409988_409988;
   reg _409989_409989 ; 
   reg __409989_409989;
   reg _409990_409990 ; 
   reg __409990_409990;
   reg _409991_409991 ; 
   reg __409991_409991;
   reg _409992_409992 ; 
   reg __409992_409992;
   reg _409993_409993 ; 
   reg __409993_409993;
   reg _409994_409994 ; 
   reg __409994_409994;
   reg _409995_409995 ; 
   reg __409995_409995;
   reg _409996_409996 ; 
   reg __409996_409996;
   reg _409997_409997 ; 
   reg __409997_409997;
   reg _409998_409998 ; 
   reg __409998_409998;
   reg _409999_409999 ; 
   reg __409999_409999;
   reg _410000_410000 ; 
   reg __410000_410000;
   reg _410001_410001 ; 
   reg __410001_410001;
   reg _410002_410002 ; 
   reg __410002_410002;
   reg _410003_410003 ; 
   reg __410003_410003;
   reg _410004_410004 ; 
   reg __410004_410004;
   reg _410005_410005 ; 
   reg __410005_410005;
   reg _410006_410006 ; 
   reg __410006_410006;
   reg _410007_410007 ; 
   reg __410007_410007;
   reg _410008_410008 ; 
   reg __410008_410008;
   reg _410009_410009 ; 
   reg __410009_410009;
   reg _410010_410010 ; 
   reg __410010_410010;
   reg _410011_410011 ; 
   reg __410011_410011;
   reg _410012_410012 ; 
   reg __410012_410012;
   reg _410013_410013 ; 
   reg __410013_410013;
   reg _410014_410014 ; 
   reg __410014_410014;
   reg _410015_410015 ; 
   reg __410015_410015;
   reg _410016_410016 ; 
   reg __410016_410016;
   reg _410017_410017 ; 
   reg __410017_410017;
   reg _410018_410018 ; 
   reg __410018_410018;
   reg _410019_410019 ; 
   reg __410019_410019;
   reg _410020_410020 ; 
   reg __410020_410020;
   reg _410021_410021 ; 
   reg __410021_410021;
   reg _410022_410022 ; 
   reg __410022_410022;
   reg _410023_410023 ; 
   reg __410023_410023;
   reg _410024_410024 ; 
   reg __410024_410024;
   reg _410025_410025 ; 
   reg __410025_410025;
   reg _410026_410026 ; 
   reg __410026_410026;
   reg _410027_410027 ; 
   reg __410027_410027;
   reg _410028_410028 ; 
   reg __410028_410028;
   reg _410029_410029 ; 
   reg __410029_410029;
   reg _410030_410030 ; 
   reg __410030_410030;
   reg _410031_410031 ; 
   reg __410031_410031;
   reg _410032_410032 ; 
   reg __410032_410032;
   reg _410033_410033 ; 
   reg __410033_410033;
   reg _410034_410034 ; 
   reg __410034_410034;
   reg _410035_410035 ; 
   reg __410035_410035;
   reg _410036_410036 ; 
   reg __410036_410036;
   reg _410037_410037 ; 
   reg __410037_410037;
   reg _410038_410038 ; 
   reg __410038_410038;
   reg _410039_410039 ; 
   reg __410039_410039;
   reg _410040_410040 ; 
   reg __410040_410040;
   reg _410041_410041 ; 
   reg __410041_410041;
   reg _410042_410042 ; 
   reg __410042_410042;
   reg _410043_410043 ; 
   reg __410043_410043;
   reg _410044_410044 ; 
   reg __410044_410044;
   reg _410045_410045 ; 
   reg __410045_410045;
   reg _410046_410046 ; 
   reg __410046_410046;
   reg _410047_410047 ; 
   reg __410047_410047;
   reg _410048_410048 ; 
   reg __410048_410048;
   reg _410049_410049 ; 
   reg __410049_410049;
   reg _410050_410050 ; 
   reg __410050_410050;
   reg _410051_410051 ; 
   reg __410051_410051;
   reg _410052_410052 ; 
   reg __410052_410052;
   reg _410053_410053 ; 
   reg __410053_410053;
   reg _410054_410054 ; 
   reg __410054_410054;
   reg _410055_410055 ; 
   reg __410055_410055;
   reg _410056_410056 ; 
   reg __410056_410056;
   reg _410057_410057 ; 
   reg __410057_410057;
   reg _410058_410058 ; 
   reg __410058_410058;
   reg _410059_410059 ; 
   reg __410059_410059;
   reg _410060_410060 ; 
   reg __410060_410060;
   reg _410061_410061 ; 
   reg __410061_410061;
   reg _410062_410062 ; 
   reg __410062_410062;
   reg _410063_410063 ; 
   reg __410063_410063;
   reg _410064_410064 ; 
   reg __410064_410064;
   reg _410065_410065 ; 
   reg __410065_410065;
   reg _410066_410066 ; 
   reg __410066_410066;
   reg _410067_410067 ; 
   reg __410067_410067;
   reg _410068_410068 ; 
   reg __410068_410068;
   reg _410069_410069 ; 
   reg __410069_410069;
   reg _410070_410070 ; 
   reg __410070_410070;
   reg _410071_410071 ; 
   reg __410071_410071;
   reg _410072_410072 ; 
   reg __410072_410072;
   reg _410073_410073 ; 
   reg __410073_410073;
   reg _410074_410074 ; 
   reg __410074_410074;
   reg _410075_410075 ; 
   reg __410075_410075;
   reg _410076_410076 ; 
   reg __410076_410076;
   reg _410077_410077 ; 
   reg __410077_410077;
   reg _410078_410078 ; 
   reg __410078_410078;
   reg _410079_410079 ; 
   reg __410079_410079;
   reg _410080_410080 ; 
   reg __410080_410080;
   reg _410081_410081 ; 
   reg __410081_410081;
   reg _410082_410082 ; 
   reg __410082_410082;
   reg _410083_410083 ; 
   reg __410083_410083;
   reg _410084_410084 ; 
   reg __410084_410084;
   reg _410085_410085 ; 
   reg __410085_410085;
   reg _410086_410086 ; 
   reg __410086_410086;
   reg _410087_410087 ; 
   reg __410087_410087;
   reg _410088_410088 ; 
   reg __410088_410088;
   reg _410089_410089 ; 
   reg __410089_410089;
   reg _410090_410090 ; 
   reg __410090_410090;
   reg _410091_410091 ; 
   reg __410091_410091;
   reg _410092_410092 ; 
   reg __410092_410092;
   reg _410093_410093 ; 
   reg __410093_410093;
   reg _410094_410094 ; 
   reg __410094_410094;
   reg _410095_410095 ; 
   reg __410095_410095;
   reg _410096_410096 ; 
   reg __410096_410096;
   reg _410097_410097 ; 
   reg __410097_410097;
   reg _410098_410098 ; 
   reg __410098_410098;
   reg _410099_410099 ; 
   reg __410099_410099;
   reg _410100_410100 ; 
   reg __410100_410100;
   reg _410101_410101 ; 
   reg __410101_410101;
   reg _410102_410102 ; 
   reg __410102_410102;
   reg _410103_410103 ; 
   reg __410103_410103;
   reg _410104_410104 ; 
   reg __410104_410104;
   reg _410105_410105 ; 
   reg __410105_410105;
   reg _410106_410106 ; 
   reg __410106_410106;
   reg _410107_410107 ; 
   reg __410107_410107;
   reg _410108_410108 ; 
   reg __410108_410108;
   reg _410109_410109 ; 
   reg __410109_410109;
   reg _410110_410110 ; 
   reg __410110_410110;
   reg _410111_410111 ; 
   reg __410111_410111;
   reg _410112_410112 ; 
   reg __410112_410112;
   reg _410113_410113 ; 
   reg __410113_410113;
   reg _410114_410114 ; 
   reg __410114_410114;
   reg _410115_410115 ; 
   reg __410115_410115;
   reg _410116_410116 ; 
   reg __410116_410116;
   reg _410117_410117 ; 
   reg __410117_410117;
   reg _410118_410118 ; 
   reg __410118_410118;
   reg _410119_410119 ; 
   reg __410119_410119;
   reg _410120_410120 ; 
   reg __410120_410120;
   reg _410121_410121 ; 
   reg __410121_410121;
   reg _410122_410122 ; 
   reg __410122_410122;
   reg _410123_410123 ; 
   reg __410123_410123;
   reg _410124_410124 ; 
   reg __410124_410124;
   reg _410125_410125 ; 
   reg __410125_410125;
   reg _410126_410126 ; 
   reg __410126_410126;
   reg _410127_410127 ; 
   reg __410127_410127;
   reg _410128_410128 ; 
   reg __410128_410128;
   reg _410129_410129 ; 
   reg __410129_410129;
   reg _410130_410130 ; 
   reg __410130_410130;
   reg _410131_410131 ; 
   reg __410131_410131;
   reg _410132_410132 ; 
   reg __410132_410132;
   reg _410133_410133 ; 
   reg __410133_410133;
   reg _410134_410134 ; 
   reg __410134_410134;
   reg _410135_410135 ; 
   reg __410135_410135;
   reg _410136_410136 ; 
   reg __410136_410136;
   reg _410137_410137 ; 
   reg __410137_410137;
   reg _410138_410138 ; 
   reg __410138_410138;
   reg _410139_410139 ; 
   reg __410139_410139;
   reg _410140_410140 ; 
   reg __410140_410140;
   reg _410141_410141 ; 
   reg __410141_410141;
   reg _410142_410142 ; 
   reg __410142_410142;
   reg _410143_410143 ; 
   reg __410143_410143;
   reg _410144_410144 ; 
   reg __410144_410144;
   reg _410145_410145 ; 
   reg __410145_410145;
   reg _410146_410146 ; 
   reg __410146_410146;
   reg _410147_410147 ; 
   reg __410147_410147;
   reg _410148_410148 ; 
   reg __410148_410148;
   reg _410149_410149 ; 
   reg __410149_410149;
   reg _410150_410150 ; 
   reg __410150_410150;
   reg _410151_410151 ; 
   reg __410151_410151;
   reg _410152_410152 ; 
   reg __410152_410152;
   reg _410153_410153 ; 
   reg __410153_410153;
   reg _410154_410154 ; 
   reg __410154_410154;
   reg _410155_410155 ; 
   reg __410155_410155;
   reg _410156_410156 ; 
   reg __410156_410156;
   reg _410157_410157 ; 
   reg __410157_410157;
   reg _410158_410158 ; 
   reg __410158_410158;
   reg _410159_410159 ; 
   reg __410159_410159;
   reg _410160_410160 ; 
   reg __410160_410160;
   reg _410161_410161 ; 
   reg __410161_410161;
   reg _410162_410162 ; 
   reg __410162_410162;
   reg _410163_410163 ; 
   reg __410163_410163;
   reg _410164_410164 ; 
   reg __410164_410164;
   reg _410165_410165 ; 
   reg __410165_410165;
   reg _410166_410166 ; 
   reg __410166_410166;
   reg _410167_410167 ; 
   reg __410167_410167;
   reg _410168_410168 ; 
   reg __410168_410168;
   reg _410169_410169 ; 
   reg __410169_410169;
   reg _410170_410170 ; 
   reg __410170_410170;
   reg _410171_410171 ; 
   reg __410171_410171;
   reg _410172_410172 ; 
   reg __410172_410172;
   reg _410173_410173 ; 
   reg __410173_410173;
   reg _410174_410174 ; 
   reg __410174_410174;
   reg _410175_410175 ; 
   reg __410175_410175;
   reg _410176_410176 ; 
   reg __410176_410176;
   reg _410177_410177 ; 
   reg __410177_410177;
   reg _410178_410178 ; 
   reg __410178_410178;
   reg _410179_410179 ; 
   reg __410179_410179;
   reg _410180_410180 ; 
   reg __410180_410180;
   reg _410181_410181 ; 
   reg __410181_410181;
   reg _410182_410182 ; 
   reg __410182_410182;
   reg _410183_410183 ; 
   reg __410183_410183;
   reg _410184_410184 ; 
   reg __410184_410184;
   reg _410185_410185 ; 
   reg __410185_410185;
   reg _410186_410186 ; 
   reg __410186_410186;
   reg _410187_410187 ; 
   reg __410187_410187;
   reg _410188_410188 ; 
   reg __410188_410188;
   reg _410189_410189 ; 
   reg __410189_410189;
   reg _410190_410190 ; 
   reg __410190_410190;
   reg _410191_410191 ; 
   reg __410191_410191;
   reg _410192_410192 ; 
   reg __410192_410192;
   reg _410193_410193 ; 
   reg __410193_410193;
   reg _410194_410194 ; 
   reg __410194_410194;
   reg _410195_410195 ; 
   reg __410195_410195;
   reg _410196_410196 ; 
   reg __410196_410196;
   reg _410197_410197 ; 
   reg __410197_410197;
   reg _410198_410198 ; 
   reg __410198_410198;
   reg _410199_410199 ; 
   reg __410199_410199;
   reg _410200_410200 ; 
   reg __410200_410200;
   reg _410201_410201 ; 
   reg __410201_410201;
   reg _410202_410202 ; 
   reg __410202_410202;
   reg _410203_410203 ; 
   reg __410203_410203;
   reg _410204_410204 ; 
   reg __410204_410204;
   reg _410205_410205 ; 
   reg __410205_410205;
   reg _410206_410206 ; 
   reg __410206_410206;
   reg _410207_410207 ; 
   reg __410207_410207;
   reg _410208_410208 ; 
   reg __410208_410208;
   reg _410209_410209 ; 
   reg __410209_410209;
   reg _410210_410210 ; 
   reg __410210_410210;
   reg _410211_410211 ; 
   reg __410211_410211;
   reg _410212_410212 ; 
   reg __410212_410212;
   reg _410213_410213 ; 
   reg __410213_410213;
   reg _410214_410214 ; 
   reg __410214_410214;
   reg _410215_410215 ; 
   reg __410215_410215;
   reg _410216_410216 ; 
   reg __410216_410216;
   reg _410217_410217 ; 
   reg __410217_410217;
   reg _410218_410218 ; 
   reg __410218_410218;
   reg _410219_410219 ; 
   reg __410219_410219;
   reg _410220_410220 ; 
   reg __410220_410220;
   reg _410221_410221 ; 
   reg __410221_410221;
   reg _410222_410222 ; 
   reg __410222_410222;
   reg _410223_410223 ; 
   reg __410223_410223;
   reg _410224_410224 ; 
   reg __410224_410224;
   reg _410225_410225 ; 
   reg __410225_410225;
   reg _410226_410226 ; 
   reg __410226_410226;
   reg _410227_410227 ; 
   reg __410227_410227;
   reg _410228_410228 ; 
   reg __410228_410228;
   reg _410229_410229 ; 
   reg __410229_410229;
   reg _410230_410230 ; 
   reg __410230_410230;
   reg _410231_410231 ; 
   reg __410231_410231;
   reg _410232_410232 ; 
   reg __410232_410232;
   reg _410233_410233 ; 
   reg __410233_410233;
   reg _410234_410234 ; 
   reg __410234_410234;
   reg _410235_410235 ; 
   reg __410235_410235;
   reg _410236_410236 ; 
   reg __410236_410236;
   reg _410237_410237 ; 
   reg __410237_410237;
   reg _410238_410238 ; 
   reg __410238_410238;
   reg _410239_410239 ; 
   reg __410239_410239;
   reg _410240_410240 ; 
   reg __410240_410240;
   reg _410241_410241 ; 
   reg __410241_410241;
   reg _410242_410242 ; 
   reg __410242_410242;
   reg _410243_410243 ; 
   reg __410243_410243;
   reg _410244_410244 ; 
   reg __410244_410244;
   reg _410245_410245 ; 
   reg __410245_410245;
   reg _410246_410246 ; 
   reg __410246_410246;
   reg _410247_410247 ; 
   reg __410247_410247;
   reg _410248_410248 ; 
   reg __410248_410248;
   reg _410249_410249 ; 
   reg __410249_410249;
   reg _410250_410250 ; 
   reg __410250_410250;
   reg _410251_410251 ; 
   reg __410251_410251;
   reg _410252_410252 ; 
   reg __410252_410252;
   reg _410253_410253 ; 
   reg __410253_410253;
   reg _410254_410254 ; 
   reg __410254_410254;
   reg _410255_410255 ; 
   reg __410255_410255;
   reg _410256_410256 ; 
   reg __410256_410256;
   reg _410257_410257 ; 
   reg __410257_410257;
   reg _410258_410258 ; 
   reg __410258_410258;
   reg _410259_410259 ; 
   reg __410259_410259;
   reg _410260_410260 ; 
   reg __410260_410260;
   reg _410261_410261 ; 
   reg __410261_410261;
   reg _410262_410262 ; 
   reg __410262_410262;
   reg _410263_410263 ; 
   reg __410263_410263;
   reg _410264_410264 ; 
   reg __410264_410264;
   reg _410265_410265 ; 
   reg __410265_410265;
   reg _410266_410266 ; 
   reg __410266_410266;
   reg _410267_410267 ; 
   reg __410267_410267;
   reg _410268_410268 ; 
   reg __410268_410268;
   reg _410269_410269 ; 
   reg __410269_410269;
   reg _410270_410270 ; 
   reg __410270_410270;
   reg _410271_410271 ; 
   reg __410271_410271;
   reg _410272_410272 ; 
   reg __410272_410272;
   reg _410273_410273 ; 
   reg __410273_410273;
   reg _410274_410274 ; 
   reg __410274_410274;
   reg _410275_410275 ; 
   reg __410275_410275;
   reg _410276_410276 ; 
   reg __410276_410276;
   reg _410277_410277 ; 
   reg __410277_410277;
   reg _410278_410278 ; 
   reg __410278_410278;
   reg _410279_410279 ; 
   reg __410279_410279;
   reg _410280_410280 ; 
   reg __410280_410280;
   reg _410281_410281 ; 
   reg __410281_410281;
   reg _410282_410282 ; 
   reg __410282_410282;
   reg _410283_410283 ; 
   reg __410283_410283;
   reg _410284_410284 ; 
   reg __410284_410284;
   reg _410285_410285 ; 
   reg __410285_410285;
   reg _410286_410286 ; 
   reg __410286_410286;
   reg _410287_410287 ; 
   reg __410287_410287;
   reg _410288_410288 ; 
   reg __410288_410288;
   reg _410289_410289 ; 
   reg __410289_410289;
   reg _410290_410290 ; 
   reg __410290_410290;
   reg _410291_410291 ; 
   reg __410291_410291;
   reg _410292_410292 ; 
   reg __410292_410292;
   reg _410293_410293 ; 
   reg __410293_410293;
   reg _410294_410294 ; 
   reg __410294_410294;
   reg _410295_410295 ; 
   reg __410295_410295;
   reg _410296_410296 ; 
   reg __410296_410296;
   reg _410297_410297 ; 
   reg __410297_410297;
   reg _410298_410298 ; 
   reg __410298_410298;
   reg _410299_410299 ; 
   reg __410299_410299;
   reg _410300_410300 ; 
   reg __410300_410300;
   reg _410301_410301 ; 
   reg __410301_410301;
   reg _410302_410302 ; 
   reg __410302_410302;
   reg _410303_410303 ; 
   reg __410303_410303;
   reg _410304_410304 ; 
   reg __410304_410304;
   reg _410305_410305 ; 
   reg __410305_410305;
   reg _410306_410306 ; 
   reg __410306_410306;
   reg _410307_410307 ; 
   reg __410307_410307;
   reg _410308_410308 ; 
   reg __410308_410308;
   reg _410309_410309 ; 
   reg __410309_410309;
   reg _410310_410310 ; 
   reg __410310_410310;
   reg _410311_410311 ; 
   reg __410311_410311;
   reg _410312_410312 ; 
   reg __410312_410312;
   reg _410313_410313 ; 
   reg __410313_410313;
   reg _410314_410314 ; 
   reg __410314_410314;
   reg _410315_410315 ; 
   reg __410315_410315;
   reg _410316_410316 ; 
   reg __410316_410316;
   reg _410317_410317 ; 
   reg __410317_410317;
   reg _410318_410318 ; 
   reg __410318_410318;
   reg _410319_410319 ; 
   reg __410319_410319;
   reg _410320_410320 ; 
   reg __410320_410320;
   reg _410321_410321 ; 
   reg __410321_410321;
   reg _410322_410322 ; 
   reg __410322_410322;
   reg _410323_410323 ; 
   reg __410323_410323;
   reg _410324_410324 ; 
   reg __410324_410324;
   reg _410325_410325 ; 
   reg __410325_410325;
   reg _410326_410326 ; 
   reg __410326_410326;
   reg _410327_410327 ; 
   reg __410327_410327;
   reg _410328_410328 ; 
   reg __410328_410328;
   reg _410329_410329 ; 
   reg __410329_410329;
   reg _410330_410330 ; 
   reg __410330_410330;
   reg _410331_410331 ; 
   reg __410331_410331;
   reg _410332_410332 ; 
   reg __410332_410332;
   reg _410333_410333 ; 
   reg __410333_410333;
   reg _410334_410334 ; 
   reg __410334_410334;
   reg _410335_410335 ; 
   reg __410335_410335;
   reg _410336_410336 ; 
   reg __410336_410336;
   reg _410337_410337 ; 
   reg __410337_410337;
   reg _410338_410338 ; 
   reg __410338_410338;
   reg _410339_410339 ; 
   reg __410339_410339;
   reg _410340_410340 ; 
   reg __410340_410340;
   reg _410341_410341 ; 
   reg __410341_410341;
   reg _410342_410342 ; 
   reg __410342_410342;
   reg _410343_410343 ; 
   reg __410343_410343;
   reg _410344_410344 ; 
   reg __410344_410344;
   reg _410345_410345 ; 
   reg __410345_410345;
   reg _410346_410346 ; 
   reg __410346_410346;
   reg _410347_410347 ; 
   reg __410347_410347;
   reg _410348_410348 ; 
   reg __410348_410348;
   reg _410349_410349 ; 
   reg __410349_410349;
   reg _410350_410350 ; 
   reg __410350_410350;
   reg _410351_410351 ; 
   reg __410351_410351;
   reg _410352_410352 ; 
   reg __410352_410352;
   reg _410353_410353 ; 
   reg __410353_410353;
   reg _410354_410354 ; 
   reg __410354_410354;
   reg _410355_410355 ; 
   reg __410355_410355;
   reg _410356_410356 ; 
   reg __410356_410356;
   reg _410357_410357 ; 
   reg __410357_410357;
   reg _410358_410358 ; 
   reg __410358_410358;
   reg _410359_410359 ; 
   reg __410359_410359;
   reg _410360_410360 ; 
   reg __410360_410360;
   reg _410361_410361 ; 
   reg __410361_410361;
   reg _410362_410362 ; 
   reg __410362_410362;
   reg _410363_410363 ; 
   reg __410363_410363;
   reg _410364_410364 ; 
   reg __410364_410364;
   reg _410365_410365 ; 
   reg __410365_410365;
   reg _410366_410366 ; 
   reg __410366_410366;
   reg _410367_410367 ; 
   reg __410367_410367;
   reg _410368_410368 ; 
   reg __410368_410368;
   reg _410369_410369 ; 
   reg __410369_410369;
   reg _410370_410370 ; 
   reg __410370_410370;
   reg _410371_410371 ; 
   reg __410371_410371;
   reg _410372_410372 ; 
   reg __410372_410372;
   reg _410373_410373 ; 
   reg __410373_410373;
   reg _410374_410374 ; 
   reg __410374_410374;
   reg _410375_410375 ; 
   reg __410375_410375;
   reg _410376_410376 ; 
   reg __410376_410376;
   reg _410377_410377 ; 
   reg __410377_410377;
   reg _410378_410378 ; 
   reg __410378_410378;
   reg _410379_410379 ; 
   reg __410379_410379;
   reg _410380_410380 ; 
   reg __410380_410380;
   reg _410381_410381 ; 
   reg __410381_410381;
   reg _410382_410382 ; 
   reg __410382_410382;
   reg _410383_410383 ; 
   reg __410383_410383;
   reg _410384_410384 ; 
   reg __410384_410384;
   reg _410385_410385 ; 
   reg __410385_410385;
   reg _410386_410386 ; 
   reg __410386_410386;
   reg _410387_410387 ; 
   reg __410387_410387;
   reg _410388_410388 ; 
   reg __410388_410388;
   reg _410389_410389 ; 
   reg __410389_410389;
   reg _410390_410390 ; 
   reg __410390_410390;
   reg _410391_410391 ; 
   reg __410391_410391;
   reg _410392_410392 ; 
   reg __410392_410392;
   reg _410393_410393 ; 
   reg __410393_410393;
   reg _410394_410394 ; 
   reg __410394_410394;
   reg _410395_410395 ; 
   reg __410395_410395;
   reg _410396_410396 ; 
   reg __410396_410396;
   reg _410397_410397 ; 
   reg __410397_410397;
   reg _410398_410398 ; 
   reg __410398_410398;
   reg _410399_410399 ; 
   reg __410399_410399;
   reg _410400_410400 ; 
   reg __410400_410400;
   reg _410401_410401 ; 
   reg __410401_410401;
   reg _410402_410402 ; 
   reg __410402_410402;
   reg _410403_410403 ; 
   reg __410403_410403;
   reg _410404_410404 ; 
   reg __410404_410404;
   reg _410405_410405 ; 
   reg __410405_410405;
   reg _410406_410406 ; 
   reg __410406_410406;
   reg _410407_410407 ; 
   reg __410407_410407;
   reg _410408_410408 ; 
   reg __410408_410408;
   reg _410409_410409 ; 
   reg __410409_410409;
   reg _410410_410410 ; 
   reg __410410_410410;
   reg _410411_410411 ; 
   reg __410411_410411;
   reg _410412_410412 ; 
   reg __410412_410412;
   reg _410413_410413 ; 
   reg __410413_410413;
   reg _410414_410414 ; 
   reg __410414_410414;
   reg _410415_410415 ; 
   reg __410415_410415;
   reg _410416_410416 ; 
   reg __410416_410416;
   reg _410417_410417 ; 
   reg __410417_410417;
   reg _410418_410418 ; 
   reg __410418_410418;
   reg _410419_410419 ; 
   reg __410419_410419;
   reg _410420_410420 ; 
   reg __410420_410420;
   reg _410421_410421 ; 
   reg __410421_410421;
   reg _410422_410422 ; 
   reg __410422_410422;
   reg _410423_410423 ; 
   reg __410423_410423;
   reg _410424_410424 ; 
   reg __410424_410424;
   reg _410425_410425 ; 
   reg __410425_410425;
   reg _410426_410426 ; 
   reg __410426_410426;
   reg _410427_410427 ; 
   reg __410427_410427;
   reg _410428_410428 ; 
   reg __410428_410428;
   reg _410429_410429 ; 
   reg __410429_410429;
   reg _410430_410430 ; 
   reg __410430_410430;
   reg _410431_410431 ; 
   reg __410431_410431;
   reg _410432_410432 ; 
   reg __410432_410432;
   reg _410433_410433 ; 
   reg __410433_410433;
   reg _410434_410434 ; 
   reg __410434_410434;
   reg _410435_410435 ; 
   reg __410435_410435;
   reg _410436_410436 ; 
   reg __410436_410436;
   reg _410437_410437 ; 
   reg __410437_410437;
   reg _410438_410438 ; 
   reg __410438_410438;
   reg _410439_410439 ; 
   reg __410439_410439;
   reg _410440_410440 ; 
   reg __410440_410440;
   reg _410441_410441 ; 
   reg __410441_410441;
   reg _410442_410442 ; 
   reg __410442_410442;
   reg _410443_410443 ; 
   reg __410443_410443;
   reg _410444_410444 ; 
   reg __410444_410444;
   reg _410445_410445 ; 
   reg __410445_410445;
   reg _410446_410446 ; 
   reg __410446_410446;
   reg _410447_410447 ; 
   reg __410447_410447;
   reg _410448_410448 ; 
   reg __410448_410448;
   reg _410449_410449 ; 
   reg __410449_410449;
   reg _410450_410450 ; 
   reg __410450_410450;
   reg _410451_410451 ; 
   reg __410451_410451;
   reg _410452_410452 ; 
   reg __410452_410452;
   reg _410453_410453 ; 
   reg __410453_410453;
   reg _410454_410454 ; 
   reg __410454_410454;
   reg _410455_410455 ; 
   reg __410455_410455;
   reg _410456_410456 ; 
   reg __410456_410456;
   reg _410457_410457 ; 
   reg __410457_410457;
   reg _410458_410458 ; 
   reg __410458_410458;
   reg _410459_410459 ; 
   reg __410459_410459;
   reg _410460_410460 ; 
   reg __410460_410460;
   reg _410461_410461 ; 
   reg __410461_410461;
   reg _410462_410462 ; 
   reg __410462_410462;
   reg _410463_410463 ; 
   reg __410463_410463;
   reg _410464_410464 ; 
   reg __410464_410464;
   reg _410465_410465 ; 
   reg __410465_410465;
   reg _410466_410466 ; 
   reg __410466_410466;
   reg _410467_410467 ; 
   reg __410467_410467;
   reg _410468_410468 ; 
   reg __410468_410468;
   reg _410469_410469 ; 
   reg __410469_410469;
   reg _410470_410470 ; 
   reg __410470_410470;
   reg _410471_410471 ; 
   reg __410471_410471;
   reg _410472_410472 ; 
   reg __410472_410472;
   reg _410473_410473 ; 
   reg __410473_410473;
   reg _410474_410474 ; 
   reg __410474_410474;
   reg _410475_410475 ; 
   reg __410475_410475;
   reg _410476_410476 ; 
   reg __410476_410476;
   reg _410477_410477 ; 
   reg __410477_410477;
   reg _410478_410478 ; 
   reg __410478_410478;
   reg _410479_410479 ; 
   reg __410479_410479;
   reg _410480_410480 ; 
   reg __410480_410480;
   reg _410481_410481 ; 
   reg __410481_410481;
   reg _410482_410482 ; 
   reg __410482_410482;
   reg _410483_410483 ; 
   reg __410483_410483;
   reg _410484_410484 ; 
   reg __410484_410484;
   reg _410485_410485 ; 
   reg __410485_410485;
   reg _410486_410486 ; 
   reg __410486_410486;
   reg _410487_410487 ; 
   reg __410487_410487;
   reg _410488_410488 ; 
   reg __410488_410488;
   reg _410489_410489 ; 
   reg __410489_410489;
   reg _410490_410490 ; 
   reg __410490_410490;
   reg _410491_410491 ; 
   reg __410491_410491;
   reg _410492_410492 ; 
   reg __410492_410492;
   reg _410493_410493 ; 
   reg __410493_410493;
   reg _410494_410494 ; 
   reg __410494_410494;
   reg _410495_410495 ; 
   reg __410495_410495;
   reg _410496_410496 ; 
   reg __410496_410496;
   reg _410497_410497 ; 
   reg __410497_410497;
   reg _410498_410498 ; 
   reg __410498_410498;
   reg _410499_410499 ; 
   reg __410499_410499;
   reg _410500_410500 ; 
   reg __410500_410500;
   reg _410501_410501 ; 
   reg __410501_410501;
   reg _410502_410502 ; 
   reg __410502_410502;
   reg _410503_410503 ; 
   reg __410503_410503;
   reg _410504_410504 ; 
   reg __410504_410504;
   reg _410505_410505 ; 
   reg __410505_410505;
   reg _410506_410506 ; 
   reg __410506_410506;
   reg _410507_410507 ; 
   reg __410507_410507;
   reg _410508_410508 ; 
   reg __410508_410508;
   reg _410509_410509 ; 
   reg __410509_410509;
   reg _410510_410510 ; 
   reg __410510_410510;
   reg _410511_410511 ; 
   reg __410511_410511;
   reg _410512_410512 ; 
   reg __410512_410512;
   reg _410513_410513 ; 
   reg __410513_410513;
   reg _410514_410514 ; 
   reg __410514_410514;
   reg _410515_410515 ; 
   reg __410515_410515;
   reg _410516_410516 ; 
   reg __410516_410516;
   reg _410517_410517 ; 
   reg __410517_410517;
   reg _410518_410518 ; 
   reg __410518_410518;
   reg _410519_410519 ; 
   reg __410519_410519;
   reg _410520_410520 ; 
   reg __410520_410520;
   reg _410521_410521 ; 
   reg __410521_410521;
   reg _410522_410522 ; 
   reg __410522_410522;
   reg _410523_410523 ; 
   reg __410523_410523;
   reg _410524_410524 ; 
   reg __410524_410524;
   reg _410525_410525 ; 
   reg __410525_410525;
   reg _410526_410526 ; 
   reg __410526_410526;
   reg _410527_410527 ; 
   reg __410527_410527;
   reg _410528_410528 ; 
   reg __410528_410528;
   reg _410529_410529 ; 
   reg __410529_410529;
   reg _410530_410530 ; 
   reg __410530_410530;
   reg _410531_410531 ; 
   reg __410531_410531;
   reg _410532_410532 ; 
   reg __410532_410532;
   reg _410533_410533 ; 
   reg __410533_410533;
   reg _410534_410534 ; 
   reg __410534_410534;
   reg _410535_410535 ; 
   reg __410535_410535;
   reg _410536_410536 ; 
   reg __410536_410536;
   reg _410537_410537 ; 
   reg __410537_410537;
   reg _410538_410538 ; 
   reg __410538_410538;
   reg _410539_410539 ; 
   reg __410539_410539;
   reg _410540_410540 ; 
   reg __410540_410540;
   reg _410541_410541 ; 
   reg __410541_410541;
   reg _410542_410542 ; 
   reg __410542_410542;
   reg _410543_410543 ; 
   reg __410543_410543;
   reg _410544_410544 ; 
   reg __410544_410544;
   reg _410545_410545 ; 
   reg __410545_410545;
   reg _410546_410546 ; 
   reg __410546_410546;
   reg _410547_410547 ; 
   reg __410547_410547;
   reg _410548_410548 ; 
   reg __410548_410548;
   reg _410549_410549 ; 
   reg __410549_410549;
   reg _410550_410550 ; 
   reg __410550_410550;
   reg _410551_410551 ; 
   reg __410551_410551;
   reg _410552_410552 ; 
   reg __410552_410552;
   reg _410553_410553 ; 
   reg __410553_410553;
   reg _410554_410554 ; 
   reg __410554_410554;
   reg _410555_410555 ; 
   reg __410555_410555;
   reg _410556_410556 ; 
   reg __410556_410556;
   reg _410557_410557 ; 
   reg __410557_410557;
   reg _410558_410558 ; 
   reg __410558_410558;
   reg _410559_410559 ; 
   reg __410559_410559;
   reg _410560_410560 ; 
   reg __410560_410560;
   reg _410561_410561 ; 
   reg __410561_410561;
   reg _410562_410562 ; 
   reg __410562_410562;
   reg _410563_410563 ; 
   reg __410563_410563;
   reg _410564_410564 ; 
   reg __410564_410564;
   reg _410565_410565 ; 
   reg __410565_410565;
   reg _410566_410566 ; 
   reg __410566_410566;
   reg _410567_410567 ; 
   reg __410567_410567;
   reg _410568_410568 ; 
   reg __410568_410568;
   reg _410569_410569 ; 
   reg __410569_410569;
   reg _410570_410570 ; 
   reg __410570_410570;
   reg _410571_410571 ; 
   reg __410571_410571;
   reg _410572_410572 ; 
   reg __410572_410572;
   reg _410573_410573 ; 
   reg __410573_410573;
   reg _410574_410574 ; 
   reg __410574_410574;
   reg _410575_410575 ; 
   reg __410575_410575;
   reg _410576_410576 ; 
   reg __410576_410576;
   reg _410577_410577 ; 
   reg __410577_410577;
   reg _410578_410578 ; 
   reg __410578_410578;
   reg _410579_410579 ; 
   reg __410579_410579;
   reg _410580_410580 ; 
   reg __410580_410580;
   reg _410581_410581 ; 
   reg __410581_410581;
   reg _410582_410582 ; 
   reg __410582_410582;
   reg _410583_410583 ; 
   reg __410583_410583;
   reg _410584_410584 ; 
   reg __410584_410584;
   reg _410585_410585 ; 
   reg __410585_410585;
   reg _410586_410586 ; 
   reg __410586_410586;
   reg _410587_410587 ; 
   reg __410587_410587;
   reg _410588_410588 ; 
   reg __410588_410588;
   reg _410589_410589 ; 
   reg __410589_410589;
   reg _410590_410590 ; 
   reg __410590_410590;
   reg _410591_410591 ; 
   reg __410591_410591;
   reg _410592_410592 ; 
   reg __410592_410592;
   reg _410593_410593 ; 
   reg __410593_410593;
   reg _410594_410594 ; 
   reg __410594_410594;
   reg _410595_410595 ; 
   reg __410595_410595;
   reg _410596_410596 ; 
   reg __410596_410596;
   reg _410597_410597 ; 
   reg __410597_410597;
   reg _410598_410598 ; 
   reg __410598_410598;
   reg _410599_410599 ; 
   reg __410599_410599;
   reg _410600_410600 ; 
   reg __410600_410600;
   reg _410601_410601 ; 
   reg __410601_410601;
   reg _410602_410602 ; 
   reg __410602_410602;
   reg _410603_410603 ; 
   reg __410603_410603;
   reg _410604_410604 ; 
   reg __410604_410604;
   reg _410605_410605 ; 
   reg __410605_410605;
   reg _410606_410606 ; 
   reg __410606_410606;
   reg _410607_410607 ; 
   reg __410607_410607;
   reg _410608_410608 ; 
   reg __410608_410608;
   reg _410609_410609 ; 
   reg __410609_410609;
   reg _410610_410610 ; 
   reg __410610_410610;
   reg _410611_410611 ; 
   reg __410611_410611;
   reg _410612_410612 ; 
   reg __410612_410612;
   reg _410613_410613 ; 
   reg __410613_410613;
   reg _410614_410614 ; 
   reg __410614_410614;
   reg _410615_410615 ; 
   reg __410615_410615;
   reg _410616_410616 ; 
   reg __410616_410616;
   reg _410617_410617 ; 
   reg __410617_410617;
   reg _410618_410618 ; 
   reg __410618_410618;
   reg _410619_410619 ; 
   reg __410619_410619;
   reg _410620_410620 ; 
   reg __410620_410620;
   reg _410621_410621 ; 
   reg __410621_410621;
   reg _410622_410622 ; 
   reg __410622_410622;
   reg _410623_410623 ; 
   reg __410623_410623;
   reg _410624_410624 ; 
   reg __410624_410624;
   reg _410625_410625 ; 
   reg __410625_410625;
   reg _410626_410626 ; 
   reg __410626_410626;
   reg _410627_410627 ; 
   reg __410627_410627;
   reg _410628_410628 ; 
   reg __410628_410628;
   reg _410629_410629 ; 
   reg __410629_410629;
   reg _410630_410630 ; 
   reg __410630_410630;
   reg _410631_410631 ; 
   reg __410631_410631;
   reg _410632_410632 ; 
   reg __410632_410632;
   reg _410633_410633 ; 
   reg __410633_410633;
   reg _410634_410634 ; 
   reg __410634_410634;
   reg _410635_410635 ; 
   reg __410635_410635;
   reg _410636_410636 ; 
   reg __410636_410636;
   reg _410637_410637 ; 
   reg __410637_410637;
   reg _410638_410638 ; 
   reg __410638_410638;
   reg _410639_410639 ; 
   reg __410639_410639;
   reg _410640_410640 ; 
   reg __410640_410640;
   reg _410641_410641 ; 
   reg __410641_410641;
   reg _410642_410642 ; 
   reg __410642_410642;
   reg _410643_410643 ; 
   reg __410643_410643;
   reg _410644_410644 ; 
   reg __410644_410644;
   reg _410645_410645 ; 
   reg __410645_410645;
   reg _410646_410646 ; 
   reg __410646_410646;
   reg _410647_410647 ; 
   reg __410647_410647;
   reg _410648_410648 ; 
   reg __410648_410648;
   reg _410649_410649 ; 
   reg __410649_410649;
   reg _410650_410650 ; 
   reg __410650_410650;
   reg _410651_410651 ; 
   reg __410651_410651;
   reg _410652_410652 ; 
   reg __410652_410652;
   reg _410653_410653 ; 
   reg __410653_410653;
   reg _410654_410654 ; 
   reg __410654_410654;
   reg _410655_410655 ; 
   reg __410655_410655;
   reg _410656_410656 ; 
   reg __410656_410656;
   reg _410657_410657 ; 
   reg __410657_410657;
   reg _410658_410658 ; 
   reg __410658_410658;
   reg _410659_410659 ; 
   reg __410659_410659;
   reg _410660_410660 ; 
   reg __410660_410660;
   reg _410661_410661 ; 
   reg __410661_410661;
   reg _410662_410662 ; 
   reg __410662_410662;
   reg _410663_410663 ; 
   reg __410663_410663;
   reg _410664_410664 ; 
   reg __410664_410664;
   reg _410665_410665 ; 
   reg __410665_410665;
   reg _410666_410666 ; 
   reg __410666_410666;
   reg _410667_410667 ; 
   reg __410667_410667;
   reg _410668_410668 ; 
   reg __410668_410668;
   reg _410669_410669 ; 
   reg __410669_410669;
   reg _410670_410670 ; 
   reg __410670_410670;
   reg _410671_410671 ; 
   reg __410671_410671;
   reg _410672_410672 ; 
   reg __410672_410672;
   reg _410673_410673 ; 
   reg __410673_410673;
   reg _410674_410674 ; 
   reg __410674_410674;
   reg _410675_410675 ; 
   reg __410675_410675;
   reg _410676_410676 ; 
   reg __410676_410676;
   reg _410677_410677 ; 
   reg __410677_410677;
   reg _410678_410678 ; 
   reg __410678_410678;
   reg _410679_410679 ; 
   reg __410679_410679;
   reg _410680_410680 ; 
   reg __410680_410680;
   reg _410681_410681 ; 
   reg __410681_410681;
   reg _410682_410682 ; 
   reg __410682_410682;
   reg _410683_410683 ; 
   reg __410683_410683;
   reg _410684_410684 ; 
   reg __410684_410684;
   reg _410685_410685 ; 
   reg __410685_410685;
   reg _410686_410686 ; 
   reg __410686_410686;
   reg _410687_410687 ; 
   reg __410687_410687;
   reg _410688_410688 ; 
   reg __410688_410688;
   reg _410689_410689 ; 
   reg __410689_410689;
   reg _410690_410690 ; 
   reg __410690_410690;
   reg _410691_410691 ; 
   reg __410691_410691;
   reg _410692_410692 ; 
   reg __410692_410692;
   reg _410693_410693 ; 
   reg __410693_410693;
   reg _410694_410694 ; 
   reg __410694_410694;
   reg _410695_410695 ; 
   reg __410695_410695;
   reg _410696_410696 ; 
   reg __410696_410696;
   reg _410697_410697 ; 
   reg __410697_410697;
   reg _410698_410698 ; 
   reg __410698_410698;
   reg _410699_410699 ; 
   reg __410699_410699;
   reg _410700_410700 ; 
   reg __410700_410700;
   reg _410701_410701 ; 
   reg __410701_410701;
   reg _410702_410702 ; 
   reg __410702_410702;
   reg _410703_410703 ; 
   reg __410703_410703;
   reg _410704_410704 ; 
   reg __410704_410704;
   reg _410705_410705 ; 
   reg __410705_410705;
   reg _410706_410706 ; 
   reg __410706_410706;
   reg _410707_410707 ; 
   reg __410707_410707;
   reg _410708_410708 ; 
   reg __410708_410708;
   reg _410709_410709 ; 
   reg __410709_410709;
   reg _410710_410710 ; 
   reg __410710_410710;
   reg _410711_410711 ; 
   reg __410711_410711;
   reg _410712_410712 ; 
   reg __410712_410712;
   reg _410713_410713 ; 
   reg __410713_410713;
   reg _410714_410714 ; 
   reg __410714_410714;
   reg _410715_410715 ; 
   reg __410715_410715;
   reg _410716_410716 ; 
   reg __410716_410716;
   reg _410717_410717 ; 
   reg __410717_410717;
   reg _410718_410718 ; 
   reg __410718_410718;
   reg _410719_410719 ; 
   reg __410719_410719;
   reg _410720_410720 ; 
   reg __410720_410720;
   reg _410721_410721 ; 
   reg __410721_410721;
   reg _410722_410722 ; 
   reg __410722_410722;
   reg _410723_410723 ; 
   reg __410723_410723;
   reg _410724_410724 ; 
   reg __410724_410724;
   reg _410725_410725 ; 
   reg __410725_410725;
   reg _410726_410726 ; 
   reg __410726_410726;
   reg _410727_410727 ; 
   reg __410727_410727;
   reg _410728_410728 ; 
   reg __410728_410728;
   reg _410729_410729 ; 
   reg __410729_410729;
   reg _410730_410730 ; 
   reg __410730_410730;
   reg _410731_410731 ; 
   reg __410731_410731;
   reg _410732_410732 ; 
   reg __410732_410732;
   reg _410733_410733 ; 
   reg __410733_410733;
   reg _410734_410734 ; 
   reg __410734_410734;
   reg _410735_410735 ; 
   reg __410735_410735;
   reg _410736_410736 ; 
   reg __410736_410736;
   reg _410737_410737 ; 
   reg __410737_410737;
   reg _410738_410738 ; 
   reg __410738_410738;
   reg _410739_410739 ; 
   reg __410739_410739;
   reg _410740_410740 ; 
   reg __410740_410740;
   reg _410741_410741 ; 
   reg __410741_410741;
   reg _410742_410742 ; 
   reg __410742_410742;
   reg _410743_410743 ; 
   reg __410743_410743;
   reg _410744_410744 ; 
   reg __410744_410744;
   reg _410745_410745 ; 
   reg __410745_410745;
   reg _410746_410746 ; 
   reg __410746_410746;
   reg _410747_410747 ; 
   reg __410747_410747;
   reg _410748_410748 ; 
   reg __410748_410748;
   reg _410749_410749 ; 
   reg __410749_410749;
   reg _410750_410750 ; 
   reg __410750_410750;
   reg _410751_410751 ; 
   reg __410751_410751;
   reg _410752_410752 ; 
   reg __410752_410752;
   reg _410753_410753 ; 
   reg __410753_410753;
   reg _410754_410754 ; 
   reg __410754_410754;
   reg _410755_410755 ; 
   reg __410755_410755;
   reg _410756_410756 ; 
   reg __410756_410756;
   reg _410757_410757 ; 
   reg __410757_410757;
   reg _410758_410758 ; 
   reg __410758_410758;
   reg _410759_410759 ; 
   reg __410759_410759;
   reg _410760_410760 ; 
   reg __410760_410760;
   reg _410761_410761 ; 
   reg __410761_410761;
   reg _410762_410762 ; 
   reg __410762_410762;
   reg _410763_410763 ; 
   reg __410763_410763;
   reg _410764_410764 ; 
   reg __410764_410764;
   reg _410765_410765 ; 
   reg __410765_410765;
   reg _410766_410766 ; 
   reg __410766_410766;
   reg _410767_410767 ; 
   reg __410767_410767;
   reg _410768_410768 ; 
   reg __410768_410768;
   reg _410769_410769 ; 
   reg __410769_410769;
   reg _410770_410770 ; 
   reg __410770_410770;
   reg _410771_410771 ; 
   reg __410771_410771;
   reg _410772_410772 ; 
   reg __410772_410772;
   reg _410773_410773 ; 
   reg __410773_410773;
   reg _410774_410774 ; 
   reg __410774_410774;
   reg _410775_410775 ; 
   reg __410775_410775;
   reg _410776_410776 ; 
   reg __410776_410776;
   reg _410777_410777 ; 
   reg __410777_410777;
   reg _410778_410778 ; 
   reg __410778_410778;
   reg _410779_410779 ; 
   reg __410779_410779;
   reg _410780_410780 ; 
   reg __410780_410780;
   reg _410781_410781 ; 
   reg __410781_410781;
   reg _410782_410782 ; 
   reg __410782_410782;
   reg _410783_410783 ; 
   reg __410783_410783;
   reg _410784_410784 ; 
   reg __410784_410784;
   reg _410785_410785 ; 
   reg __410785_410785;
   reg _410786_410786 ; 
   reg __410786_410786;
   reg _410787_410787 ; 
   reg __410787_410787;
   reg _410788_410788 ; 
   reg __410788_410788;
   reg _410789_410789 ; 
   reg __410789_410789;
   reg _410790_410790 ; 
   reg __410790_410790;
   reg _410791_410791 ; 
   reg __410791_410791;
   reg _410792_410792 ; 
   reg __410792_410792;
   reg _410793_410793 ; 
   reg __410793_410793;
   reg _410794_410794 ; 
   reg __410794_410794;
   reg _410795_410795 ; 
   reg __410795_410795;
   reg _410796_410796 ; 
   reg __410796_410796;
   reg _410797_410797 ; 
   reg __410797_410797;
   reg _410798_410798 ; 
   reg __410798_410798;
   reg _410799_410799 ; 
   reg __410799_410799;
   reg _410800_410800 ; 
   reg __410800_410800;
   reg _410801_410801 ; 
   reg __410801_410801;
   reg _410802_410802 ; 
   reg __410802_410802;
   reg _410803_410803 ; 
   reg __410803_410803;
   reg _410804_410804 ; 
   reg __410804_410804;
   reg _410805_410805 ; 
   reg __410805_410805;
   reg _410806_410806 ; 
   reg __410806_410806;
   reg _410807_410807 ; 
   reg __410807_410807;
   reg _410808_410808 ; 
   reg __410808_410808;
   reg _410809_410809 ; 
   reg __410809_410809;
   reg _410810_410810 ; 
   reg __410810_410810;
   reg _410811_410811 ; 
   reg __410811_410811;
   reg _410812_410812 ; 
   reg __410812_410812;
   reg _410813_410813 ; 
   reg __410813_410813;
   reg _410814_410814 ; 
   reg __410814_410814;
   reg _410815_410815 ; 
   reg __410815_410815;
   reg _410816_410816 ; 
   reg __410816_410816;
   reg _410817_410817 ; 
   reg __410817_410817;
   reg _410818_410818 ; 
   reg __410818_410818;
   reg _410819_410819 ; 
   reg __410819_410819;
   reg _410820_410820 ; 
   reg __410820_410820;
   reg _410821_410821 ; 
   reg __410821_410821;
   reg _410822_410822 ; 
   reg __410822_410822;
   reg _410823_410823 ; 
   reg __410823_410823;
   reg _410824_410824 ; 
   reg __410824_410824;
   reg _410825_410825 ; 
   reg __410825_410825;
   reg _410826_410826 ; 
   reg __410826_410826;
   reg _410827_410827 ; 
   reg __410827_410827;
   reg _410828_410828 ; 
   reg __410828_410828;
   reg _410829_410829 ; 
   reg __410829_410829;
   reg _410830_410830 ; 
   reg __410830_410830;
   reg _410831_410831 ; 
   reg __410831_410831;
   reg _410832_410832 ; 
   reg __410832_410832;
   reg _410833_410833 ; 
   reg __410833_410833;
   reg _410834_410834 ; 
   reg __410834_410834;
   reg _410835_410835 ; 
   reg __410835_410835;
   reg _410836_410836 ; 
   reg __410836_410836;
   reg _410837_410837 ; 
   reg __410837_410837;
   reg _410838_410838 ; 
   reg __410838_410838;
   reg _410839_410839 ; 
   reg __410839_410839;
   reg _410840_410840 ; 
   reg __410840_410840;
   reg _410841_410841 ; 
   reg __410841_410841;
   reg _410842_410842 ; 
   reg __410842_410842;
   reg _410843_410843 ; 
   reg __410843_410843;
   reg _410844_410844 ; 
   reg __410844_410844;
   reg _410845_410845 ; 
   reg __410845_410845;
   reg _410846_410846 ; 
   reg __410846_410846;
   reg _410847_410847 ; 
   reg __410847_410847;
   reg _410848_410848 ; 
   reg __410848_410848;
   reg _410849_410849 ; 
   reg __410849_410849;
   reg _410850_410850 ; 
   reg __410850_410850;
   reg _410851_410851 ; 
   reg __410851_410851;
   reg _410852_410852 ; 
   reg __410852_410852;
   reg _410853_410853 ; 
   reg __410853_410853;
   reg _410854_410854 ; 
   reg __410854_410854;
   reg _410855_410855 ; 
   reg __410855_410855;
   reg _410856_410856 ; 
   reg __410856_410856;
   reg _410857_410857 ; 
   reg __410857_410857;
   reg _410858_410858 ; 
   reg __410858_410858;
   reg _410859_410859 ; 
   reg __410859_410859;
   reg _410860_410860 ; 
   reg __410860_410860;
   reg _410861_410861 ; 
   reg __410861_410861;
   reg _410862_410862 ; 
   reg __410862_410862;
   reg _410863_410863 ; 
   reg __410863_410863;
   reg _410864_410864 ; 
   reg __410864_410864;
   reg _410865_410865 ; 
   reg __410865_410865;
   reg _410866_410866 ; 
   reg __410866_410866;
   reg _410867_410867 ; 
   reg __410867_410867;
   reg _410868_410868 ; 
   reg __410868_410868;
   reg _410869_410869 ; 
   reg __410869_410869;
   reg _410870_410870 ; 
   reg __410870_410870;
   reg _410871_410871 ; 
   reg __410871_410871;
   reg _410872_410872 ; 
   reg __410872_410872;
   reg _410873_410873 ; 
   reg __410873_410873;
   reg _410874_410874 ; 
   reg __410874_410874;
   reg _410875_410875 ; 
   reg __410875_410875;
   reg _410876_410876 ; 
   reg __410876_410876;
   reg _410877_410877 ; 
   reg __410877_410877;
   reg _410878_410878 ; 
   reg __410878_410878;
   reg _410879_410879 ; 
   reg __410879_410879;
   reg _410880_410880 ; 
   reg __410880_410880;
   reg _410881_410881 ; 
   reg __410881_410881;
   reg _410882_410882 ; 
   reg __410882_410882;
   reg _410883_410883 ; 
   reg __410883_410883;
   reg _410884_410884 ; 
   reg __410884_410884;
   reg _410885_410885 ; 
   reg __410885_410885;
   reg _410886_410886 ; 
   reg __410886_410886;
   reg _410887_410887 ; 
   reg __410887_410887;
   reg _410888_410888 ; 
   reg __410888_410888;
   reg _410889_410889 ; 
   reg __410889_410889;
   reg _410890_410890 ; 
   reg __410890_410890;
   reg _410891_410891 ; 
   reg __410891_410891;
   reg _410892_410892 ; 
   reg __410892_410892;
   reg _410893_410893 ; 
   reg __410893_410893;
   reg _410894_410894 ; 
   reg __410894_410894;
   reg _410895_410895 ; 
   reg __410895_410895;
   reg _410896_410896 ; 
   reg __410896_410896;
   reg _410897_410897 ; 
   reg __410897_410897;
   reg _410898_410898 ; 
   reg __410898_410898;
   reg _410899_410899 ; 
   reg __410899_410899;
   reg _410900_410900 ; 
   reg __410900_410900;
   reg _410901_410901 ; 
   reg __410901_410901;
   reg _410902_410902 ; 
   reg __410902_410902;
   reg _410903_410903 ; 
   reg __410903_410903;
   reg _410904_410904 ; 
   reg __410904_410904;
   reg _410905_410905 ; 
   reg __410905_410905;
   reg _410906_410906 ; 
   reg __410906_410906;
   reg _410907_410907 ; 
   reg __410907_410907;
   reg _410908_410908 ; 
   reg __410908_410908;
   reg _410909_410909 ; 
   reg __410909_410909;
   reg _410910_410910 ; 
   reg __410910_410910;
   reg _410911_410911 ; 
   reg __410911_410911;
   reg _410912_410912 ; 
   reg __410912_410912;
   reg _410913_410913 ; 
   reg __410913_410913;
   reg _410914_410914 ; 
   reg __410914_410914;
   reg _410915_410915 ; 
   reg __410915_410915;
   reg _410916_410916 ; 
   reg __410916_410916;
   reg _410917_410917 ; 
   reg __410917_410917;
   reg _410918_410918 ; 
   reg __410918_410918;
   reg _410919_410919 ; 
   reg __410919_410919;
   reg _410920_410920 ; 
   reg __410920_410920;
   reg _410921_410921 ; 
   reg __410921_410921;
   reg _410922_410922 ; 
   reg __410922_410922;
   reg _410923_410923 ; 
   reg __410923_410923;
   reg _410924_410924 ; 
   reg __410924_410924;
   reg _410925_410925 ; 
   reg __410925_410925;
   reg _410926_410926 ; 
   reg __410926_410926;
   reg _410927_410927 ; 
   reg __410927_410927;
   reg _410928_410928 ; 
   reg __410928_410928;
   reg _410929_410929 ; 
   reg __410929_410929;
   reg _410930_410930 ; 
   reg __410930_410930;
   reg _410931_410931 ; 
   reg __410931_410931;
   reg _410932_410932 ; 
   reg __410932_410932;
   reg _410933_410933 ; 
   reg __410933_410933;
   reg _410934_410934 ; 
   reg __410934_410934;
   reg _410935_410935 ; 
   reg __410935_410935;
   reg _410936_410936 ; 
   reg __410936_410936;
   reg _410937_410937 ; 
   reg __410937_410937;
   reg _410938_410938 ; 
   reg __410938_410938;
   reg _410939_410939 ; 
   reg __410939_410939;
   reg _410940_410940 ; 
   reg __410940_410940;
   reg _410941_410941 ; 
   reg __410941_410941;
   reg _410942_410942 ; 
   reg __410942_410942;
   reg _410943_410943 ; 
   reg __410943_410943;
   reg _410944_410944 ; 
   reg __410944_410944;
   reg _410945_410945 ; 
   reg __410945_410945;
   reg _410946_410946 ; 
   reg __410946_410946;
   reg _410947_410947 ; 
   reg __410947_410947;
   reg _410948_410948 ; 
   reg __410948_410948;
   reg _410949_410949 ; 
   reg __410949_410949;
   reg _410950_410950 ; 
   reg __410950_410950;
   reg _410951_410951 ; 
   reg __410951_410951;
   reg _410952_410952 ; 
   reg __410952_410952;
   reg _410953_410953 ; 
   reg __410953_410953;
   reg _410954_410954 ; 
   reg __410954_410954;
   reg _410955_410955 ; 
   reg __410955_410955;
   reg _410956_410956 ; 
   reg __410956_410956;
   reg _410957_410957 ; 
   reg __410957_410957;
   reg _410958_410958 ; 
   reg __410958_410958;
   reg _410959_410959 ; 
   reg __410959_410959;
   reg _410960_410960 ; 
   reg __410960_410960;
   reg _410961_410961 ; 
   reg __410961_410961;
   reg _410962_410962 ; 
   reg __410962_410962;
   reg _410963_410963 ; 
   reg __410963_410963;
   reg _410964_410964 ; 
   reg __410964_410964;
   reg _410965_410965 ; 
   reg __410965_410965;
   reg _410966_410966 ; 
   reg __410966_410966;
   reg _410967_410967 ; 
   reg __410967_410967;
   reg _410968_410968 ; 
   reg __410968_410968;
   reg _410969_410969 ; 
   reg __410969_410969;
   reg _410970_410970 ; 
   reg __410970_410970;
   reg _410971_410971 ; 
   reg __410971_410971;
   reg _410972_410972 ; 
   reg __410972_410972;
   reg _410973_410973 ; 
   reg __410973_410973;
   reg _410974_410974 ; 
   reg __410974_410974;
   reg _410975_410975 ; 
   reg __410975_410975;
   reg _410976_410976 ; 
   reg __410976_410976;
   reg _410977_410977 ; 
   reg __410977_410977;
   reg _410978_410978 ; 
   reg __410978_410978;
   reg _410979_410979 ; 
   reg __410979_410979;
   reg _410980_410980 ; 
   reg __410980_410980;
   reg _410981_410981 ; 
   reg __410981_410981;
   reg _410982_410982 ; 
   reg __410982_410982;
   reg _410983_410983 ; 
   reg __410983_410983;
   reg _410984_410984 ; 
   reg __410984_410984;
   reg _410985_410985 ; 
   reg __410985_410985;
   reg _410986_410986 ; 
   reg __410986_410986;
   reg _410987_410987 ; 
   reg __410987_410987;
   reg _410988_410988 ; 
   reg __410988_410988;
   reg _410989_410989 ; 
   reg __410989_410989;
   reg _410990_410990 ; 
   reg __410990_410990;
   reg _410991_410991 ; 
   reg __410991_410991;
   reg _410992_410992 ; 
   reg __410992_410992;
   reg _410993_410993 ; 
   reg __410993_410993;
   reg _410994_410994 ; 
   reg __410994_410994;
   reg _410995_410995 ; 
   reg __410995_410995;
   reg _410996_410996 ; 
   reg __410996_410996;
   reg _410997_410997 ; 
   reg __410997_410997;
   reg _410998_410998 ; 
   reg __410998_410998;
   reg _410999_410999 ; 
   reg __410999_410999;
   reg _411000_411000 ; 
   reg __411000_411000;
   reg _411001_411001 ; 
   reg __411001_411001;
   reg _411002_411002 ; 
   reg __411002_411002;
   reg _411003_411003 ; 
   reg __411003_411003;
   reg _411004_411004 ; 
   reg __411004_411004;
   reg _411005_411005 ; 
   reg __411005_411005;
   reg _411006_411006 ; 
   reg __411006_411006;
   reg _411007_411007 ; 
   reg __411007_411007;
   reg _411008_411008 ; 
   reg __411008_411008;
   reg _411009_411009 ; 
   reg __411009_411009;
   reg _411010_411010 ; 
   reg __411010_411010;
   reg _411011_411011 ; 
   reg __411011_411011;
   reg _411012_411012 ; 
   reg __411012_411012;
   reg _411013_411013 ; 
   reg __411013_411013;
   reg _411014_411014 ; 
   reg __411014_411014;
   reg _411015_411015 ; 
   reg __411015_411015;
   reg _411016_411016 ; 
   reg __411016_411016;
   reg _411017_411017 ; 
   reg __411017_411017;
   reg _411018_411018 ; 
   reg __411018_411018;
   reg _411019_411019 ; 
   reg __411019_411019;
   reg _411020_411020 ; 
   reg __411020_411020;
   reg _411021_411021 ; 
   reg __411021_411021;
   reg _411022_411022 ; 
   reg __411022_411022;
   reg _411023_411023 ; 
   reg __411023_411023;
   reg _411024_411024 ; 
   reg __411024_411024;
   reg _411025_411025 ; 
   reg __411025_411025;
   reg _411026_411026 ; 
   reg __411026_411026;
   reg _411027_411027 ; 
   reg __411027_411027;
   reg _411028_411028 ; 
   reg __411028_411028;
   reg _411029_411029 ; 
   reg __411029_411029;
   reg _411030_411030 ; 
   reg __411030_411030;
   reg _411031_411031 ; 
   reg __411031_411031;
   reg _411032_411032 ; 
   reg __411032_411032;
   reg _411033_411033 ; 
   reg __411033_411033;
   reg _411034_411034 ; 
   reg __411034_411034;
   reg _411035_411035 ; 
   reg __411035_411035;
   reg _411036_411036 ; 
   reg __411036_411036;
   reg _411037_411037 ; 
   reg __411037_411037;
   reg _411038_411038 ; 
   reg __411038_411038;
   reg _411039_411039 ; 
   reg __411039_411039;
   reg _411040_411040 ; 
   reg __411040_411040;
   reg _411041_411041 ; 
   reg __411041_411041;
   reg _411042_411042 ; 
   reg __411042_411042;
   reg _411043_411043 ; 
   reg __411043_411043;
   reg _411044_411044 ; 
   reg __411044_411044;
   reg _411045_411045 ; 
   reg __411045_411045;
   reg _411046_411046 ; 
   reg __411046_411046;
   reg _411047_411047 ; 
   reg __411047_411047;
   reg _411048_411048 ; 
   reg __411048_411048;
   reg _411049_411049 ; 
   reg __411049_411049;
   reg _411050_411050 ; 
   reg __411050_411050;
   reg _411051_411051 ; 
   reg __411051_411051;
   reg _411052_411052 ; 
   reg __411052_411052;
   reg _411053_411053 ; 
   reg __411053_411053;
   reg _411054_411054 ; 
   reg __411054_411054;
   reg _411055_411055 ; 
   reg __411055_411055;
   reg _411056_411056 ; 
   reg __411056_411056;
   reg _411057_411057 ; 
   reg __411057_411057;
   reg _411058_411058 ; 
   reg __411058_411058;
   reg _411059_411059 ; 
   reg __411059_411059;
   reg _411060_411060 ; 
   reg __411060_411060;
   reg _411061_411061 ; 
   reg __411061_411061;
   reg _411062_411062 ; 
   reg __411062_411062;
   reg _411063_411063 ; 
   reg __411063_411063;
   reg _411064_411064 ; 
   reg __411064_411064;
   reg _411065_411065 ; 
   reg __411065_411065;
   reg _411066_411066 ; 
   reg __411066_411066;
   reg _411067_411067 ; 
   reg __411067_411067;
   reg _411068_411068 ; 
   reg __411068_411068;
   reg _411069_411069 ; 
   reg __411069_411069;
   reg _411070_411070 ; 
   reg __411070_411070;
   reg _411071_411071 ; 
   reg __411071_411071;
   reg _411072_411072 ; 
   reg __411072_411072;
   reg _411073_411073 ; 
   reg __411073_411073;
   reg _411074_411074 ; 
   reg __411074_411074;
   reg _411075_411075 ; 
   reg __411075_411075;
   reg _411076_411076 ; 
   reg __411076_411076;
   reg _411077_411077 ; 
   reg __411077_411077;
   reg _411078_411078 ; 
   reg __411078_411078;
   reg _411079_411079 ; 
   reg __411079_411079;
   reg _411080_411080 ; 
   reg __411080_411080;
   reg _411081_411081 ; 
   reg __411081_411081;
   reg _411082_411082 ; 
   reg __411082_411082;
   reg _411083_411083 ; 
   reg __411083_411083;
   reg _411084_411084 ; 
   reg __411084_411084;
   reg _411085_411085 ; 
   reg __411085_411085;
   reg _411086_411086 ; 
   reg __411086_411086;
   reg _411087_411087 ; 
   reg __411087_411087;
   reg _411088_411088 ; 
   reg __411088_411088;
   reg _411089_411089 ; 
   reg __411089_411089;
   reg _411090_411090 ; 
   reg __411090_411090;
   reg _411091_411091 ; 
   reg __411091_411091;
   reg _411092_411092 ; 
   reg __411092_411092;
   reg _411093_411093 ; 
   reg __411093_411093;
   reg _411094_411094 ; 
   reg __411094_411094;
   reg _411095_411095 ; 
   reg __411095_411095;
   reg _411096_411096 ; 
   reg __411096_411096;
   reg _411097_411097 ; 
   reg __411097_411097;
   reg _411098_411098 ; 
   reg __411098_411098;
   reg _411099_411099 ; 
   reg __411099_411099;
   reg _411100_411100 ; 
   reg __411100_411100;
   reg _411101_411101 ; 
   reg __411101_411101;
   reg _411102_411102 ; 
   reg __411102_411102;
   reg _411103_411103 ; 
   reg __411103_411103;
   reg _411104_411104 ; 
   reg __411104_411104;
   reg _411105_411105 ; 
   reg __411105_411105;
   reg _411106_411106 ; 
   reg __411106_411106;
   reg _411107_411107 ; 
   reg __411107_411107;
   reg _411108_411108 ; 
   reg __411108_411108;
   reg _411109_411109 ; 
   reg __411109_411109;
   reg _411110_411110 ; 
   reg __411110_411110;
   reg _411111_411111 ; 
   reg __411111_411111;
   reg _411112_411112 ; 
   reg __411112_411112;
   reg _411113_411113 ; 
   reg __411113_411113;
   reg _411114_411114 ; 
   reg __411114_411114;
   reg _411115_411115 ; 
   reg __411115_411115;
   reg _411116_411116 ; 
   reg __411116_411116;
   reg _411117_411117 ; 
   reg __411117_411117;
   reg _411118_411118 ; 
   reg __411118_411118;
   reg _411119_411119 ; 
   reg __411119_411119;
   reg _411120_411120 ; 
   reg __411120_411120;
   reg _411121_411121 ; 
   reg __411121_411121;
   reg _411122_411122 ; 
   reg __411122_411122;
   reg _411123_411123 ; 
   reg __411123_411123;
   reg _411124_411124 ; 
   reg __411124_411124;
   reg _411125_411125 ; 
   reg __411125_411125;
   reg _411126_411126 ; 
   reg __411126_411126;
   reg _411127_411127 ; 
   reg __411127_411127;
   reg _411128_411128 ; 
   reg __411128_411128;
   reg _411129_411129 ; 
   reg __411129_411129;
   reg _411130_411130 ; 
   reg __411130_411130;
   reg _411131_411131 ; 
   reg __411131_411131;
   reg _411132_411132 ; 
   reg __411132_411132;
   reg _411133_411133 ; 
   reg __411133_411133;
   reg _411134_411134 ; 
   reg __411134_411134;
   reg _411135_411135 ; 
   reg __411135_411135;
   reg _411136_411136 ; 
   reg __411136_411136;
   reg _411137_411137 ; 
   reg __411137_411137;
   reg _411138_411138 ; 
   reg __411138_411138;
   reg _411139_411139 ; 
   reg __411139_411139;
   reg _411140_411140 ; 
   reg __411140_411140;
   reg _411141_411141 ; 
   reg __411141_411141;
   reg _411142_411142 ; 
   reg __411142_411142;
   reg _411143_411143 ; 
   reg __411143_411143;
   reg _411144_411144 ; 
   reg __411144_411144;
   reg _411145_411145 ; 
   reg __411145_411145;
   reg _411146_411146 ; 
   reg __411146_411146;
   reg _411147_411147 ; 
   reg __411147_411147;
   reg _411148_411148 ; 
   reg __411148_411148;
   reg _411149_411149 ; 
   reg __411149_411149;
   reg _411150_411150 ; 
   reg __411150_411150;
   reg _411151_411151 ; 
   reg __411151_411151;
   reg _411152_411152 ; 
   reg __411152_411152;
   reg _411153_411153 ; 
   reg __411153_411153;
   reg _411154_411154 ; 
   reg __411154_411154;
   reg _411155_411155 ; 
   reg __411155_411155;
   reg _411156_411156 ; 
   reg __411156_411156;
   reg _411157_411157 ; 
   reg __411157_411157;
   reg _411158_411158 ; 
   reg __411158_411158;
   reg _411159_411159 ; 
   reg __411159_411159;
   reg _411160_411160 ; 
   reg __411160_411160;
   reg _411161_411161 ; 
   reg __411161_411161;
   reg _411162_411162 ; 
   reg __411162_411162;
   reg _411163_411163 ; 
   reg __411163_411163;
   reg _411164_411164 ; 
   reg __411164_411164;
   reg _411165_411165 ; 
   reg __411165_411165;
   reg _411166_411166 ; 
   reg __411166_411166;
   reg _411167_411167 ; 
   reg __411167_411167;
   reg _411168_411168 ; 
   reg __411168_411168;
   reg _411169_411169 ; 
   reg __411169_411169;
   reg _411170_411170 ; 
   reg __411170_411170;
   reg _411171_411171 ; 
   reg __411171_411171;
   reg _411172_411172 ; 
   reg __411172_411172;
   reg _411173_411173 ; 
   reg __411173_411173;
   reg _411174_411174 ; 
   reg __411174_411174;
   reg _411175_411175 ; 
   reg __411175_411175;
   reg _411176_411176 ; 
   reg __411176_411176;
   reg _411177_411177 ; 
   reg __411177_411177;
   reg _411178_411178 ; 
   reg __411178_411178;
   reg _411179_411179 ; 
   reg __411179_411179;
   reg _411180_411180 ; 
   reg __411180_411180;
   reg _411181_411181 ; 
   reg __411181_411181;
   reg _411182_411182 ; 
   reg __411182_411182;
   reg _411183_411183 ; 
   reg __411183_411183;
   reg _411184_411184 ; 
   reg __411184_411184;
   reg _411185_411185 ; 
   reg __411185_411185;
   reg _411186_411186 ; 
   reg __411186_411186;
   reg _411187_411187 ; 
   reg __411187_411187;
   reg _411188_411188 ; 
   reg __411188_411188;
   reg _411189_411189 ; 
   reg __411189_411189;
   reg _411190_411190 ; 
   reg __411190_411190;
   reg _411191_411191 ; 
   reg __411191_411191;
   reg _411192_411192 ; 
   reg __411192_411192;
   reg _411193_411193 ; 
   reg __411193_411193;
   reg _411194_411194 ; 
   reg __411194_411194;
   reg _411195_411195 ; 
   reg __411195_411195;
   reg _411196_411196 ; 
   reg __411196_411196;
   reg _411197_411197 ; 
   reg __411197_411197;
   reg _411198_411198 ; 
   reg __411198_411198;
   reg _411199_411199 ; 
   reg __411199_411199;
   reg _411200_411200 ; 
   reg __411200_411200;
   reg _411201_411201 ; 
   reg __411201_411201;
   reg _411202_411202 ; 
   reg __411202_411202;
   reg _411203_411203 ; 
   reg __411203_411203;
   reg _411204_411204 ; 
   reg __411204_411204;
   reg _411205_411205 ; 
   reg __411205_411205;
   reg _411206_411206 ; 
   reg __411206_411206;
   reg _411207_411207 ; 
   reg __411207_411207;
   reg _411208_411208 ; 
   reg __411208_411208;
   reg _411209_411209 ; 
   reg __411209_411209;
   reg _411210_411210 ; 
   reg __411210_411210;
   reg _411211_411211 ; 
   reg __411211_411211;
   reg _411212_411212 ; 
   reg __411212_411212;
   reg _411213_411213 ; 
   reg __411213_411213;
   reg _411214_411214 ; 
   reg __411214_411214;
   reg _411215_411215 ; 
   reg __411215_411215;
   reg _411216_411216 ; 
   reg __411216_411216;
   reg _411217_411217 ; 
   reg __411217_411217;
   reg _411218_411218 ; 
   reg __411218_411218;
   reg _411219_411219 ; 
   reg __411219_411219;
   reg _411220_411220 ; 
   reg __411220_411220;
   reg _411221_411221 ; 
   reg __411221_411221;
   reg _411222_411222 ; 
   reg __411222_411222;
   reg _411223_411223 ; 
   reg __411223_411223;
   reg _411224_411224 ; 
   reg __411224_411224;
   reg _411225_411225 ; 
   reg __411225_411225;
   reg _411226_411226 ; 
   reg __411226_411226;
   reg _411227_411227 ; 
   reg __411227_411227;
   reg _411228_411228 ; 
   reg __411228_411228;
   reg _411229_411229 ; 
   reg __411229_411229;
   reg _411230_411230 ; 
   reg __411230_411230;
   reg _411231_411231 ; 
   reg __411231_411231;
   reg _411232_411232 ; 
   reg __411232_411232;
   reg _411233_411233 ; 
   reg __411233_411233;
   reg _411234_411234 ; 
   reg __411234_411234;
   reg _411235_411235 ; 
   reg __411235_411235;
   reg _411236_411236 ; 
   reg __411236_411236;
   reg _411237_411237 ; 
   reg __411237_411237;
   reg _411238_411238 ; 
   reg __411238_411238;
   reg _411239_411239 ; 
   reg __411239_411239;
   reg _411240_411240 ; 
   reg __411240_411240;
   reg _411241_411241 ; 
   reg __411241_411241;
   reg _411242_411242 ; 
   reg __411242_411242;
   reg _411243_411243 ; 
   reg __411243_411243;
   reg _411244_411244 ; 
   reg __411244_411244;
   reg _411245_411245 ; 
   reg __411245_411245;
   reg _411246_411246 ; 
   reg __411246_411246;
   reg _411247_411247 ; 
   reg __411247_411247;
   reg _411248_411248 ; 
   reg __411248_411248;
   reg _411249_411249 ; 
   reg __411249_411249;
   reg _411250_411250 ; 
   reg __411250_411250;
   reg _411251_411251 ; 
   reg __411251_411251;
   reg _411252_411252 ; 
   reg __411252_411252;
   reg _411253_411253 ; 
   reg __411253_411253;
   reg _411254_411254 ; 
   reg __411254_411254;
   reg _411255_411255 ; 
   reg __411255_411255;
   reg _411256_411256 ; 
   reg __411256_411256;
   reg _411257_411257 ; 
   reg __411257_411257;
   reg _411258_411258 ; 
   reg __411258_411258;
   reg _411259_411259 ; 
   reg __411259_411259;
   reg _411260_411260 ; 
   reg __411260_411260;
   reg _411261_411261 ; 
   reg __411261_411261;
   reg _411262_411262 ; 
   reg __411262_411262;
   reg _411263_411263 ; 
   reg __411263_411263;
   reg _411264_411264 ; 
   reg __411264_411264;
   reg _411265_411265 ; 
   reg __411265_411265;
   reg _411266_411266 ; 
   reg __411266_411266;
   reg _411267_411267 ; 
   reg __411267_411267;
   reg _411268_411268 ; 
   reg __411268_411268;
   reg _411269_411269 ; 
   reg __411269_411269;
   reg _411270_411270 ; 
   reg __411270_411270;
   reg _411271_411271 ; 
   reg __411271_411271;
   reg _411272_411272 ; 
   reg __411272_411272;
   reg _411273_411273 ; 
   reg __411273_411273;
   reg _411274_411274 ; 
   reg __411274_411274;
   reg _411275_411275 ; 
   reg __411275_411275;
   reg _411276_411276 ; 
   reg __411276_411276;
   reg _411277_411277 ; 
   reg __411277_411277;
   reg _411278_411278 ; 
   reg __411278_411278;
   reg _411279_411279 ; 
   reg __411279_411279;
   reg _411280_411280 ; 
   reg __411280_411280;
   reg _411281_411281 ; 
   reg __411281_411281;
   reg _411282_411282 ; 
   reg __411282_411282;
   reg _411283_411283 ; 
   reg __411283_411283;
   reg _411284_411284 ; 
   reg __411284_411284;
   reg _411285_411285 ; 
   reg __411285_411285;
   reg _411286_411286 ; 
   reg __411286_411286;
   reg _411287_411287 ; 
   reg __411287_411287;
   reg _411288_411288 ; 
   reg __411288_411288;
   reg _411289_411289 ; 
   reg __411289_411289;
   reg _411290_411290 ; 
   reg __411290_411290;
   reg _411291_411291 ; 
   reg __411291_411291;
   reg _411292_411292 ; 
   reg __411292_411292;
   reg _411293_411293 ; 
   reg __411293_411293;
   reg _411294_411294 ; 
   reg __411294_411294;
   reg _411295_411295 ; 
   reg __411295_411295;
   reg _411296_411296 ; 
   reg __411296_411296;
   reg _411297_411297 ; 
   reg __411297_411297;
   reg _411298_411298 ; 
   reg __411298_411298;
   reg _411299_411299 ; 
   reg __411299_411299;
   reg _411300_411300 ; 
   reg __411300_411300;
   reg _411301_411301 ; 
   reg __411301_411301;
   reg _411302_411302 ; 
   reg __411302_411302;
   reg _411303_411303 ; 
   reg __411303_411303;
   reg _411304_411304 ; 
   reg __411304_411304;
   reg _411305_411305 ; 
   reg __411305_411305;
   reg _411306_411306 ; 
   reg __411306_411306;
   reg _411307_411307 ; 
   reg __411307_411307;
   reg _411308_411308 ; 
   reg __411308_411308;
   reg _411309_411309 ; 
   reg __411309_411309;
   reg _411310_411310 ; 
   reg __411310_411310;
   reg _411311_411311 ; 
   reg __411311_411311;
   reg _411312_411312 ; 
   reg __411312_411312;
   reg _411313_411313 ; 
   reg __411313_411313;
   reg _411314_411314 ; 
   reg __411314_411314;
   reg _411315_411315 ; 
   reg __411315_411315;
   reg _411316_411316 ; 
   reg __411316_411316;
   reg _411317_411317 ; 
   reg __411317_411317;
   reg _411318_411318 ; 
   reg __411318_411318;
   reg _411319_411319 ; 
   reg __411319_411319;
   reg _411320_411320 ; 
   reg __411320_411320;
   reg _411321_411321 ; 
   reg __411321_411321;
   reg _411322_411322 ; 
   reg __411322_411322;
   reg _411323_411323 ; 
   reg __411323_411323;
   reg _411324_411324 ; 
   reg __411324_411324;
   reg _411325_411325 ; 
   reg __411325_411325;
   reg _411326_411326 ; 
   reg __411326_411326;
   reg _411327_411327 ; 
   reg __411327_411327;
   reg _411328_411328 ; 
   reg __411328_411328;
   reg _411329_411329 ; 
   reg __411329_411329;
   reg _411330_411330 ; 
   reg __411330_411330;
   reg _411331_411331 ; 
   reg __411331_411331;
   reg _411332_411332 ; 
   reg __411332_411332;
   reg _411333_411333 ; 
   reg __411333_411333;
   reg _411334_411334 ; 
   reg __411334_411334;
   reg _411335_411335 ; 
   reg __411335_411335;
   reg _411336_411336 ; 
   reg __411336_411336;
   reg _411337_411337 ; 
   reg __411337_411337;
   reg _411338_411338 ; 
   reg __411338_411338;
   reg _411339_411339 ; 
   reg __411339_411339;
   reg _411340_411340 ; 
   reg __411340_411340;
   reg _411341_411341 ; 
   reg __411341_411341;
   reg _411342_411342 ; 
   reg __411342_411342;
   reg _411343_411343 ; 
   reg __411343_411343;
   reg _411344_411344 ; 
   reg __411344_411344;
   reg _411345_411345 ; 
   reg __411345_411345;
   reg _411346_411346 ; 
   reg __411346_411346;
   reg _411347_411347 ; 
   reg __411347_411347;
   reg _411348_411348 ; 
   reg __411348_411348;
   reg _411349_411349 ; 
   reg __411349_411349;
   reg _411350_411350 ; 
   reg __411350_411350;
   reg _411351_411351 ; 
   reg __411351_411351;
   reg _411352_411352 ; 
   reg __411352_411352;
   reg _411353_411353 ; 
   reg __411353_411353;
   reg _411354_411354 ; 
   reg __411354_411354;
   reg _411355_411355 ; 
   reg __411355_411355;
   reg _411356_411356 ; 
   reg __411356_411356;
   reg _411357_411357 ; 
   reg __411357_411357;
   reg _411358_411358 ; 
   reg __411358_411358;
   reg _411359_411359 ; 
   reg __411359_411359;
   reg _411360_411360 ; 
   reg __411360_411360;
   reg _411361_411361 ; 
   reg __411361_411361;
   reg _411362_411362 ; 
   reg __411362_411362;
   reg _411363_411363 ; 
   reg __411363_411363;
   reg _411364_411364 ; 
   reg __411364_411364;
   reg _411365_411365 ; 
   reg __411365_411365;
   reg _411366_411366 ; 
   reg __411366_411366;
   reg _411367_411367 ; 
   reg __411367_411367;
   reg _411368_411368 ; 
   reg __411368_411368;
   reg _411369_411369 ; 
   reg __411369_411369;
   reg _411370_411370 ; 
   reg __411370_411370;
   reg _411371_411371 ; 
   reg __411371_411371;
   reg _411372_411372 ; 
   reg __411372_411372;
   reg _411373_411373 ; 
   reg __411373_411373;
   reg _411374_411374 ; 
   reg __411374_411374;
   reg _411375_411375 ; 
   reg __411375_411375;
   reg _411376_411376 ; 
   reg __411376_411376;
   reg _411377_411377 ; 
   reg __411377_411377;
   reg _411378_411378 ; 
   reg __411378_411378;
   reg _411379_411379 ; 
   reg __411379_411379;
   reg _411380_411380 ; 
   reg __411380_411380;
   reg _411381_411381 ; 
   reg __411381_411381;
   reg _411382_411382 ; 
   reg __411382_411382;
   reg _411383_411383 ; 
   reg __411383_411383;
   reg _411384_411384 ; 
   reg __411384_411384;
   reg _411385_411385 ; 
   reg __411385_411385;
   reg _411386_411386 ; 
   reg __411386_411386;
   reg _411387_411387 ; 
   reg __411387_411387;
   reg _411388_411388 ; 
   reg __411388_411388;
   reg _411389_411389 ; 
   reg __411389_411389;
   reg _411390_411390 ; 
   reg __411390_411390;
   reg _411391_411391 ; 
   reg __411391_411391;
   reg _411392_411392 ; 
   reg __411392_411392;
   reg _411393_411393 ; 
   reg __411393_411393;
   reg _411394_411394 ; 
   reg __411394_411394;
   reg _411395_411395 ; 
   reg __411395_411395;
   reg _411396_411396 ; 
   reg __411396_411396;
   reg _411397_411397 ; 
   reg __411397_411397;
   reg _411398_411398 ; 
   reg __411398_411398;
   reg _411399_411399 ; 
   reg __411399_411399;
   reg _411400_411400 ; 
   reg __411400_411400;
   reg _411401_411401 ; 
   reg __411401_411401;
   reg _411402_411402 ; 
   reg __411402_411402;
   reg _411403_411403 ; 
   reg __411403_411403;
   reg _411404_411404 ; 
   reg __411404_411404;
   reg _411405_411405 ; 
   reg __411405_411405;
   reg _411406_411406 ; 
   reg __411406_411406;
   reg _411407_411407 ; 
   reg __411407_411407;
   reg _411408_411408 ; 
   reg __411408_411408;
   reg _411409_411409 ; 
   reg __411409_411409;
   reg _411410_411410 ; 
   reg __411410_411410;
   reg _411411_411411 ; 
   reg __411411_411411;
   reg _411412_411412 ; 
   reg __411412_411412;
   reg _411413_411413 ; 
   reg __411413_411413;
   reg _411414_411414 ; 
   reg __411414_411414;
   reg _411415_411415 ; 
   reg __411415_411415;
   reg _411416_411416 ; 
   reg __411416_411416;
   reg _411417_411417 ; 
   reg __411417_411417;
   reg _411418_411418 ; 
   reg __411418_411418;
   reg _411419_411419 ; 
   reg __411419_411419;
   reg _411420_411420 ; 
   reg __411420_411420;
   reg _411421_411421 ; 
   reg __411421_411421;
   reg _411422_411422 ; 
   reg __411422_411422;
   reg _411423_411423 ; 
   reg __411423_411423;
   reg _411424_411424 ; 
   reg __411424_411424;
   reg _411425_411425 ; 
   reg __411425_411425;
   reg _411426_411426 ; 
   reg __411426_411426;
   reg _411427_411427 ; 
   reg __411427_411427;
   reg _411428_411428 ; 
   reg __411428_411428;
   reg _411429_411429 ; 
   reg __411429_411429;
   reg _411430_411430 ; 
   reg __411430_411430;
   reg _411431_411431 ; 
   reg __411431_411431;
   reg _411432_411432 ; 
   reg __411432_411432;
   reg _411433_411433 ; 
   reg __411433_411433;
   reg _411434_411434 ; 
   reg __411434_411434;
   reg _411435_411435 ; 
   reg __411435_411435;
   reg _411436_411436 ; 
   reg __411436_411436;
   reg _411437_411437 ; 
   reg __411437_411437;
   reg _411438_411438 ; 
   reg __411438_411438;
   reg _411439_411439 ; 
   reg __411439_411439;
   reg _411440_411440 ; 
   reg __411440_411440;
   reg _411441_411441 ; 
   reg __411441_411441;
   reg _411442_411442 ; 
   reg __411442_411442;
   reg _411443_411443 ; 
   reg __411443_411443;
   reg _411444_411444 ; 
   reg __411444_411444;
   reg _411445_411445 ; 
   reg __411445_411445;
   reg _411446_411446 ; 
   reg __411446_411446;
   reg _411447_411447 ; 
   reg __411447_411447;
   reg _411448_411448 ; 
   reg __411448_411448;
   reg _411449_411449 ; 
   reg __411449_411449;
   reg _411450_411450 ; 
   reg __411450_411450;
   reg _411451_411451 ; 
   reg __411451_411451;
   reg _411452_411452 ; 
   reg __411452_411452;
   reg _411453_411453 ; 
   reg __411453_411453;
   reg _411454_411454 ; 
   reg __411454_411454;
   reg _411455_411455 ; 
   reg __411455_411455;
   reg _411456_411456 ; 
   reg __411456_411456;
   reg _411457_411457 ; 
   reg __411457_411457;
   reg _411458_411458 ; 
   reg __411458_411458;
   reg _411459_411459 ; 
   reg __411459_411459;
   reg _411460_411460 ; 
   reg __411460_411460;
   reg _411461_411461 ; 
   reg __411461_411461;
   reg _411462_411462 ; 
   reg __411462_411462;
   reg _411463_411463 ; 
   reg __411463_411463;
   reg _411464_411464 ; 
   reg __411464_411464;
   reg _411465_411465 ; 
   reg __411465_411465;
   reg _411466_411466 ; 
   reg __411466_411466;
   reg _411467_411467 ; 
   reg __411467_411467;
   reg _411468_411468 ; 
   reg __411468_411468;
   reg _411469_411469 ; 
   reg __411469_411469;
   reg _411470_411470 ; 
   reg __411470_411470;
   reg _411471_411471 ; 
   reg __411471_411471;
   reg _411472_411472 ; 
   reg __411472_411472;
   reg _411473_411473 ; 
   reg __411473_411473;
   reg _411474_411474 ; 
   reg __411474_411474;
   reg _411475_411475 ; 
   reg __411475_411475;
   reg _411476_411476 ; 
   reg __411476_411476;
   reg _411477_411477 ; 
   reg __411477_411477;
   reg _411478_411478 ; 
   reg __411478_411478;
   reg _411479_411479 ; 
   reg __411479_411479;
   reg _411480_411480 ; 
   reg __411480_411480;
   reg _411481_411481 ; 
   reg __411481_411481;
   reg _411482_411482 ; 
   reg __411482_411482;
   reg _411483_411483 ; 
   reg __411483_411483;
   reg _411484_411484 ; 
   reg __411484_411484;
   reg _411485_411485 ; 
   reg __411485_411485;
   reg _411486_411486 ; 
   reg __411486_411486;
   reg _411487_411487 ; 
   reg __411487_411487;
   reg _411488_411488 ; 
   reg __411488_411488;
   reg _411489_411489 ; 
   reg __411489_411489;
   reg _411490_411490 ; 
   reg __411490_411490;
   reg _411491_411491 ; 
   reg __411491_411491;
   reg _411492_411492 ; 
   reg __411492_411492;
   reg _411493_411493 ; 
   reg __411493_411493;
   reg _411494_411494 ; 
   reg __411494_411494;
   reg _411495_411495 ; 
   reg __411495_411495;
   reg _411496_411496 ; 
   reg __411496_411496;
   reg _411497_411497 ; 
   reg __411497_411497;
   reg _411498_411498 ; 
   reg __411498_411498;
   reg _411499_411499 ; 
   reg __411499_411499;
   reg _411500_411500 ; 
   reg __411500_411500;
   reg _411501_411501 ; 
   reg __411501_411501;
   reg _411502_411502 ; 
   reg __411502_411502;
   reg _411503_411503 ; 
   reg __411503_411503;
   reg _411504_411504 ; 
   reg __411504_411504;
   reg _411505_411505 ; 
   reg __411505_411505;
   reg _411506_411506 ; 
   reg __411506_411506;
   reg _411507_411507 ; 
   reg __411507_411507;
   reg _411508_411508 ; 
   reg __411508_411508;
   reg _411509_411509 ; 
   reg __411509_411509;
   reg _411510_411510 ; 
   reg __411510_411510;
   reg _411511_411511 ; 
   reg __411511_411511;
   reg _411512_411512 ; 
   reg __411512_411512;
   reg _411513_411513 ; 
   reg __411513_411513;
   reg _411514_411514 ; 
   reg __411514_411514;
   reg _411515_411515 ; 
   reg __411515_411515;
   reg _411516_411516 ; 
   reg __411516_411516;
   reg _411517_411517 ; 
   reg __411517_411517;
   reg _411518_411518 ; 
   reg __411518_411518;
   reg _411519_411519 ; 
   reg __411519_411519;
   reg _411520_411520 ; 
   reg __411520_411520;
   reg _411521_411521 ; 
   reg __411521_411521;
   reg _411522_411522 ; 
   reg __411522_411522;
   reg _411523_411523 ; 
   reg __411523_411523;
   reg _411524_411524 ; 
   reg __411524_411524;
   reg _411525_411525 ; 
   reg __411525_411525;
   reg _411526_411526 ; 
   reg __411526_411526;
   reg _411527_411527 ; 
   reg __411527_411527;
   reg _411528_411528 ; 
   reg __411528_411528;
   reg _411529_411529 ; 
   reg __411529_411529;
   reg _411530_411530 ; 
   reg __411530_411530;
   reg _411531_411531 ; 
   reg __411531_411531;
   reg _411532_411532 ; 
   reg __411532_411532;
   reg _411533_411533 ; 
   reg __411533_411533;
   reg _411534_411534 ; 
   reg __411534_411534;
   reg _411535_411535 ; 
   reg __411535_411535;
   reg _411536_411536 ; 
   reg __411536_411536;
   reg _411537_411537 ; 
   reg __411537_411537;
   reg _411538_411538 ; 
   reg __411538_411538;
   reg _411539_411539 ; 
   reg __411539_411539;
   reg _411540_411540 ; 
   reg __411540_411540;
   reg _411541_411541 ; 
   reg __411541_411541;
   reg _411542_411542 ; 
   reg __411542_411542;
   reg _411543_411543 ; 
   reg __411543_411543;
   reg _411544_411544 ; 
   reg __411544_411544;
   reg _411545_411545 ; 
   reg __411545_411545;
   reg _411546_411546 ; 
   reg __411546_411546;
   reg _411547_411547 ; 
   reg __411547_411547;
   reg _411548_411548 ; 
   reg __411548_411548;
   reg _411549_411549 ; 
   reg __411549_411549;
   reg _411550_411550 ; 
   reg __411550_411550;
   reg _411551_411551 ; 
   reg __411551_411551;
   reg _411552_411552 ; 
   reg __411552_411552;
   reg _411553_411553 ; 
   reg __411553_411553;
   reg _411554_411554 ; 
   reg __411554_411554;
   reg _411555_411555 ; 
   reg __411555_411555;
   reg _411556_411556 ; 
   reg __411556_411556;
   reg _411557_411557 ; 
   reg __411557_411557;
   reg _411558_411558 ; 
   reg __411558_411558;
   reg _411559_411559 ; 
   reg __411559_411559;
   reg _411560_411560 ; 
   reg __411560_411560;
   reg _411561_411561 ; 
   reg __411561_411561;
   reg _411562_411562 ; 
   reg __411562_411562;
   reg _411563_411563 ; 
   reg __411563_411563;
   reg _411564_411564 ; 
   reg __411564_411564;
   reg _411565_411565 ; 
   reg __411565_411565;
   reg _411566_411566 ; 
   reg __411566_411566;
   reg _411567_411567 ; 
   reg __411567_411567;
   reg _411568_411568 ; 
   reg __411568_411568;
   reg _411569_411569 ; 
   reg __411569_411569;
   reg _411570_411570 ; 
   reg __411570_411570;
   reg _411571_411571 ; 
   reg __411571_411571;
   reg _411572_411572 ; 
   reg __411572_411572;
   reg _411573_411573 ; 
   reg __411573_411573;
   reg _411574_411574 ; 
   reg __411574_411574;
   reg _411575_411575 ; 
   reg __411575_411575;
   reg _411576_411576 ; 
   reg __411576_411576;
   reg _411577_411577 ; 
   reg __411577_411577;
   reg _411578_411578 ; 
   reg __411578_411578;
   reg _411579_411579 ; 
   reg __411579_411579;
   reg _411580_411580 ; 
   reg __411580_411580;
   reg _411581_411581 ; 
   reg __411581_411581;
   reg _411582_411582 ; 
   reg __411582_411582;
   reg _411583_411583 ; 
   reg __411583_411583;
   reg _411584_411584 ; 
   reg __411584_411584;
   reg _411585_411585 ; 
   reg __411585_411585;
   reg _411586_411586 ; 
   reg __411586_411586;
   reg _411587_411587 ; 
   reg __411587_411587;
   reg _411588_411588 ; 
   reg __411588_411588;
   reg _411589_411589 ; 
   reg __411589_411589;
   reg _411590_411590 ; 
   reg __411590_411590;
   reg _411591_411591 ; 
   reg __411591_411591;
   reg _411592_411592 ; 
   reg __411592_411592;
   reg _411593_411593 ; 
   reg __411593_411593;
   reg _411594_411594 ; 
   reg __411594_411594;
   reg _411595_411595 ; 
   reg __411595_411595;
   reg _411596_411596 ; 
   reg __411596_411596;
   reg _411597_411597 ; 
   reg __411597_411597;
   reg _411598_411598 ; 
   reg __411598_411598;
   reg _411599_411599 ; 
   reg __411599_411599;
   reg _411600_411600 ; 
   reg __411600_411600;
   reg _411601_411601 ; 
   reg __411601_411601;
   reg _411602_411602 ; 
   reg __411602_411602;
   reg _411603_411603 ; 
   reg __411603_411603;
   reg _411604_411604 ; 
   reg __411604_411604;
   reg _411605_411605 ; 
   reg __411605_411605;
   reg _411606_411606 ; 
   reg __411606_411606;
   reg _411607_411607 ; 
   reg __411607_411607;
   reg _411608_411608 ; 
   reg __411608_411608;
   reg _411609_411609 ; 
   reg __411609_411609;
   reg _411610_411610 ; 
   reg __411610_411610;
   reg _411611_411611 ; 
   reg __411611_411611;
   reg _411612_411612 ; 
   reg __411612_411612;
   reg _411613_411613 ; 
   reg __411613_411613;
   reg _411614_411614 ; 
   reg __411614_411614;
   reg _411615_411615 ; 
   reg __411615_411615;
   reg _411616_411616 ; 
   reg __411616_411616;
   reg _411617_411617 ; 
   reg __411617_411617;
   reg _411618_411618 ; 
   reg __411618_411618;
   reg _411619_411619 ; 
   reg __411619_411619;
   reg _411620_411620 ; 
   reg __411620_411620;
   reg _411621_411621 ; 
   reg __411621_411621;
   reg _411622_411622 ; 
   reg __411622_411622;
   reg _411623_411623 ; 
   reg __411623_411623;
   reg _411624_411624 ; 
   reg __411624_411624;
   reg _411625_411625 ; 
   reg __411625_411625;
   reg _411626_411626 ; 
   reg __411626_411626;
   reg _411627_411627 ; 
   reg __411627_411627;
   reg _411628_411628 ; 
   reg __411628_411628;
   reg _411629_411629 ; 
   reg __411629_411629;
   reg _411630_411630 ; 
   reg __411630_411630;
   reg _411631_411631 ; 
   reg __411631_411631;
   reg _411632_411632 ; 
   reg __411632_411632;
   reg _411633_411633 ; 
   reg __411633_411633;
   reg _411634_411634 ; 
   reg __411634_411634;
   reg _411635_411635 ; 
   reg __411635_411635;
   reg _411636_411636 ; 
   reg __411636_411636;
   reg _411637_411637 ; 
   reg __411637_411637;
   reg _411638_411638 ; 
   reg __411638_411638;
   reg _411639_411639 ; 
   reg __411639_411639;
   reg _411640_411640 ; 
   reg __411640_411640;
   reg _411641_411641 ; 
   reg __411641_411641;
   reg _411642_411642 ; 
   reg __411642_411642;
   reg _411643_411643 ; 
   reg __411643_411643;
   reg _411644_411644 ; 
   reg __411644_411644;
   reg _411645_411645 ; 
   reg __411645_411645;
   reg _411646_411646 ; 
   reg __411646_411646;
   reg _411647_411647 ; 
   reg __411647_411647;
   reg _411648_411648 ; 
   reg __411648_411648;
   reg _411649_411649 ; 
   reg __411649_411649;
   reg _411650_411650 ; 
   reg __411650_411650;
   reg _411651_411651 ; 
   reg __411651_411651;
   reg _411652_411652 ; 
   reg __411652_411652;
   reg _411653_411653 ; 
   reg __411653_411653;
   reg _411654_411654 ; 
   reg __411654_411654;
   reg _411655_411655 ; 
   reg __411655_411655;
   reg _411656_411656 ; 
   reg __411656_411656;
   reg _411657_411657 ; 
   reg __411657_411657;
   reg _411658_411658 ; 
   reg __411658_411658;
   reg _411659_411659 ; 
   reg __411659_411659;
   reg _411660_411660 ; 
   reg __411660_411660;
   reg _411661_411661 ; 
   reg __411661_411661;
   reg _411662_411662 ; 
   reg __411662_411662;
   reg _411663_411663 ; 
   reg __411663_411663;
   reg _411664_411664 ; 
   reg __411664_411664;
   reg _411665_411665 ; 
   reg __411665_411665;
   reg _411666_411666 ; 
   reg __411666_411666;
   reg _411667_411667 ; 
   reg __411667_411667;
   reg _411668_411668 ; 
   reg __411668_411668;
   reg _411669_411669 ; 
   reg __411669_411669;
   reg _411670_411670 ; 
   reg __411670_411670;
   reg _411671_411671 ; 
   reg __411671_411671;
   reg _411672_411672 ; 
   reg __411672_411672;
   reg _411673_411673 ; 
   reg __411673_411673;
   reg _411674_411674 ; 
   reg __411674_411674;
   reg _411675_411675 ; 
   reg __411675_411675;
   reg _411676_411676 ; 
   reg __411676_411676;
   reg _411677_411677 ; 
   reg __411677_411677;
   reg _411678_411678 ; 
   reg __411678_411678;
   reg _411679_411679 ; 
   reg __411679_411679;
   reg _411680_411680 ; 
   reg __411680_411680;
   reg _411681_411681 ; 
   reg __411681_411681;
   reg _411682_411682 ; 
   reg __411682_411682;
   reg _411683_411683 ; 
   reg __411683_411683;
   reg _411684_411684 ; 
   reg __411684_411684;
   reg _411685_411685 ; 
   reg __411685_411685;
   reg _411686_411686 ; 
   reg __411686_411686;
   reg _411687_411687 ; 
   reg __411687_411687;
   reg _411688_411688 ; 
   reg __411688_411688;
   reg _411689_411689 ; 
   reg __411689_411689;
   reg _411690_411690 ; 
   reg __411690_411690;
   reg _411691_411691 ; 
   reg __411691_411691;
   reg _411692_411692 ; 
   reg __411692_411692;
   reg _411693_411693 ; 
   reg __411693_411693;
   reg _411694_411694 ; 
   reg __411694_411694;
   reg _411695_411695 ; 
   reg __411695_411695;
   reg _411696_411696 ; 
   reg __411696_411696;
   reg _411697_411697 ; 
   reg __411697_411697;
   reg _411698_411698 ; 
   reg __411698_411698;
   reg _411699_411699 ; 
   reg __411699_411699;
   reg _411700_411700 ; 
   reg __411700_411700;
   reg _411701_411701 ; 
   reg __411701_411701;
   reg _411702_411702 ; 
   reg __411702_411702;
   reg _411703_411703 ; 
   reg __411703_411703;
   reg _411704_411704 ; 
   reg __411704_411704;
   reg _411705_411705 ; 
   reg __411705_411705;
   reg _411706_411706 ; 
   reg __411706_411706;
   reg _411707_411707 ; 
   reg __411707_411707;
   reg _411708_411708 ; 
   reg __411708_411708;
   reg _411709_411709 ; 
   reg __411709_411709;
   reg _411710_411710 ; 
   reg __411710_411710;
   reg _411711_411711 ; 
   reg __411711_411711;
   reg _411712_411712 ; 
   reg __411712_411712;
   reg _411713_411713 ; 
   reg __411713_411713;
   reg _411714_411714 ; 
   reg __411714_411714;
   reg _411715_411715 ; 
   reg __411715_411715;
   reg _411716_411716 ; 
   reg __411716_411716;
   reg _411717_411717 ; 
   reg __411717_411717;
   reg _411718_411718 ; 
   reg __411718_411718;
   reg _411719_411719 ; 
   reg __411719_411719;
   reg _411720_411720 ; 
   reg __411720_411720;
   reg _411721_411721 ; 
   reg __411721_411721;
   reg _411722_411722 ; 
   reg __411722_411722;
   reg _411723_411723 ; 
   reg __411723_411723;
   reg _411724_411724 ; 
   reg __411724_411724;
   reg _411725_411725 ; 
   reg __411725_411725;
   reg _411726_411726 ; 
   reg __411726_411726;
   reg _411727_411727 ; 
   reg __411727_411727;
   reg _411728_411728 ; 
   reg __411728_411728;
   reg _411729_411729 ; 
   reg __411729_411729;
   reg _411730_411730 ; 
   reg __411730_411730;
   reg _411731_411731 ; 
   reg __411731_411731;
   reg _411732_411732 ; 
   reg __411732_411732;
   reg _411733_411733 ; 
   reg __411733_411733;
   reg _411734_411734 ; 
   reg __411734_411734;
   reg _411735_411735 ; 
   reg __411735_411735;
   reg _411736_411736 ; 
   reg __411736_411736;
   reg _411737_411737 ; 
   reg __411737_411737;
   reg _411738_411738 ; 
   reg __411738_411738;
   reg _411739_411739 ; 
   reg __411739_411739;
   reg _411740_411740 ; 
   reg __411740_411740;
   reg _411741_411741 ; 
   reg __411741_411741;
   reg _411742_411742 ; 
   reg __411742_411742;
   reg _411743_411743 ; 
   reg __411743_411743;
   reg _411744_411744 ; 
   reg __411744_411744;
   reg _411745_411745 ; 
   reg __411745_411745;
   reg _411746_411746 ; 
   reg __411746_411746;
   reg _411747_411747 ; 
   reg __411747_411747;
   reg _411748_411748 ; 
   reg __411748_411748;
   reg _411749_411749 ; 
   reg __411749_411749;
   reg _411750_411750 ; 
   reg __411750_411750;
   reg _411751_411751 ; 
   reg __411751_411751;
   reg _411752_411752 ; 
   reg __411752_411752;
   reg _411753_411753 ; 
   reg __411753_411753;
   reg _411754_411754 ; 
   reg __411754_411754;
   reg _411755_411755 ; 
   reg __411755_411755;
   reg _411756_411756 ; 
   reg __411756_411756;
   reg _411757_411757 ; 
   reg __411757_411757;
   reg _411758_411758 ; 
   reg __411758_411758;
   reg _411759_411759 ; 
   reg __411759_411759;
   reg _411760_411760 ; 
   reg __411760_411760;
   reg _411761_411761 ; 
   reg __411761_411761;
   reg _411762_411762 ; 
   reg __411762_411762;
   reg _411763_411763 ; 
   reg __411763_411763;
   reg _411764_411764 ; 
   reg __411764_411764;
   reg _411765_411765 ; 
   reg __411765_411765;
   reg _411766_411766 ; 
   reg __411766_411766;
   reg _411767_411767 ; 
   reg __411767_411767;
   reg _411768_411768 ; 
   reg __411768_411768;
   reg _411769_411769 ; 
   reg __411769_411769;
   reg _411770_411770 ; 
   reg __411770_411770;
   reg _411771_411771 ; 
   reg __411771_411771;
   reg _411772_411772 ; 
   reg __411772_411772;
   reg _411773_411773 ; 
   reg __411773_411773;
   reg _411774_411774 ; 
   reg __411774_411774;
   reg _411775_411775 ; 
   reg __411775_411775;
   reg _411776_411776 ; 
   reg __411776_411776;
   reg _411777_411777 ; 
   reg __411777_411777;
   reg _411778_411778 ; 
   reg __411778_411778;
   reg _411779_411779 ; 
   reg __411779_411779;
   reg _411780_411780 ; 
   reg __411780_411780;
   reg _411781_411781 ; 
   reg __411781_411781;
   reg _411782_411782 ; 
   reg __411782_411782;
   reg _411783_411783 ; 
   reg __411783_411783;
   reg _411784_411784 ; 
   reg __411784_411784;
   reg _411785_411785 ; 
   reg __411785_411785;
   reg _411786_411786 ; 
   reg __411786_411786;
   reg _411787_411787 ; 
   reg __411787_411787;
   reg _411788_411788 ; 
   reg __411788_411788;
   reg _411789_411789 ; 
   reg __411789_411789;
   reg _411790_411790 ; 
   reg __411790_411790;
   reg _411791_411791 ; 
   reg __411791_411791;
   reg _411792_411792 ; 
   reg __411792_411792;
   reg _411793_411793 ; 
   reg __411793_411793;
   reg _411794_411794 ; 
   reg __411794_411794;
   reg _411795_411795 ; 
   reg __411795_411795;
   reg _411796_411796 ; 
   reg __411796_411796;
   reg _411797_411797 ; 
   reg __411797_411797;
   reg _411798_411798 ; 
   reg __411798_411798;
   reg _411799_411799 ; 
   reg __411799_411799;
   reg _411800_411800 ; 
   reg __411800_411800;
   reg _411801_411801 ; 
   reg __411801_411801;
   reg _411802_411802 ; 
   reg __411802_411802;
   reg _411803_411803 ; 
   reg __411803_411803;
   reg _411804_411804 ; 
   reg __411804_411804;
   reg _411805_411805 ; 
   reg __411805_411805;
   reg _411806_411806 ; 
   reg __411806_411806;
   reg _411807_411807 ; 
   reg __411807_411807;
   reg _411808_411808 ; 
   reg __411808_411808;
   reg _411809_411809 ; 
   reg __411809_411809;
   reg _411810_411810 ; 
   reg __411810_411810;
   reg _411811_411811 ; 
   reg __411811_411811;
   reg _411812_411812 ; 
   reg __411812_411812;
   reg _411813_411813 ; 
   reg __411813_411813;
   reg _411814_411814 ; 
   reg __411814_411814;
   reg _411815_411815 ; 
   reg __411815_411815;
   reg _411816_411816 ; 
   reg __411816_411816;
   reg _411817_411817 ; 
   reg __411817_411817;
   reg _411818_411818 ; 
   reg __411818_411818;
   reg _411819_411819 ; 
   reg __411819_411819;
   reg _411820_411820 ; 
   reg __411820_411820;
   reg _411821_411821 ; 
   reg __411821_411821;
   reg _411822_411822 ; 
   reg __411822_411822;
   reg _411823_411823 ; 
   reg __411823_411823;
   reg _411824_411824 ; 
   reg __411824_411824;
   reg _411825_411825 ; 
   reg __411825_411825;
   reg _411826_411826 ; 
   reg __411826_411826;
   reg _411827_411827 ; 
   reg __411827_411827;
   reg _411828_411828 ; 
   reg __411828_411828;
   reg _411829_411829 ; 
   reg __411829_411829;
   reg _411830_411830 ; 
   reg __411830_411830;
   reg _411831_411831 ; 
   reg __411831_411831;
   reg _411832_411832 ; 
   reg __411832_411832;
   reg _411833_411833 ; 
   reg __411833_411833;
   reg _411834_411834 ; 
   reg __411834_411834;
   reg _411835_411835 ; 
   reg __411835_411835;
   reg _411836_411836 ; 
   reg __411836_411836;
   reg _411837_411837 ; 
   reg __411837_411837;
   reg _411838_411838 ; 
   reg __411838_411838;
   reg _411839_411839 ; 
   reg __411839_411839;
   reg _411840_411840 ; 
   reg __411840_411840;
   reg _411841_411841 ; 
   reg __411841_411841;
   reg _411842_411842 ; 
   reg __411842_411842;
   reg _411843_411843 ; 
   reg __411843_411843;
   reg _411844_411844 ; 
   reg __411844_411844;
   reg _411845_411845 ; 
   reg __411845_411845;
   reg _411846_411846 ; 
   reg __411846_411846;
   reg _411847_411847 ; 
   reg __411847_411847;
   reg _411848_411848 ; 
   reg __411848_411848;
   reg _411849_411849 ; 
   reg __411849_411849;
   reg _411850_411850 ; 
   reg __411850_411850;
   reg _411851_411851 ; 
   reg __411851_411851;
   reg _411852_411852 ; 
   reg __411852_411852;
   reg _411853_411853 ; 
   reg __411853_411853;
   reg _411854_411854 ; 
   reg __411854_411854;
   reg _411855_411855 ; 
   reg __411855_411855;
   reg _411856_411856 ; 
   reg __411856_411856;
   reg _411857_411857 ; 
   reg __411857_411857;
   reg _411858_411858 ; 
   reg __411858_411858;
   reg _411859_411859 ; 
   reg __411859_411859;
   reg _411860_411860 ; 
   reg __411860_411860;
   reg _411861_411861 ; 
   reg __411861_411861;
   reg _411862_411862 ; 
   reg __411862_411862;
   reg _411863_411863 ; 
   reg __411863_411863;
   reg _411864_411864 ; 
   reg __411864_411864;
   reg _411865_411865 ; 
   reg __411865_411865;
   reg _411866_411866 ; 
   reg __411866_411866;
   reg _411867_411867 ; 
   reg __411867_411867;
   reg _411868_411868 ; 
   reg __411868_411868;
   reg _411869_411869 ; 
   reg __411869_411869;
   reg _411870_411870 ; 
   reg __411870_411870;
   reg _411871_411871 ; 
   reg __411871_411871;
   reg _411872_411872 ; 
   reg __411872_411872;
   reg _411873_411873 ; 
   reg __411873_411873;
   reg _411874_411874 ; 
   reg __411874_411874;
   reg _411875_411875 ; 
   reg __411875_411875;
   reg _411876_411876 ; 
   reg __411876_411876;
   reg _411877_411877 ; 
   reg __411877_411877;
   reg _411878_411878 ; 
   reg __411878_411878;
   reg _411879_411879 ; 
   reg __411879_411879;
   reg _411880_411880 ; 
   reg __411880_411880;
   reg _411881_411881 ; 
   reg __411881_411881;
   reg _411882_411882 ; 
   reg __411882_411882;
   reg _411883_411883 ; 
   reg __411883_411883;
   reg _411884_411884 ; 
   reg __411884_411884;
   reg _411885_411885 ; 
   reg __411885_411885;
   reg _411886_411886 ; 
   reg __411886_411886;
   reg _411887_411887 ; 
   reg __411887_411887;
   reg _411888_411888 ; 
   reg __411888_411888;
   reg _411889_411889 ; 
   reg __411889_411889;
   reg _411890_411890 ; 
   reg __411890_411890;
   reg _411891_411891 ; 
   reg __411891_411891;
   reg _411892_411892 ; 
   reg __411892_411892;
   reg _411893_411893 ; 
   reg __411893_411893;
   reg _411894_411894 ; 
   reg __411894_411894;
   reg _411895_411895 ; 
   reg __411895_411895;
   reg _411896_411896 ; 
   reg __411896_411896;
   reg _411897_411897 ; 
   reg __411897_411897;
   reg _411898_411898 ; 
   reg __411898_411898;
   reg _411899_411899 ; 
   reg __411899_411899;
   reg _411900_411900 ; 
   reg __411900_411900;
   reg _411901_411901 ; 
   reg __411901_411901;
   reg _411902_411902 ; 
   reg __411902_411902;
   reg _411903_411903 ; 
   reg __411903_411903;
   reg _411904_411904 ; 
   reg __411904_411904;
   reg _411905_411905 ; 
   reg __411905_411905;
   reg _411906_411906 ; 
   reg __411906_411906;
   reg _411907_411907 ; 
   reg __411907_411907;
   reg _411908_411908 ; 
   reg __411908_411908;
   reg _411909_411909 ; 
   reg __411909_411909;
   reg _411910_411910 ; 
   reg __411910_411910;
   reg _411911_411911 ; 
   reg __411911_411911;
   reg _411912_411912 ; 
   reg __411912_411912;
   reg _411913_411913 ; 
   reg __411913_411913;
   reg _411914_411914 ; 
   reg __411914_411914;
   reg _411915_411915 ; 
   reg __411915_411915;
   reg _411916_411916 ; 
   reg __411916_411916;
   reg _411917_411917 ; 
   reg __411917_411917;
   reg _411918_411918 ; 
   reg __411918_411918;
   reg _411919_411919 ; 
   reg __411919_411919;
   reg _411920_411920 ; 
   reg __411920_411920;
   reg _411921_411921 ; 
   reg __411921_411921;
   reg _411922_411922 ; 
   reg __411922_411922;
   reg _411923_411923 ; 
   reg __411923_411923;
   reg _411924_411924 ; 
   reg __411924_411924;
   reg _411925_411925 ; 
   reg __411925_411925;
   reg _411926_411926 ; 
   reg __411926_411926;
   reg _411927_411927 ; 
   reg __411927_411927;
   reg _411928_411928 ; 
   reg __411928_411928;
   reg _411929_411929 ; 
   reg __411929_411929;
   reg _411930_411930 ; 
   reg __411930_411930;
   reg _411931_411931 ; 
   reg __411931_411931;
   reg _411932_411932 ; 
   reg __411932_411932;
   reg _411933_411933 ; 
   reg __411933_411933;
   reg _411934_411934 ; 
   reg __411934_411934;
   reg _411935_411935 ; 
   reg __411935_411935;
   reg _411936_411936 ; 
   reg __411936_411936;
   reg _411937_411937 ; 
   reg __411937_411937;
   reg _411938_411938 ; 
   reg __411938_411938;
   reg _411939_411939 ; 
   reg __411939_411939;
   reg _411940_411940 ; 
   reg __411940_411940;
   reg _411941_411941 ; 
   reg __411941_411941;
   reg _411942_411942 ; 
   reg __411942_411942;
   reg _411943_411943 ; 
   reg __411943_411943;
   reg _411944_411944 ; 
   reg __411944_411944;
   reg _411945_411945 ; 
   reg __411945_411945;
   reg _411946_411946 ; 
   reg __411946_411946;
   reg _411947_411947 ; 
   reg __411947_411947;
   reg _411948_411948 ; 
   reg __411948_411948;
   reg _411949_411949 ; 
   reg __411949_411949;
   reg _411950_411950 ; 
   reg __411950_411950;
   reg _411951_411951 ; 
   reg __411951_411951;
   reg _411952_411952 ; 
   reg __411952_411952;
   reg _411953_411953 ; 
   reg __411953_411953;
   reg _411954_411954 ; 
   reg __411954_411954;
   reg _411955_411955 ; 
   reg __411955_411955;
   reg _411956_411956 ; 
   reg __411956_411956;
   reg _411957_411957 ; 
   reg __411957_411957;
   reg _411958_411958 ; 
   reg __411958_411958;
   reg _411959_411959 ; 
   reg __411959_411959;
   reg _411960_411960 ; 
   reg __411960_411960;
   reg _411961_411961 ; 
   reg __411961_411961;
   reg _411962_411962 ; 
   reg __411962_411962;
   reg _411963_411963 ; 
   reg __411963_411963;
   reg _411964_411964 ; 
   reg __411964_411964;
   reg _411965_411965 ; 
   reg __411965_411965;
   reg _411966_411966 ; 
   reg __411966_411966;
   reg _411967_411967 ; 
   reg __411967_411967;
   reg _411968_411968 ; 
   reg __411968_411968;
   reg _411969_411969 ; 
   reg __411969_411969;
   reg _411970_411970 ; 
   reg __411970_411970;
   reg _411971_411971 ; 
   reg __411971_411971;
   reg _411972_411972 ; 
   reg __411972_411972;
   reg _411973_411973 ; 
   reg __411973_411973;
   reg _411974_411974 ; 
   reg __411974_411974;
   reg _411975_411975 ; 
   reg __411975_411975;
   reg _411976_411976 ; 
   reg __411976_411976;
   reg _411977_411977 ; 
   reg __411977_411977;
   reg _411978_411978 ; 
   reg __411978_411978;
   reg _411979_411979 ; 
   reg __411979_411979;
   reg _411980_411980 ; 
   reg __411980_411980;
   reg _411981_411981 ; 
   reg __411981_411981;
   reg _411982_411982 ; 
   reg __411982_411982;
   reg _411983_411983 ; 
   reg __411983_411983;
   reg _411984_411984 ; 
   reg __411984_411984;
   reg _411985_411985 ; 
   reg __411985_411985;
   reg _411986_411986 ; 
   reg __411986_411986;
   reg _411987_411987 ; 
   reg __411987_411987;
   reg _411988_411988 ; 
   reg __411988_411988;
   reg _411989_411989 ; 
   reg __411989_411989;
   reg _411990_411990 ; 
   reg __411990_411990;
   reg _411991_411991 ; 
   reg __411991_411991;
   reg _411992_411992 ; 
   reg __411992_411992;
   reg _411993_411993 ; 
   reg __411993_411993;
   reg _411994_411994 ; 
   reg __411994_411994;
   reg _411995_411995 ; 
   reg __411995_411995;
   reg _411996_411996 ; 
   reg __411996_411996;
   reg _411997_411997 ; 
   reg __411997_411997;
   reg _411998_411998 ; 
   reg __411998_411998;
   reg _411999_411999 ; 
   reg __411999_411999;
   reg _412000_412000 ; 
   reg __412000_412000;
   reg _412001_412001 ; 
   reg __412001_412001;
   reg _412002_412002 ; 
   reg __412002_412002;
   reg _412003_412003 ; 
   reg __412003_412003;
   reg _412004_412004 ; 
   reg __412004_412004;
   reg _412005_412005 ; 
   reg __412005_412005;
   reg _412006_412006 ; 
   reg __412006_412006;
   reg _412007_412007 ; 
   reg __412007_412007;
   reg _412008_412008 ; 
   reg __412008_412008;
   reg _412009_412009 ; 
   reg __412009_412009;
   reg _412010_412010 ; 
   reg __412010_412010;
   reg _412011_412011 ; 
   reg __412011_412011;
   reg _412012_412012 ; 
   reg __412012_412012;
   reg _412013_412013 ; 
   reg __412013_412013;
   reg _412014_412014 ; 
   reg __412014_412014;
   reg _412015_412015 ; 
   reg __412015_412015;
   reg _412016_412016 ; 
   reg __412016_412016;
   reg _412017_412017 ; 
   reg __412017_412017;
   reg _412018_412018 ; 
   reg __412018_412018;
   reg _412019_412019 ; 
   reg __412019_412019;
   reg _412020_412020 ; 
   reg __412020_412020;
   reg _412021_412021 ; 
   reg __412021_412021;
   reg _412022_412022 ; 
   reg __412022_412022;
   reg _412023_412023 ; 
   reg __412023_412023;
   reg _412024_412024 ; 
   reg __412024_412024;
   reg _412025_412025 ; 
   reg __412025_412025;
   reg _412026_412026 ; 
   reg __412026_412026;
   reg _412027_412027 ; 
   reg __412027_412027;
   reg _412028_412028 ; 
   reg __412028_412028;
   reg _412029_412029 ; 
   reg __412029_412029;
   reg _412030_412030 ; 
   reg __412030_412030;
   reg _412031_412031 ; 
   reg __412031_412031;
   reg _412032_412032 ; 
   reg __412032_412032;
   reg _412033_412033 ; 
   reg __412033_412033;
   reg _412034_412034 ; 
   reg __412034_412034;
   reg _412035_412035 ; 
   reg __412035_412035;
   reg _412036_412036 ; 
   reg __412036_412036;
   reg _412037_412037 ; 
   reg __412037_412037;
   reg _412038_412038 ; 
   reg __412038_412038;
   reg _412039_412039 ; 
   reg __412039_412039;
   reg _412040_412040 ; 
   reg __412040_412040;
   reg _412041_412041 ; 
   reg __412041_412041;
   reg _412042_412042 ; 
   reg __412042_412042;
   reg _412043_412043 ; 
   reg __412043_412043;
   reg _412044_412044 ; 
   reg __412044_412044;
   reg _412045_412045 ; 
   reg __412045_412045;
   reg _412046_412046 ; 
   reg __412046_412046;
   reg _412047_412047 ; 
   reg __412047_412047;
   reg _412048_412048 ; 
   reg __412048_412048;
   reg _412049_412049 ; 
   reg __412049_412049;
   reg _412050_412050 ; 
   reg __412050_412050;
   reg _412051_412051 ; 
   reg __412051_412051;
   reg _412052_412052 ; 
   reg __412052_412052;
   reg _412053_412053 ; 
   reg __412053_412053;
   reg _412054_412054 ; 
   reg __412054_412054;
   reg _412055_412055 ; 
   reg __412055_412055;
   reg _412056_412056 ; 
   reg __412056_412056;
   reg _412057_412057 ; 
   reg __412057_412057;
   reg _412058_412058 ; 
   reg __412058_412058;
   reg _412059_412059 ; 
   reg __412059_412059;
   reg _412060_412060 ; 
   reg __412060_412060;
   reg _412061_412061 ; 
   reg __412061_412061;
   reg _412062_412062 ; 
   reg __412062_412062;
   reg _412063_412063 ; 
   reg __412063_412063;
   reg _412064_412064 ; 
   reg __412064_412064;
   reg _412065_412065 ; 
   reg __412065_412065;
   reg _412066_412066 ; 
   reg __412066_412066;
   reg _412067_412067 ; 
   reg __412067_412067;
   reg _412068_412068 ; 
   reg __412068_412068;
   reg _412069_412069 ; 
   reg __412069_412069;
   reg _412070_412070 ; 
   reg __412070_412070;
   reg _412071_412071 ; 
   reg __412071_412071;
   reg _412072_412072 ; 
   reg __412072_412072;
   reg _412073_412073 ; 
   reg __412073_412073;
   reg _412074_412074 ; 
   reg __412074_412074;
   reg _412075_412075 ; 
   reg __412075_412075;
   reg _412076_412076 ; 
   reg __412076_412076;
   reg _412077_412077 ; 
   reg __412077_412077;
   reg _412078_412078 ; 
   reg __412078_412078;
   reg _412079_412079 ; 
   reg __412079_412079;
   reg _412080_412080 ; 
   reg __412080_412080;
   reg _412081_412081 ; 
   reg __412081_412081;
   reg _412082_412082 ; 
   reg __412082_412082;
   reg _412083_412083 ; 
   reg __412083_412083;
   reg _412084_412084 ; 
   reg __412084_412084;
   reg _412085_412085 ; 
   reg __412085_412085;
   reg _412086_412086 ; 
   reg __412086_412086;
   reg _412087_412087 ; 
   reg __412087_412087;
   reg _412088_412088 ; 
   reg __412088_412088;
   reg _412089_412089 ; 
   reg __412089_412089;
   reg _412090_412090 ; 
   reg __412090_412090;
   reg _412091_412091 ; 
   reg __412091_412091;
   reg _412092_412092 ; 
   reg __412092_412092;
   reg _412093_412093 ; 
   reg __412093_412093;
   reg _412094_412094 ; 
   reg __412094_412094;
   reg _412095_412095 ; 
   reg __412095_412095;
   reg _412096_412096 ; 
   reg __412096_412096;
   reg _412097_412097 ; 
   reg __412097_412097;
   reg _412098_412098 ; 
   reg __412098_412098;
   reg _412099_412099 ; 
   reg __412099_412099;
   reg _412100_412100 ; 
   reg __412100_412100;
   reg _412101_412101 ; 
   reg __412101_412101;
   reg _412102_412102 ; 
   reg __412102_412102;
   reg _412103_412103 ; 
   reg __412103_412103;
   reg _412104_412104 ; 
   reg __412104_412104;
   reg _412105_412105 ; 
   reg __412105_412105;
   reg _412106_412106 ; 
   reg __412106_412106;
   reg _412107_412107 ; 
   reg __412107_412107;
   reg _412108_412108 ; 
   reg __412108_412108;
   reg _412109_412109 ; 
   reg __412109_412109;
   reg _412110_412110 ; 
   reg __412110_412110;
   reg _412111_412111 ; 
   reg __412111_412111;
   reg _412112_412112 ; 
   reg __412112_412112;
   reg _412113_412113 ; 
   reg __412113_412113;
   reg _412114_412114 ; 
   reg __412114_412114;
   reg _412115_412115 ; 
   reg __412115_412115;
   reg _412116_412116 ; 
   reg __412116_412116;
   reg _412117_412117 ; 
   reg __412117_412117;
   reg _412118_412118 ; 
   reg __412118_412118;
   reg _412119_412119 ; 
   reg __412119_412119;
   reg _412120_412120 ; 
   reg __412120_412120;
   reg _412121_412121 ; 
   reg __412121_412121;
   reg _412122_412122 ; 
   reg __412122_412122;
   reg _412123_412123 ; 
   reg __412123_412123;
   reg _412124_412124 ; 
   reg __412124_412124;
   reg _412125_412125 ; 
   reg __412125_412125;
   reg _412126_412126 ; 
   reg __412126_412126;
   reg _412127_412127 ; 
   reg __412127_412127;
   reg _412128_412128 ; 
   reg __412128_412128;
   reg _412129_412129 ; 
   reg __412129_412129;
   reg _412130_412130 ; 
   reg __412130_412130;
   reg _412131_412131 ; 
   reg __412131_412131;
   reg _412132_412132 ; 
   reg __412132_412132;
   reg _412133_412133 ; 
   reg __412133_412133;
   reg _412134_412134 ; 
   reg __412134_412134;
   reg _412135_412135 ; 
   reg __412135_412135;
   reg _412136_412136 ; 
   reg __412136_412136;
   reg _412137_412137 ; 
   reg __412137_412137;
   reg _412138_412138 ; 
   reg __412138_412138;
   reg _412139_412139 ; 
   reg __412139_412139;
   reg _412140_412140 ; 
   reg __412140_412140;
   reg _412141_412141 ; 
   reg __412141_412141;
   reg _412142_412142 ; 
   reg __412142_412142;
   reg _412143_412143 ; 
   reg __412143_412143;
   reg _412144_412144 ; 
   reg __412144_412144;
   reg _412145_412145 ; 
   reg __412145_412145;
   reg _412146_412146 ; 
   reg __412146_412146;
   reg _412147_412147 ; 
   reg __412147_412147;
   reg _412148_412148 ; 
   reg __412148_412148;
   reg _412149_412149 ; 
   reg __412149_412149;
   reg _412150_412150 ; 
   reg __412150_412150;
   reg _412151_412151 ; 
   reg __412151_412151;
   reg _412152_412152 ; 
   reg __412152_412152;
   reg _412153_412153 ; 
   reg __412153_412153;
   reg _412154_412154 ; 
   reg __412154_412154;
   reg _412155_412155 ; 
   reg __412155_412155;
   reg _412156_412156 ; 
   reg __412156_412156;
   reg _412157_412157 ; 
   reg __412157_412157;
   reg _412158_412158 ; 
   reg __412158_412158;
   reg _412159_412159 ; 
   reg __412159_412159;
   reg _412160_412160 ; 
   reg __412160_412160;
   reg _412161_412161 ; 
   reg __412161_412161;
   reg _412162_412162 ; 
   reg __412162_412162;
   reg _412163_412163 ; 
   reg __412163_412163;
   reg _412164_412164 ; 
   reg __412164_412164;
   reg _412165_412165 ; 
   reg __412165_412165;
   reg _412166_412166 ; 
   reg __412166_412166;
   reg _412167_412167 ; 
   reg __412167_412167;
   reg _412168_412168 ; 
   reg __412168_412168;
   reg _412169_412169 ; 
   reg __412169_412169;
   reg _412170_412170 ; 
   reg __412170_412170;
   reg _412171_412171 ; 
   reg __412171_412171;
   reg _412172_412172 ; 
   reg __412172_412172;
   reg _412173_412173 ; 
   reg __412173_412173;
   reg _412174_412174 ; 
   reg __412174_412174;
   reg _412175_412175 ; 
   reg __412175_412175;
   reg _412176_412176 ; 
   reg __412176_412176;
   reg _412177_412177 ; 
   reg __412177_412177;
   reg _412178_412178 ; 
   reg __412178_412178;
   reg _412179_412179 ; 
   reg __412179_412179;
   reg _412180_412180 ; 
   reg __412180_412180;
   reg _412181_412181 ; 
   reg __412181_412181;
   reg _412182_412182 ; 
   reg __412182_412182;
   reg _412183_412183 ; 
   reg __412183_412183;
   reg _412184_412184 ; 
   reg __412184_412184;
   reg _412185_412185 ; 
   reg __412185_412185;
   reg _412186_412186 ; 
   reg __412186_412186;
   reg _412187_412187 ; 
   reg __412187_412187;
   reg _412188_412188 ; 
   reg __412188_412188;
   reg _412189_412189 ; 
   reg __412189_412189;
   reg _412190_412190 ; 
   reg __412190_412190;
   reg _412191_412191 ; 
   reg __412191_412191;
   reg _412192_412192 ; 
   reg __412192_412192;
   reg _412193_412193 ; 
   reg __412193_412193;
   reg _412194_412194 ; 
   reg __412194_412194;
   reg _412195_412195 ; 
   reg __412195_412195;
   reg _412196_412196 ; 
   reg __412196_412196;
   reg _412197_412197 ; 
   reg __412197_412197;
   reg _412198_412198 ; 
   reg __412198_412198;
   reg _412199_412199 ; 
   reg __412199_412199;
   reg _412200_412200 ; 
   reg __412200_412200;
   reg _412201_412201 ; 
   reg __412201_412201;
   reg _412202_412202 ; 
   reg __412202_412202;
   reg _412203_412203 ; 
   reg __412203_412203;
   reg _412204_412204 ; 
   reg __412204_412204;
   reg _412205_412205 ; 
   reg __412205_412205;
   reg _412206_412206 ; 
   reg __412206_412206;
   reg _412207_412207 ; 
   reg __412207_412207;
   reg _412208_412208 ; 
   reg __412208_412208;
   reg _412209_412209 ; 
   reg __412209_412209;
   reg _412210_412210 ; 
   reg __412210_412210;
   reg _412211_412211 ; 
   reg __412211_412211;
   reg _412212_412212 ; 
   reg __412212_412212;
   reg _412213_412213 ; 
   reg __412213_412213;
   reg _412214_412214 ; 
   reg __412214_412214;
   reg _412215_412215 ; 
   reg __412215_412215;
   reg _412216_412216 ; 
   reg __412216_412216;
   reg _412217_412217 ; 
   reg __412217_412217;
   reg _412218_412218 ; 
   reg __412218_412218;
   reg _412219_412219 ; 
   reg __412219_412219;
   reg _412220_412220 ; 
   reg __412220_412220;
   reg _412221_412221 ; 
   reg __412221_412221;
   reg _412222_412222 ; 
   reg __412222_412222;
   reg _412223_412223 ; 
   reg __412223_412223;
   reg _412224_412224 ; 
   reg __412224_412224;
   reg _412225_412225 ; 
   reg __412225_412225;
   reg _412226_412226 ; 
   reg __412226_412226;
   reg _412227_412227 ; 
   reg __412227_412227;
   reg _412228_412228 ; 
   reg __412228_412228;
   reg _412229_412229 ; 
   reg __412229_412229;
   reg _412230_412230 ; 
   reg __412230_412230;
   reg _412231_412231 ; 
   reg __412231_412231;
   reg _412232_412232 ; 
   reg __412232_412232;
   reg _412233_412233 ; 
   reg __412233_412233;
   reg _412234_412234 ; 
   reg __412234_412234;
   reg _412235_412235 ; 
   reg __412235_412235;
   reg _412236_412236 ; 
   reg __412236_412236;
   reg _412237_412237 ; 
   reg __412237_412237;
   reg _412238_412238 ; 
   reg __412238_412238;
   reg _412239_412239 ; 
   reg __412239_412239;
   reg _412240_412240 ; 
   reg __412240_412240;
   reg _412241_412241 ; 
   reg __412241_412241;
   reg _412242_412242 ; 
   reg __412242_412242;
   reg _412243_412243 ; 
   reg __412243_412243;
   reg _412244_412244 ; 
   reg __412244_412244;
   reg _412245_412245 ; 
   reg __412245_412245;
   reg _412246_412246 ; 
   reg __412246_412246;
   reg _412247_412247 ; 
   reg __412247_412247;
   reg _412248_412248 ; 
   reg __412248_412248;
   reg _412249_412249 ; 
   reg __412249_412249;
   reg _412250_412250 ; 
   reg __412250_412250;
   reg _412251_412251 ; 
   reg __412251_412251;
   reg _412252_412252 ; 
   reg __412252_412252;
   reg _412253_412253 ; 
   reg __412253_412253;
   reg _412254_412254 ; 
   reg __412254_412254;
   reg _412255_412255 ; 
   reg __412255_412255;
   reg _412256_412256 ; 
   reg __412256_412256;
   reg _412257_412257 ; 
   reg __412257_412257;
   reg _412258_412258 ; 
   reg __412258_412258;
   reg _412259_412259 ; 
   reg __412259_412259;
   reg _412260_412260 ; 
   reg __412260_412260;
   reg _412261_412261 ; 
   reg __412261_412261;
   reg _412262_412262 ; 
   reg __412262_412262;
   reg _412263_412263 ; 
   reg __412263_412263;
   reg _412264_412264 ; 
   reg __412264_412264;
   reg _412265_412265 ; 
   reg __412265_412265;
   reg _412266_412266 ; 
   reg __412266_412266;
   reg _412267_412267 ; 
   reg __412267_412267;
   reg _412268_412268 ; 
   reg __412268_412268;
   reg _412269_412269 ; 
   reg __412269_412269;
   reg _412270_412270 ; 
   reg __412270_412270;
   reg _412271_412271 ; 
   reg __412271_412271;
   reg _412272_412272 ; 
   reg __412272_412272;
   reg _412273_412273 ; 
   reg __412273_412273;
   reg _412274_412274 ; 
   reg __412274_412274;
   reg _412275_412275 ; 
   reg __412275_412275;
   reg _412276_412276 ; 
   reg __412276_412276;
   reg _412277_412277 ; 
   reg __412277_412277;
   reg _412278_412278 ; 
   reg __412278_412278;
   reg _412279_412279 ; 
   reg __412279_412279;
   reg _412280_412280 ; 
   reg __412280_412280;
   reg _412281_412281 ; 
   reg __412281_412281;
   reg _412282_412282 ; 
   reg __412282_412282;
   reg _412283_412283 ; 
   reg __412283_412283;
   reg _412284_412284 ; 
   reg __412284_412284;
   reg _412285_412285 ; 
   reg __412285_412285;
   reg _412286_412286 ; 
   reg __412286_412286;
   reg _412287_412287 ; 
   reg __412287_412287;
   reg _412288_412288 ; 
   reg __412288_412288;
   reg _412289_412289 ; 
   reg __412289_412289;
   reg _412290_412290 ; 
   reg __412290_412290;
   reg _412291_412291 ; 
   reg __412291_412291;
   reg _412292_412292 ; 
   reg __412292_412292;
   reg _412293_412293 ; 
   reg __412293_412293;
   reg _412294_412294 ; 
   reg __412294_412294;
   reg _412295_412295 ; 
   reg __412295_412295;
   reg _412296_412296 ; 
   reg __412296_412296;
   reg _412297_412297 ; 
   reg __412297_412297;
   reg _412298_412298 ; 
   reg __412298_412298;
   reg _412299_412299 ; 
   reg __412299_412299;
   reg _412300_412300 ; 
   reg __412300_412300;
   reg _412301_412301 ; 
   reg __412301_412301;
   reg _412302_412302 ; 
   reg __412302_412302;
   reg _412303_412303 ; 
   reg __412303_412303;
   reg _412304_412304 ; 
   reg __412304_412304;
   reg _412305_412305 ; 
   reg __412305_412305;
   reg _412306_412306 ; 
   reg __412306_412306;
   reg _412307_412307 ; 
   reg __412307_412307;
   reg _412308_412308 ; 
   reg __412308_412308;
   reg _412309_412309 ; 
   reg __412309_412309;
   reg _412310_412310 ; 
   reg __412310_412310;
   reg _412311_412311 ; 
   reg __412311_412311;
   reg _412312_412312 ; 
   reg __412312_412312;
   reg _412313_412313 ; 
   reg __412313_412313;
   reg _412314_412314 ; 
   reg __412314_412314;
   reg _412315_412315 ; 
   reg __412315_412315;
   reg _412316_412316 ; 
   reg __412316_412316;
   reg _412317_412317 ; 
   reg __412317_412317;
   reg _412318_412318 ; 
   reg __412318_412318;
   reg _412319_412319 ; 
   reg __412319_412319;
   reg _412320_412320 ; 
   reg __412320_412320;
   reg _412321_412321 ; 
   reg __412321_412321;
   reg _412322_412322 ; 
   reg __412322_412322;
   reg _412323_412323 ; 
   reg __412323_412323;
   reg _412324_412324 ; 
   reg __412324_412324;
   reg _412325_412325 ; 
   reg __412325_412325;
   reg _412326_412326 ; 
   reg __412326_412326;
   reg _412327_412327 ; 
   reg __412327_412327;
   reg _412328_412328 ; 
   reg __412328_412328;
   reg _412329_412329 ; 
   reg __412329_412329;
   reg _412330_412330 ; 
   reg __412330_412330;
   reg _412331_412331 ; 
   reg __412331_412331;
   reg _412332_412332 ; 
   reg __412332_412332;
   reg _412333_412333 ; 
   reg __412333_412333;
   reg _412334_412334 ; 
   reg __412334_412334;
   reg _412335_412335 ; 
   reg __412335_412335;
   reg _412336_412336 ; 
   reg __412336_412336;
   reg _412337_412337 ; 
   reg __412337_412337;
   reg _412338_412338 ; 
   reg __412338_412338;
   reg _412339_412339 ; 
   reg __412339_412339;
   reg _412340_412340 ; 
   reg __412340_412340;
   reg _412341_412341 ; 
   reg __412341_412341;
   reg _412342_412342 ; 
   reg __412342_412342;
   reg _412343_412343 ; 
   reg __412343_412343;
   reg _412344_412344 ; 
   reg __412344_412344;
   reg _412345_412345 ; 
   reg __412345_412345;
   reg _412346_412346 ; 
   reg __412346_412346;
   reg _412347_412347 ; 
   reg __412347_412347;
   reg _412348_412348 ; 
   reg __412348_412348;
   reg _412349_412349 ; 
   reg __412349_412349;
   reg _412350_412350 ; 
   reg __412350_412350;
   reg _412351_412351 ; 
   reg __412351_412351;
   reg _412352_412352 ; 
   reg __412352_412352;
   reg _412353_412353 ; 
   reg __412353_412353;
   reg _412354_412354 ; 
   reg __412354_412354;
   reg _412355_412355 ; 
   reg __412355_412355;
   reg _412356_412356 ; 
   reg __412356_412356;
   reg _412357_412357 ; 
   reg __412357_412357;
   reg _412358_412358 ; 
   reg __412358_412358;
   reg _412359_412359 ; 
   reg __412359_412359;
   reg _412360_412360 ; 
   reg __412360_412360;
   reg _412361_412361 ; 
   reg __412361_412361;
   reg _412362_412362 ; 
   reg __412362_412362;
   reg _412363_412363 ; 
   reg __412363_412363;
   reg _412364_412364 ; 
   reg __412364_412364;
   reg _412365_412365 ; 
   reg __412365_412365;
   reg _412366_412366 ; 
   reg __412366_412366;
   reg _412367_412367 ; 
   reg __412367_412367;
   reg _412368_412368 ; 
   reg __412368_412368;
   reg _412369_412369 ; 
   reg __412369_412369;
   reg _412370_412370 ; 
   reg __412370_412370;
   reg _412371_412371 ; 
   reg __412371_412371;
   reg _412372_412372 ; 
   reg __412372_412372;
   reg _412373_412373 ; 
   reg __412373_412373;
   reg _412374_412374 ; 
   reg __412374_412374;
   reg _412375_412375 ; 
   reg __412375_412375;
   reg _412376_412376 ; 
   reg __412376_412376;
   reg _412377_412377 ; 
   reg __412377_412377;
   reg _412378_412378 ; 
   reg __412378_412378;
   reg _412379_412379 ; 
   reg __412379_412379;
   reg _412380_412380 ; 
   reg __412380_412380;
   reg _412381_412381 ; 
   reg __412381_412381;
   reg _412382_412382 ; 
   reg __412382_412382;
   reg _412383_412383 ; 
   reg __412383_412383;
   reg _412384_412384 ; 
   reg __412384_412384;
   reg _412385_412385 ; 
   reg __412385_412385;
   reg _412386_412386 ; 
   reg __412386_412386;
   reg _412387_412387 ; 
   reg __412387_412387;
   reg _412388_412388 ; 
   reg __412388_412388;
   reg _412389_412389 ; 
   reg __412389_412389;
   reg _412390_412390 ; 
   reg __412390_412390;
   reg _412391_412391 ; 
   reg __412391_412391;
   reg _412392_412392 ; 
   reg __412392_412392;
   reg _412393_412393 ; 
   reg __412393_412393;
   reg _412394_412394 ; 
   reg __412394_412394;
   reg _412395_412395 ; 
   reg __412395_412395;
   reg _412396_412396 ; 
   reg __412396_412396;
   reg _412397_412397 ; 
   reg __412397_412397;
   reg _412398_412398 ; 
   reg __412398_412398;
   reg _412399_412399 ; 
   reg __412399_412399;
   reg _412400_412400 ; 
   reg __412400_412400;
   reg _412401_412401 ; 
   reg __412401_412401;
   reg _412402_412402 ; 
   reg __412402_412402;
   reg _412403_412403 ; 
   reg __412403_412403;
   reg _412404_412404 ; 
   reg __412404_412404;
   reg _412405_412405 ; 
   reg __412405_412405;
   reg _412406_412406 ; 
   reg __412406_412406;
   reg _412407_412407 ; 
   reg __412407_412407;
   reg _412408_412408 ; 
   reg __412408_412408;
   reg _412409_412409 ; 
   reg __412409_412409;
   reg _412410_412410 ; 
   reg __412410_412410;
   reg _412411_412411 ; 
   reg __412411_412411;
   reg _412412_412412 ; 
   reg __412412_412412;
   reg _412413_412413 ; 
   reg __412413_412413;
   reg _412414_412414 ; 
   reg __412414_412414;
   reg _412415_412415 ; 
   reg __412415_412415;
   reg _412416_412416 ; 
   reg __412416_412416;
   reg _412417_412417 ; 
   reg __412417_412417;
   reg _412418_412418 ; 
   reg __412418_412418;
   reg _412419_412419 ; 
   reg __412419_412419;
   reg _412420_412420 ; 
   reg __412420_412420;
   reg _412421_412421 ; 
   reg __412421_412421;
   reg _412422_412422 ; 
   reg __412422_412422;
   reg _412423_412423 ; 
   reg __412423_412423;
   reg _412424_412424 ; 
   reg __412424_412424;
   reg _412425_412425 ; 
   reg __412425_412425;
   reg _412426_412426 ; 
   reg __412426_412426;
   reg _412427_412427 ; 
   reg __412427_412427;
   reg _412428_412428 ; 
   reg __412428_412428;
   reg _412429_412429 ; 
   reg __412429_412429;
   reg _412430_412430 ; 
   reg __412430_412430;
   reg _412431_412431 ; 
   reg __412431_412431;
   reg _412432_412432 ; 
   reg __412432_412432;
   reg _412433_412433 ; 
   reg __412433_412433;
   reg _412434_412434 ; 
   reg __412434_412434;
   reg _412435_412435 ; 
   reg __412435_412435;
   reg _412436_412436 ; 
   reg __412436_412436;
   reg _412437_412437 ; 
   reg __412437_412437;
   reg _412438_412438 ; 
   reg __412438_412438;
   reg _412439_412439 ; 
   reg __412439_412439;
   reg _412440_412440 ; 
   reg __412440_412440;
   reg _412441_412441 ; 
   reg __412441_412441;
   reg _412442_412442 ; 
   reg __412442_412442;
   reg _412443_412443 ; 
   reg __412443_412443;
   reg _412444_412444 ; 
   reg __412444_412444;
   reg _412445_412445 ; 
   reg __412445_412445;
   reg _412446_412446 ; 
   reg __412446_412446;
   reg _412447_412447 ; 
   reg __412447_412447;
   reg _412448_412448 ; 
   reg __412448_412448;
   reg _412449_412449 ; 
   reg __412449_412449;
   reg _412450_412450 ; 
   reg __412450_412450;
   reg _412451_412451 ; 
   reg __412451_412451;
   reg _412452_412452 ; 
   reg __412452_412452;
   reg _412453_412453 ; 
   reg __412453_412453;
   reg _412454_412454 ; 
   reg __412454_412454;
   reg _412455_412455 ; 
   reg __412455_412455;
   reg _412456_412456 ; 
   reg __412456_412456;
   reg _412457_412457 ; 
   reg __412457_412457;
   reg _412458_412458 ; 
   reg __412458_412458;
   reg _412459_412459 ; 
   reg __412459_412459;
   reg _412460_412460 ; 
   reg __412460_412460;
   reg _412461_412461 ; 
   reg __412461_412461;
   reg _412462_412462 ; 
   reg __412462_412462;
   reg _412463_412463 ; 
   reg __412463_412463;
   reg _412464_412464 ; 
   reg __412464_412464;
   reg _412465_412465 ; 
   reg __412465_412465;
   reg _412466_412466 ; 
   reg __412466_412466;
   reg _412467_412467 ; 
   reg __412467_412467;
   reg _412468_412468 ; 
   reg __412468_412468;
   reg _412469_412469 ; 
   reg __412469_412469;
   reg _412470_412470 ; 
   reg __412470_412470;
   reg _412471_412471 ; 
   reg __412471_412471;
   reg _412472_412472 ; 
   reg __412472_412472;
   reg _412473_412473 ; 
   reg __412473_412473;
   reg _412474_412474 ; 
   reg __412474_412474;
   reg _412475_412475 ; 
   reg __412475_412475;
   reg _412476_412476 ; 
   reg __412476_412476;
   reg _412477_412477 ; 
   reg __412477_412477;
   reg _412478_412478 ; 
   reg __412478_412478;
   reg _412479_412479 ; 
   reg __412479_412479;
   reg _412480_412480 ; 
   reg __412480_412480;
   reg _412481_412481 ; 
   reg __412481_412481;
   reg _412482_412482 ; 
   reg __412482_412482;
   reg _412483_412483 ; 
   reg __412483_412483;
   reg _412484_412484 ; 
   reg __412484_412484;
   reg _412485_412485 ; 
   reg __412485_412485;
   reg _412486_412486 ; 
   reg __412486_412486;
   reg _412487_412487 ; 
   reg __412487_412487;
   reg _412488_412488 ; 
   reg __412488_412488;
   reg _412489_412489 ; 
   reg __412489_412489;
   reg _412490_412490 ; 
   reg __412490_412490;
   reg _412491_412491 ; 
   reg __412491_412491;
   reg _412492_412492 ; 
   reg __412492_412492;
   reg _412493_412493 ; 
   reg __412493_412493;
   reg _412494_412494 ; 
   reg __412494_412494;
   reg _412495_412495 ; 
   reg __412495_412495;
   reg _412496_412496 ; 
   reg __412496_412496;
   reg _412497_412497 ; 
   reg __412497_412497;
   reg _412498_412498 ; 
   reg __412498_412498;
   reg _412499_412499 ; 
   reg __412499_412499;
   reg _412500_412500 ; 
   reg __412500_412500;
   reg _412501_412501 ; 
   reg __412501_412501;
   reg _412502_412502 ; 
   reg __412502_412502;
   reg _412503_412503 ; 
   reg __412503_412503;
   reg _412504_412504 ; 
   reg __412504_412504;
   reg _412505_412505 ; 
   reg __412505_412505;
   reg _412506_412506 ; 
   reg __412506_412506;
   reg _412507_412507 ; 
   reg __412507_412507;
   reg _412508_412508 ; 
   reg __412508_412508;
   reg _412509_412509 ; 
   reg __412509_412509;
   reg _412510_412510 ; 
   reg __412510_412510;
   reg _412511_412511 ; 
   reg __412511_412511;
   reg _412512_412512 ; 
   reg __412512_412512;
   reg _412513_412513 ; 
   reg __412513_412513;
   reg _412514_412514 ; 
   reg __412514_412514;
   reg _412515_412515 ; 
   reg __412515_412515;
   reg _412516_412516 ; 
   reg __412516_412516;
   reg _412517_412517 ; 
   reg __412517_412517;
   reg _412518_412518 ; 
   reg __412518_412518;
   reg _412519_412519 ; 
   reg __412519_412519;
   reg _412520_412520 ; 
   reg __412520_412520;
   reg _412521_412521 ; 
   reg __412521_412521;
   reg _412522_412522 ; 
   reg __412522_412522;
   reg _412523_412523 ; 
   reg __412523_412523;
   reg _412524_412524 ; 
   reg __412524_412524;
   reg _412525_412525 ; 
   reg __412525_412525;
   reg _412526_412526 ; 
   reg __412526_412526;
   reg _412527_412527 ; 
   reg __412527_412527;
   reg _412528_412528 ; 
   reg __412528_412528;
   reg _412529_412529 ; 
   reg __412529_412529;
   reg _412530_412530 ; 
   reg __412530_412530;
   reg _412531_412531 ; 
   reg __412531_412531;
   reg _412532_412532 ; 
   reg __412532_412532;
   reg _412533_412533 ; 
   reg __412533_412533;
   reg _412534_412534 ; 
   reg __412534_412534;
   reg _412535_412535 ; 
   reg __412535_412535;
   reg _412536_412536 ; 
   reg __412536_412536;
   reg _412537_412537 ; 
   reg __412537_412537;
   reg _412538_412538 ; 
   reg __412538_412538;
   reg _412539_412539 ; 
   reg __412539_412539;
   reg _412540_412540 ; 
   reg __412540_412540;
   reg _412541_412541 ; 
   reg __412541_412541;
   reg _412542_412542 ; 
   reg __412542_412542;
   reg _412543_412543 ; 
   reg __412543_412543;
   reg _412544_412544 ; 
   reg __412544_412544;
   reg _412545_412545 ; 
   reg __412545_412545;
   reg _412546_412546 ; 
   reg __412546_412546;
   reg _412547_412547 ; 
   reg __412547_412547;
   reg _412548_412548 ; 
   reg __412548_412548;
   reg _412549_412549 ; 
   reg __412549_412549;
   reg _412550_412550 ; 
   reg __412550_412550;
   reg _412551_412551 ; 
   reg __412551_412551;
   reg _412552_412552 ; 
   reg __412552_412552;
   reg _412553_412553 ; 
   reg __412553_412553;
   reg _412554_412554 ; 
   reg __412554_412554;
   reg _412555_412555 ; 
   reg __412555_412555;
   reg _412556_412556 ; 
   reg __412556_412556;
   reg _412557_412557 ; 
   reg __412557_412557;
   reg _412558_412558 ; 
   reg __412558_412558;
   reg _412559_412559 ; 
   reg __412559_412559;
   reg _412560_412560 ; 
   reg __412560_412560;
   reg _412561_412561 ; 
   reg __412561_412561;
   reg _412562_412562 ; 
   reg __412562_412562;
   reg _412563_412563 ; 
   reg __412563_412563;
   reg _412564_412564 ; 
   reg __412564_412564;
   reg _412565_412565 ; 
   reg __412565_412565;
   reg _412566_412566 ; 
   reg __412566_412566;
   reg _412567_412567 ; 
   reg __412567_412567;
   reg _412568_412568 ; 
   reg __412568_412568;
   reg _412569_412569 ; 
   reg __412569_412569;
   reg _412570_412570 ; 
   reg __412570_412570;
   reg _412571_412571 ; 
   reg __412571_412571;
   reg _412572_412572 ; 
   reg __412572_412572;
   reg _412573_412573 ; 
   reg __412573_412573;
   reg _412574_412574 ; 
   reg __412574_412574;
   reg _412575_412575 ; 
   reg __412575_412575;
   reg _412576_412576 ; 
   reg __412576_412576;
   reg _412577_412577 ; 
   reg __412577_412577;
   reg _412578_412578 ; 
   reg __412578_412578;
   reg _412579_412579 ; 
   reg __412579_412579;
   reg _412580_412580 ; 
   reg __412580_412580;
   reg _412581_412581 ; 
   reg __412581_412581;
   reg _412582_412582 ; 
   reg __412582_412582;
   reg _412583_412583 ; 
   reg __412583_412583;
   reg _412584_412584 ; 
   reg __412584_412584;
   reg _412585_412585 ; 
   reg __412585_412585;
   reg _412586_412586 ; 
   reg __412586_412586;
   reg _412587_412587 ; 
   reg __412587_412587;
   reg _412588_412588 ; 
   reg __412588_412588;
   reg _412589_412589 ; 
   reg __412589_412589;
   reg _412590_412590 ; 
   reg __412590_412590;
   reg _412591_412591 ; 
   reg __412591_412591;
   reg _412592_412592 ; 
   reg __412592_412592;
   reg _412593_412593 ; 
   reg __412593_412593;
   reg _412594_412594 ; 
   reg __412594_412594;
   reg _412595_412595 ; 
   reg __412595_412595;
   reg _412596_412596 ; 
   reg __412596_412596;
   reg _412597_412597 ; 
   reg __412597_412597;
   reg _412598_412598 ; 
   reg __412598_412598;
   reg _412599_412599 ; 
   reg __412599_412599;
   reg _412600_412600 ; 
   reg __412600_412600;
   reg _412601_412601 ; 
   reg __412601_412601;
   reg _412602_412602 ; 
   reg __412602_412602;
   reg _412603_412603 ; 
   reg __412603_412603;
   reg _412604_412604 ; 
   reg __412604_412604;
   reg _412605_412605 ; 
   reg __412605_412605;
   reg _412606_412606 ; 
   reg __412606_412606;
   reg _412607_412607 ; 
   reg __412607_412607;
   reg _412608_412608 ; 
   reg __412608_412608;
   reg _412609_412609 ; 
   reg __412609_412609;
   reg _412610_412610 ; 
   reg __412610_412610;
   reg _412611_412611 ; 
   reg __412611_412611;
   reg _412612_412612 ; 
   reg __412612_412612;
   reg _412613_412613 ; 
   reg __412613_412613;
   reg _412614_412614 ; 
   reg __412614_412614;
   reg _412615_412615 ; 
   reg __412615_412615;
   reg _412616_412616 ; 
   reg __412616_412616;
   reg _412617_412617 ; 
   reg __412617_412617;
   reg _412618_412618 ; 
   reg __412618_412618;
   reg _412619_412619 ; 
   reg __412619_412619;
   reg _412620_412620 ; 
   reg __412620_412620;
   reg _412621_412621 ; 
   reg __412621_412621;
   reg _412622_412622 ; 
   reg __412622_412622;
   reg _412623_412623 ; 
   reg __412623_412623;
   reg _412624_412624 ; 
   reg __412624_412624;
   reg _412625_412625 ; 
   reg __412625_412625;
   reg _412626_412626 ; 
   reg __412626_412626;
   reg _412627_412627 ; 
   reg __412627_412627;
   reg _412628_412628 ; 
   reg __412628_412628;
   reg _412629_412629 ; 
   reg __412629_412629;
   reg _412630_412630 ; 
   reg __412630_412630;
   reg _412631_412631 ; 
   reg __412631_412631;
   reg _412632_412632 ; 
   reg __412632_412632;
   reg _412633_412633 ; 
   reg __412633_412633;
   reg _412634_412634 ; 
   reg __412634_412634;
   reg _412635_412635 ; 
   reg __412635_412635;
   reg _412636_412636 ; 
   reg __412636_412636;
   reg _412637_412637 ; 
   reg __412637_412637;
   reg _412638_412638 ; 
   reg __412638_412638;
   reg _412639_412639 ; 
   reg __412639_412639;
   reg _412640_412640 ; 
   reg __412640_412640;
   reg _412641_412641 ; 
   reg __412641_412641;
   reg _412642_412642 ; 
   reg __412642_412642;
   reg _412643_412643 ; 
   reg __412643_412643;
   reg _412644_412644 ; 
   reg __412644_412644;
   reg _412645_412645 ; 
   reg __412645_412645;
   reg _412646_412646 ; 
   reg __412646_412646;
   reg _412647_412647 ; 
   reg __412647_412647;
   reg _412648_412648 ; 
   reg __412648_412648;
   reg _412649_412649 ; 
   reg __412649_412649;
   reg _412650_412650 ; 
   reg __412650_412650;
   reg _412651_412651 ; 
   reg __412651_412651;
   reg _412652_412652 ; 
   reg __412652_412652;
   reg _412653_412653 ; 
   reg __412653_412653;
   reg _412654_412654 ; 
   reg __412654_412654;
   reg _412655_412655 ; 
   reg __412655_412655;
   reg _412656_412656 ; 
   reg __412656_412656;
   reg _412657_412657 ; 
   reg __412657_412657;
   reg _412658_412658 ; 
   reg __412658_412658;
   reg _412659_412659 ; 
   reg __412659_412659;
   reg _412660_412660 ; 
   reg __412660_412660;
   reg _412661_412661 ; 
   reg __412661_412661;
   reg _412662_412662 ; 
   reg __412662_412662;
   reg _412663_412663 ; 
   reg __412663_412663;
   reg _412664_412664 ; 
   reg __412664_412664;
   reg _412665_412665 ; 
   reg __412665_412665;
   reg _412666_412666 ; 
   reg __412666_412666;
   reg _412667_412667 ; 
   reg __412667_412667;
   reg _412668_412668 ; 
   reg __412668_412668;
   reg _412669_412669 ; 
   reg __412669_412669;
   reg _412670_412670 ; 
   reg __412670_412670;
   reg _412671_412671 ; 
   reg __412671_412671;
   reg _412672_412672 ; 
   reg __412672_412672;
   reg _412673_412673 ; 
   reg __412673_412673;
   reg _412674_412674 ; 
   reg __412674_412674;
   reg _412675_412675 ; 
   reg __412675_412675;
   reg _412676_412676 ; 
   reg __412676_412676;
   reg _412677_412677 ; 
   reg __412677_412677;
   reg _412678_412678 ; 
   reg __412678_412678;
   reg _412679_412679 ; 
   reg __412679_412679;
   reg _412680_412680 ; 
   reg __412680_412680;
   reg _412681_412681 ; 
   reg __412681_412681;
   reg _412682_412682 ; 
   reg __412682_412682;
   reg _412683_412683 ; 
   reg __412683_412683;
   reg _412684_412684 ; 
   reg __412684_412684;
   reg _412685_412685 ; 
   reg __412685_412685;
   reg _412686_412686 ; 
   reg __412686_412686;
   reg _412687_412687 ; 
   reg __412687_412687;
   reg _412688_412688 ; 
   reg __412688_412688;
   reg _412689_412689 ; 
   reg __412689_412689;
   reg _412690_412690 ; 
   reg __412690_412690;
   reg _412691_412691 ; 
   reg __412691_412691;
   reg _412692_412692 ; 
   reg __412692_412692;
   reg _412693_412693 ; 
   reg __412693_412693;
   reg _412694_412694 ; 
   reg __412694_412694;
   reg _412695_412695 ; 
   reg __412695_412695;
   reg _412696_412696 ; 
   reg __412696_412696;
   reg _412697_412697 ; 
   reg __412697_412697;
   reg _412698_412698 ; 
   reg __412698_412698;
   reg _412699_412699 ; 
   reg __412699_412699;
   reg _412700_412700 ; 
   reg __412700_412700;
   reg _412701_412701 ; 
   reg __412701_412701;
   reg _412702_412702 ; 
   reg __412702_412702;
   reg _412703_412703 ; 
   reg __412703_412703;
   reg _412704_412704 ; 
   reg __412704_412704;
   reg _412705_412705 ; 
   reg __412705_412705;
   reg _412706_412706 ; 
   reg __412706_412706;
   reg _412707_412707 ; 
   reg __412707_412707;
   reg _412708_412708 ; 
   reg __412708_412708;
   reg _412709_412709 ; 
   reg __412709_412709;
   reg _412710_412710 ; 
   reg __412710_412710;
   reg _412711_412711 ; 
   reg __412711_412711;
   reg _412712_412712 ; 
   reg __412712_412712;
   reg _412713_412713 ; 
   reg __412713_412713;
   reg _412714_412714 ; 
   reg __412714_412714;
   reg _412715_412715 ; 
   reg __412715_412715;
   reg _412716_412716 ; 
   reg __412716_412716;
   reg _412717_412717 ; 
   reg __412717_412717;
   reg _412718_412718 ; 
   reg __412718_412718;
   reg _412719_412719 ; 
   reg __412719_412719;
   reg _412720_412720 ; 
   reg __412720_412720;
   reg _412721_412721 ; 
   reg __412721_412721;
   reg _412722_412722 ; 
   reg __412722_412722;
   reg _412723_412723 ; 
   reg __412723_412723;
   reg _412724_412724 ; 
   reg __412724_412724;
   reg _412725_412725 ; 
   reg __412725_412725;
   reg _412726_412726 ; 
   reg __412726_412726;
   reg _412727_412727 ; 
   reg __412727_412727;
   reg _412728_412728 ; 
   reg __412728_412728;
   reg _412729_412729 ; 
   reg __412729_412729;
   reg _412730_412730 ; 
   reg __412730_412730;
   reg _412731_412731 ; 
   reg __412731_412731;
   reg _412732_412732 ; 
   reg __412732_412732;
   reg _412733_412733 ; 
   reg __412733_412733;
   reg _412734_412734 ; 
   reg __412734_412734;
   reg _412735_412735 ; 
   reg __412735_412735;
   reg _412736_412736 ; 
   reg __412736_412736;
   reg _412737_412737 ; 
   reg __412737_412737;
   reg _412738_412738 ; 
   reg __412738_412738;
   reg _412739_412739 ; 
   reg __412739_412739;
   reg _412740_412740 ; 
   reg __412740_412740;
   reg _412741_412741 ; 
   reg __412741_412741;
   reg _412742_412742 ; 
   reg __412742_412742;
   reg _412743_412743 ; 
   reg __412743_412743;
   reg _412744_412744 ; 
   reg __412744_412744;
   reg _412745_412745 ; 
   reg __412745_412745;
   reg _412746_412746 ; 
   reg __412746_412746;
   reg _412747_412747 ; 
   reg __412747_412747;
   reg _412748_412748 ; 
   reg __412748_412748;
   reg _412749_412749 ; 
   reg __412749_412749;
   reg _412750_412750 ; 
   reg __412750_412750;
   reg _412751_412751 ; 
   reg __412751_412751;
   reg _412752_412752 ; 
   reg __412752_412752;
   reg _412753_412753 ; 
   reg __412753_412753;
   reg _412754_412754 ; 
   reg __412754_412754;
   reg _412755_412755 ; 
   reg __412755_412755;
   reg _412756_412756 ; 
   reg __412756_412756;
   reg _412757_412757 ; 
   reg __412757_412757;
   reg _412758_412758 ; 
   reg __412758_412758;
   reg _412759_412759 ; 
   reg __412759_412759;
   reg _412760_412760 ; 
   reg __412760_412760;
   reg _412761_412761 ; 
   reg __412761_412761;
   reg _412762_412762 ; 
   reg __412762_412762;
   reg _412763_412763 ; 
   reg __412763_412763;
   reg _412764_412764 ; 
   reg __412764_412764;
   reg _412765_412765 ; 
   reg __412765_412765;
   reg _412766_412766 ; 
   reg __412766_412766;
   reg _412767_412767 ; 
   reg __412767_412767;
   reg _412768_412768 ; 
   reg __412768_412768;
   reg _412769_412769 ; 
   reg __412769_412769;
   reg _412770_412770 ; 
   reg __412770_412770;
   reg _412771_412771 ; 
   reg __412771_412771;
   reg _412772_412772 ; 
   reg __412772_412772;
   reg _412773_412773 ; 
   reg __412773_412773;
   reg _412774_412774 ; 
   reg __412774_412774;
   reg _412775_412775 ; 
   reg __412775_412775;
   reg _412776_412776 ; 
   reg __412776_412776;
   reg _412777_412777 ; 
   reg __412777_412777;
   reg _412778_412778 ; 
   reg __412778_412778;
   reg _412779_412779 ; 
   reg __412779_412779;
   reg _412780_412780 ; 
   reg __412780_412780;
   reg _412781_412781 ; 
   reg __412781_412781;
   reg _412782_412782 ; 
   reg __412782_412782;
   reg _412783_412783 ; 
   reg __412783_412783;
   reg _412784_412784 ; 
   reg __412784_412784;
   reg _412785_412785 ; 
   reg __412785_412785;
   reg _412786_412786 ; 
   reg __412786_412786;
   reg _412787_412787 ; 
   reg __412787_412787;
   reg _412788_412788 ; 
   reg __412788_412788;
   reg _412789_412789 ; 
   reg __412789_412789;
   reg _412790_412790 ; 
   reg __412790_412790;
   reg _412791_412791 ; 
   reg __412791_412791;
   reg _412792_412792 ; 
   reg __412792_412792;
   reg _412793_412793 ; 
   reg __412793_412793;
   reg _412794_412794 ; 
   reg __412794_412794;
   reg _412795_412795 ; 
   reg __412795_412795;
   reg _412796_412796 ; 
   reg __412796_412796;
   reg _412797_412797 ; 
   reg __412797_412797;
   reg _412798_412798 ; 
   reg __412798_412798;
   reg _412799_412799 ; 
   reg __412799_412799;
   reg _412800_412800 ; 
   reg __412800_412800;
   reg _412801_412801 ; 
   reg __412801_412801;
   reg _412802_412802 ; 
   reg __412802_412802;
   reg _412803_412803 ; 
   reg __412803_412803;
   reg _412804_412804 ; 
   reg __412804_412804;
   reg _412805_412805 ; 
   reg __412805_412805;
   reg _412806_412806 ; 
   reg __412806_412806;
   reg _412807_412807 ; 
   reg __412807_412807;
   reg _412808_412808 ; 
   reg __412808_412808;
   reg _412809_412809 ; 
   reg __412809_412809;
   reg _412810_412810 ; 
   reg __412810_412810;
   reg _412811_412811 ; 
   reg __412811_412811;
   reg _412812_412812 ; 
   reg __412812_412812;
   reg _412813_412813 ; 
   reg __412813_412813;
   reg _412814_412814 ; 
   reg __412814_412814;
   reg _412815_412815 ; 
   reg __412815_412815;
   reg _412816_412816 ; 
   reg __412816_412816;
   reg _412817_412817 ; 
   reg __412817_412817;
   reg _412818_412818 ; 
   reg __412818_412818;
   reg _412819_412819 ; 
   reg __412819_412819;
   reg _412820_412820 ; 
   reg __412820_412820;
   reg _412821_412821 ; 
   reg __412821_412821;
   reg _412822_412822 ; 
   reg __412822_412822;
   reg _412823_412823 ; 
   reg __412823_412823;
   reg _412824_412824 ; 
   reg __412824_412824;
   reg _412825_412825 ; 
   reg __412825_412825;
   reg _412826_412826 ; 
   reg __412826_412826;
   reg _412827_412827 ; 
   reg __412827_412827;
   reg _412828_412828 ; 
   reg __412828_412828;
   reg _412829_412829 ; 
   reg __412829_412829;
   reg _412830_412830 ; 
   reg __412830_412830;
   reg _412831_412831 ; 
   reg __412831_412831;
   reg _412832_412832 ; 
   reg __412832_412832;
   reg _412833_412833 ; 
   reg __412833_412833;
   reg _412834_412834 ; 
   reg __412834_412834;
   reg _412835_412835 ; 
   reg __412835_412835;
   reg _412836_412836 ; 
   reg __412836_412836;
   reg _412837_412837 ; 
   reg __412837_412837;
   reg _412838_412838 ; 
   reg __412838_412838;
   reg _412839_412839 ; 
   reg __412839_412839;
   reg _412840_412840 ; 
   reg __412840_412840;
   reg _412841_412841 ; 
   reg __412841_412841;
   reg _412842_412842 ; 
   reg __412842_412842;
   reg _412843_412843 ; 
   reg __412843_412843;
   reg _412844_412844 ; 
   reg __412844_412844;
   reg _412845_412845 ; 
   reg __412845_412845;
   reg _412846_412846 ; 
   reg __412846_412846;
   reg _412847_412847 ; 
   reg __412847_412847;
   reg _412848_412848 ; 
   reg __412848_412848;
   reg _412849_412849 ; 
   reg __412849_412849;
   reg _412850_412850 ; 
   reg __412850_412850;
   reg _412851_412851 ; 
   reg __412851_412851;
   reg _412852_412852 ; 
   reg __412852_412852;
   reg _412853_412853 ; 
   reg __412853_412853;
   reg _412854_412854 ; 
   reg __412854_412854;
   reg _412855_412855 ; 
   reg __412855_412855;
   reg _412856_412856 ; 
   reg __412856_412856;
   reg _412857_412857 ; 
   reg __412857_412857;
   reg _412858_412858 ; 
   reg __412858_412858;
   reg _412859_412859 ; 
   reg __412859_412859;
   reg _412860_412860 ; 
   reg __412860_412860;
   reg _412861_412861 ; 
   reg __412861_412861;
   reg _412862_412862 ; 
   reg __412862_412862;
   reg _412863_412863 ; 
   reg __412863_412863;
   reg _412864_412864 ; 
   reg __412864_412864;
   reg _412865_412865 ; 
   reg __412865_412865;
   reg _412866_412866 ; 
   reg __412866_412866;
   reg _412867_412867 ; 
   reg __412867_412867;
   reg _412868_412868 ; 
   reg __412868_412868;
   reg _412869_412869 ; 
   reg __412869_412869;
   reg _412870_412870 ; 
   reg __412870_412870;
   reg _412871_412871 ; 
   reg __412871_412871;
   reg _412872_412872 ; 
   reg __412872_412872;
   reg _412873_412873 ; 
   reg __412873_412873;
   reg _412874_412874 ; 
   reg __412874_412874;
   reg _412875_412875 ; 
   reg __412875_412875;
   reg _412876_412876 ; 
   reg __412876_412876;
   reg _412877_412877 ; 
   reg __412877_412877;
   reg _412878_412878 ; 
   reg __412878_412878;
   reg _412879_412879 ; 
   reg __412879_412879;
   reg _412880_412880 ; 
   reg __412880_412880;
   reg _412881_412881 ; 
   reg __412881_412881;
   reg _412882_412882 ; 
   reg __412882_412882;
   reg _412883_412883 ; 
   reg __412883_412883;
   reg _412884_412884 ; 
   reg __412884_412884;
   reg _412885_412885 ; 
   reg __412885_412885;
   reg _412886_412886 ; 
   reg __412886_412886;
   reg _412887_412887 ; 
   reg __412887_412887;
   reg _412888_412888 ; 
   reg __412888_412888;
   reg _412889_412889 ; 
   reg __412889_412889;
   reg _412890_412890 ; 
   reg __412890_412890;
   reg _412891_412891 ; 
   reg __412891_412891;
   reg _412892_412892 ; 
   reg __412892_412892;
   reg _412893_412893 ; 
   reg __412893_412893;
   reg _412894_412894 ; 
   reg __412894_412894;
   reg _412895_412895 ; 
   reg __412895_412895;
   reg _412896_412896 ; 
   reg __412896_412896;
   reg _412897_412897 ; 
   reg __412897_412897;
   reg _412898_412898 ; 
   reg __412898_412898;
   reg _412899_412899 ; 
   reg __412899_412899;
   reg _412900_412900 ; 
   reg __412900_412900;
   reg _412901_412901 ; 
   reg __412901_412901;
   reg _412902_412902 ; 
   reg __412902_412902;
   reg _412903_412903 ; 
   reg __412903_412903;
   reg _412904_412904 ; 
   reg __412904_412904;
   reg _412905_412905 ; 
   reg __412905_412905;
   reg _412906_412906 ; 
   reg __412906_412906;
   reg _412907_412907 ; 
   reg __412907_412907;
   reg _412908_412908 ; 
   reg __412908_412908;
   reg _412909_412909 ; 
   reg __412909_412909;
   reg _412910_412910 ; 
   reg __412910_412910;
   reg _412911_412911 ; 
   reg __412911_412911;
   reg _412912_412912 ; 
   reg __412912_412912;
   reg _412913_412913 ; 
   reg __412913_412913;
   reg _412914_412914 ; 
   reg __412914_412914;
   reg _412915_412915 ; 
   reg __412915_412915;
   reg _412916_412916 ; 
   reg __412916_412916;
   reg _412917_412917 ; 
   reg __412917_412917;
   reg _412918_412918 ; 
   reg __412918_412918;
   reg _412919_412919 ; 
   reg __412919_412919;
   reg _412920_412920 ; 
   reg __412920_412920;
   reg _412921_412921 ; 
   reg __412921_412921;
   reg _412922_412922 ; 
   reg __412922_412922;
   reg _412923_412923 ; 
   reg __412923_412923;
   reg _412924_412924 ; 
   reg __412924_412924;
   reg _412925_412925 ; 
   reg __412925_412925;
   reg _412926_412926 ; 
   reg __412926_412926;
   reg _412927_412927 ; 
   reg __412927_412927;
   reg _412928_412928 ; 
   reg __412928_412928;
   reg _412929_412929 ; 
   reg __412929_412929;
   reg _412930_412930 ; 
   reg __412930_412930;
   reg _412931_412931 ; 
   reg __412931_412931;
   reg _412932_412932 ; 
   reg __412932_412932;
   reg _412933_412933 ; 
   reg __412933_412933;
   reg _412934_412934 ; 
   reg __412934_412934;
   reg _412935_412935 ; 
   reg __412935_412935;
   reg _412936_412936 ; 
   reg __412936_412936;
   reg _412937_412937 ; 
   reg __412937_412937;
   reg _412938_412938 ; 
   reg __412938_412938;
   reg _412939_412939 ; 
   reg __412939_412939;
   reg _412940_412940 ; 
   reg __412940_412940;
   reg _412941_412941 ; 
   reg __412941_412941;
   reg _412942_412942 ; 
   reg __412942_412942;
   reg _412943_412943 ; 
   reg __412943_412943;
   reg _412944_412944 ; 
   reg __412944_412944;
   reg _412945_412945 ; 
   reg __412945_412945;
   reg _412946_412946 ; 
   reg __412946_412946;
   reg _412947_412947 ; 
   reg __412947_412947;
   reg _412948_412948 ; 
   reg __412948_412948;
   reg _412949_412949 ; 
   reg __412949_412949;
   reg _412950_412950 ; 
   reg __412950_412950;
   reg _412951_412951 ; 
   reg __412951_412951;
   reg _412952_412952 ; 
   reg __412952_412952;
   reg _412953_412953 ; 
   reg __412953_412953;
   reg _412954_412954 ; 
   reg __412954_412954;
   reg _412955_412955 ; 
   reg __412955_412955;
   reg _412956_412956 ; 
   reg __412956_412956;
   reg _412957_412957 ; 
   reg __412957_412957;
   reg _412958_412958 ; 
   reg __412958_412958;
   reg _412959_412959 ; 
   reg __412959_412959;
   reg _412960_412960 ; 
   reg __412960_412960;
   reg _412961_412961 ; 
   reg __412961_412961;
   reg _412962_412962 ; 
   reg __412962_412962;
   reg _412963_412963 ; 
   reg __412963_412963;
   reg _412964_412964 ; 
   reg __412964_412964;
   reg _412965_412965 ; 
   reg __412965_412965;
   reg _412966_412966 ; 
   reg __412966_412966;
   reg _412967_412967 ; 
   reg __412967_412967;
   reg _412968_412968 ; 
   reg __412968_412968;
   reg _412969_412969 ; 
   reg __412969_412969;
   reg _412970_412970 ; 
   reg __412970_412970;
   reg _412971_412971 ; 
   reg __412971_412971;
   reg _412972_412972 ; 
   reg __412972_412972;
   reg _412973_412973 ; 
   reg __412973_412973;
   reg _412974_412974 ; 
   reg __412974_412974;
   reg _412975_412975 ; 
   reg __412975_412975;
   reg _412976_412976 ; 
   reg __412976_412976;
   reg _412977_412977 ; 
   reg __412977_412977;
   reg _412978_412978 ; 
   reg __412978_412978;
   reg _412979_412979 ; 
   reg __412979_412979;
   reg _412980_412980 ; 
   reg __412980_412980;
   reg _412981_412981 ; 
   reg __412981_412981;
   reg _412982_412982 ; 
   reg __412982_412982;
   reg _412983_412983 ; 
   reg __412983_412983;
   reg _412984_412984 ; 
   reg __412984_412984;
   reg _412985_412985 ; 
   reg __412985_412985;
   reg _412986_412986 ; 
   reg __412986_412986;
   reg _412987_412987 ; 
   reg __412987_412987;
   reg _412988_412988 ; 
   reg __412988_412988;
   reg _412989_412989 ; 
   reg __412989_412989;
   reg _412990_412990 ; 
   reg __412990_412990;
   reg _412991_412991 ; 
   reg __412991_412991;
   reg _412992_412992 ; 
   reg __412992_412992;
   reg _412993_412993 ; 
   reg __412993_412993;
   reg _412994_412994 ; 
   reg __412994_412994;
   reg _412995_412995 ; 
   reg __412995_412995;
   reg _412996_412996 ; 
   reg __412996_412996;
   reg _412997_412997 ; 
   reg __412997_412997;
   reg _412998_412998 ; 
   reg __412998_412998;
   reg _412999_412999 ; 
   reg __412999_412999;
   reg _413000_413000 ; 
   reg __413000_413000;
   reg _413001_413001 ; 
   reg __413001_413001;
   reg _413002_413002 ; 
   reg __413002_413002;
   reg _413003_413003 ; 
   reg __413003_413003;
   reg _413004_413004 ; 
   reg __413004_413004;
   reg _413005_413005 ; 
   reg __413005_413005;
   reg _413006_413006 ; 
   reg __413006_413006;
   reg _413007_413007 ; 
   reg __413007_413007;
   reg _413008_413008 ; 
   reg __413008_413008;
   reg _413009_413009 ; 
   reg __413009_413009;
   reg _413010_413010 ; 
   reg __413010_413010;
   reg _413011_413011 ; 
   reg __413011_413011;
   reg _413012_413012 ; 
   reg __413012_413012;
   reg _413013_413013 ; 
   reg __413013_413013;
   reg _413014_413014 ; 
   reg __413014_413014;
   reg _413015_413015 ; 
   reg __413015_413015;
   reg _413016_413016 ; 
   reg __413016_413016;
   reg _413017_413017 ; 
   reg __413017_413017;
   reg _413018_413018 ; 
   reg __413018_413018;
   reg _413019_413019 ; 
   reg __413019_413019;
   reg _413020_413020 ; 
   reg __413020_413020;
   reg _413021_413021 ; 
   reg __413021_413021;
   reg _413022_413022 ; 
   reg __413022_413022;
   reg _413023_413023 ; 
   reg __413023_413023;
   reg _413024_413024 ; 
   reg __413024_413024;
   reg _413025_413025 ; 
   reg __413025_413025;
   reg _413026_413026 ; 
   reg __413026_413026;
   reg _413027_413027 ; 
   reg __413027_413027;
   reg _413028_413028 ; 
   reg __413028_413028;
   reg _413029_413029 ; 
   reg __413029_413029;
   reg _413030_413030 ; 
   reg __413030_413030;
   reg _413031_413031 ; 
   reg __413031_413031;
   reg _413032_413032 ; 
   reg __413032_413032;
   reg _413033_413033 ; 
   reg __413033_413033;
   reg _413034_413034 ; 
   reg __413034_413034;
   reg _413035_413035 ; 
   reg __413035_413035;
   reg _413036_413036 ; 
   reg __413036_413036;
   reg _413037_413037 ; 
   reg __413037_413037;
   reg _413038_413038 ; 
   reg __413038_413038;
   reg _413039_413039 ; 
   reg __413039_413039;
   reg _413040_413040 ; 
   reg __413040_413040;
   reg _413041_413041 ; 
   reg __413041_413041;
   reg _413042_413042 ; 
   reg __413042_413042;
   reg _413043_413043 ; 
   reg __413043_413043;
   reg _413044_413044 ; 
   reg __413044_413044;
   reg _413045_413045 ; 
   reg __413045_413045;
   reg _413046_413046 ; 
   reg __413046_413046;
   reg _413047_413047 ; 
   reg __413047_413047;
   reg _413048_413048 ; 
   reg __413048_413048;
   reg _413049_413049 ; 
   reg __413049_413049;
   reg _413050_413050 ; 
   reg __413050_413050;
   reg _413051_413051 ; 
   reg __413051_413051;
   reg _413052_413052 ; 
   reg __413052_413052;
   reg _413053_413053 ; 
   reg __413053_413053;
   reg _413054_413054 ; 
   reg __413054_413054;
   reg _413055_413055 ; 
   reg __413055_413055;
   reg _413056_413056 ; 
   reg __413056_413056;
   reg _413057_413057 ; 
   reg __413057_413057;
   reg _413058_413058 ; 
   reg __413058_413058;
   reg _413059_413059 ; 
   reg __413059_413059;
   reg _413060_413060 ; 
   reg __413060_413060;
   reg _413061_413061 ; 
   reg __413061_413061;
   reg _413062_413062 ; 
   reg __413062_413062;
   reg _413063_413063 ; 
   reg __413063_413063;
   reg _413064_413064 ; 
   reg __413064_413064;
   reg _413065_413065 ; 
   reg __413065_413065;
   reg _413066_413066 ; 
   reg __413066_413066;
   reg _413067_413067 ; 
   reg __413067_413067;
   reg _413068_413068 ; 
   reg __413068_413068;
   reg _413069_413069 ; 
   reg __413069_413069;
   reg _413070_413070 ; 
   reg __413070_413070;
   reg _413071_413071 ; 
   reg __413071_413071;
   reg _413072_413072 ; 
   reg __413072_413072;
   reg _413073_413073 ; 
   reg __413073_413073;
   reg _413074_413074 ; 
   reg __413074_413074;
   reg _413075_413075 ; 
   reg __413075_413075;
   reg _413076_413076 ; 
   reg __413076_413076;
   reg _413077_413077 ; 
   reg __413077_413077;
   reg _413078_413078 ; 
   reg __413078_413078;
   reg _413079_413079 ; 
   reg __413079_413079;
   reg _413080_413080 ; 
   reg __413080_413080;
   reg _413081_413081 ; 
   reg __413081_413081;
   reg _413082_413082 ; 
   reg __413082_413082;
   reg _413083_413083 ; 
   reg __413083_413083;
   reg _413084_413084 ; 
   reg __413084_413084;
   reg _413085_413085 ; 
   reg __413085_413085;
   reg _413086_413086 ; 
   reg __413086_413086;
   reg _413087_413087 ; 
   reg __413087_413087;
   reg _413088_413088 ; 
   reg __413088_413088;
   reg _413089_413089 ; 
   reg __413089_413089;
   reg _413090_413090 ; 
   reg __413090_413090;
   reg _413091_413091 ; 
   reg __413091_413091;
   reg _413092_413092 ; 
   reg __413092_413092;
   reg _413093_413093 ; 
   reg __413093_413093;
   reg _413094_413094 ; 
   reg __413094_413094;
   reg _413095_413095 ; 
   reg __413095_413095;
   reg _413096_413096 ; 
   reg __413096_413096;
   reg _413097_413097 ; 
   reg __413097_413097;
   reg _413098_413098 ; 
   reg __413098_413098;
   reg _413099_413099 ; 
   reg __413099_413099;
   reg _413100_413100 ; 
   reg __413100_413100;
   reg _413101_413101 ; 
   reg __413101_413101;
   reg _413102_413102 ; 
   reg __413102_413102;
   reg _413103_413103 ; 
   reg __413103_413103;
   reg _413104_413104 ; 
   reg __413104_413104;
   reg _413105_413105 ; 
   reg __413105_413105;
   reg _413106_413106 ; 
   reg __413106_413106;
   reg _413107_413107 ; 
   reg __413107_413107;
   reg _413108_413108 ; 
   reg __413108_413108;
   reg _413109_413109 ; 
   reg __413109_413109;
   reg _413110_413110 ; 
   reg __413110_413110;
   reg _413111_413111 ; 
   reg __413111_413111;
   reg _413112_413112 ; 
   reg __413112_413112;
   reg _413113_413113 ; 
   reg __413113_413113;
   reg _413114_413114 ; 
   reg __413114_413114;
   reg _413115_413115 ; 
   reg __413115_413115;
   reg _413116_413116 ; 
   reg __413116_413116;
   reg _413117_413117 ; 
   reg __413117_413117;
   reg _413118_413118 ; 
   reg __413118_413118;
   reg _413119_413119 ; 
   reg __413119_413119;
   reg _413120_413120 ; 
   reg __413120_413120;
   reg _413121_413121 ; 
   reg __413121_413121;
   reg _413122_413122 ; 
   reg __413122_413122;
   reg _413123_413123 ; 
   reg __413123_413123;
   reg _413124_413124 ; 
   reg __413124_413124;
   reg _413125_413125 ; 
   reg __413125_413125;
   reg _413126_413126 ; 
   reg __413126_413126;
   reg _413127_413127 ; 
   reg __413127_413127;
   reg _413128_413128 ; 
   reg __413128_413128;
   reg _413129_413129 ; 
   reg __413129_413129;
   reg _413130_413130 ; 
   reg __413130_413130;
   reg _413131_413131 ; 
   reg __413131_413131;
   reg _413132_413132 ; 
   reg __413132_413132;
   reg _413133_413133 ; 
   reg __413133_413133;
   reg _413134_413134 ; 
   reg __413134_413134;
   reg _413135_413135 ; 
   reg __413135_413135;
   reg _413136_413136 ; 
   reg __413136_413136;
   reg _413137_413137 ; 
   reg __413137_413137;
   reg _413138_413138 ; 
   reg __413138_413138;
   reg _413139_413139 ; 
   reg __413139_413139;
   reg _413140_413140 ; 
   reg __413140_413140;
   reg _413141_413141 ; 
   reg __413141_413141;
   reg _413142_413142 ; 
   reg __413142_413142;
   reg _413143_413143 ; 
   reg __413143_413143;
   reg _413144_413144 ; 
   reg __413144_413144;
   reg _413145_413145 ; 
   reg __413145_413145;
   reg _413146_413146 ; 
   reg __413146_413146;
   reg _413147_413147 ; 
   reg __413147_413147;
   reg _413148_413148 ; 
   reg __413148_413148;
   reg _413149_413149 ; 
   reg __413149_413149;
   reg _413150_413150 ; 
   reg __413150_413150;
   reg _413151_413151 ; 
   reg __413151_413151;
   reg _413152_413152 ; 
   reg __413152_413152;
   reg _413153_413153 ; 
   reg __413153_413153;
   reg _413154_413154 ; 
   reg __413154_413154;
   reg _413155_413155 ; 
   reg __413155_413155;
   reg _413156_413156 ; 
   reg __413156_413156;
   reg _413157_413157 ; 
   reg __413157_413157;
   reg _413158_413158 ; 
   reg __413158_413158;
   reg _413159_413159 ; 
   reg __413159_413159;
   reg _413160_413160 ; 
   reg __413160_413160;
   reg _413161_413161 ; 
   reg __413161_413161;
   reg _413162_413162 ; 
   reg __413162_413162;
   reg _413163_413163 ; 
   reg __413163_413163;
   reg _413164_413164 ; 
   reg __413164_413164;
   reg _413165_413165 ; 
   reg __413165_413165;
   reg _413166_413166 ; 
   reg __413166_413166;
   reg _413167_413167 ; 
   reg __413167_413167;
   reg _413168_413168 ; 
   reg __413168_413168;
   reg _413169_413169 ; 
   reg __413169_413169;
   reg _413170_413170 ; 
   reg __413170_413170;
   reg _413171_413171 ; 
   reg __413171_413171;
   reg _413172_413172 ; 
   reg __413172_413172;
   reg _413173_413173 ; 
   reg __413173_413173;
   reg _413174_413174 ; 
   reg __413174_413174;
   reg _413175_413175 ; 
   reg __413175_413175;
   reg _413176_413176 ; 
   reg __413176_413176;
   reg _413177_413177 ; 
   reg __413177_413177;
   reg _413178_413178 ; 
   reg __413178_413178;
   reg _413179_413179 ; 
   reg __413179_413179;
   reg _413180_413180 ; 
   reg __413180_413180;
   reg _413181_413181 ; 
   reg __413181_413181;
   reg _413182_413182 ; 
   reg __413182_413182;
   reg _413183_413183 ; 
   reg __413183_413183;
   reg _413184_413184 ; 
   reg __413184_413184;
   reg _413185_413185 ; 
   reg __413185_413185;
   reg _413186_413186 ; 
   reg __413186_413186;
   reg _413187_413187 ; 
   reg __413187_413187;
   reg _413188_413188 ; 
   reg __413188_413188;
   reg _413189_413189 ; 
   reg __413189_413189;
   reg _413190_413190 ; 
   reg __413190_413190;
   reg _413191_413191 ; 
   reg __413191_413191;
   reg _413192_413192 ; 
   reg __413192_413192;
   reg _413193_413193 ; 
   reg __413193_413193;
   reg _413194_413194 ; 
   reg __413194_413194;
   reg _413195_413195 ; 
   reg __413195_413195;
   reg _413196_413196 ; 
   reg __413196_413196;
   reg _413197_413197 ; 
   reg __413197_413197;
   reg _413198_413198 ; 
   reg __413198_413198;
   reg _413199_413199 ; 
   reg __413199_413199;
   reg _413200_413200 ; 
   reg __413200_413200;
   reg _413201_413201 ; 
   reg __413201_413201;
   reg _413202_413202 ; 
   reg __413202_413202;
   reg _413203_413203 ; 
   reg __413203_413203;
   reg _413204_413204 ; 
   reg __413204_413204;
   reg _413205_413205 ; 
   reg __413205_413205;
   reg _413206_413206 ; 
   reg __413206_413206;
   reg _413207_413207 ; 
   reg __413207_413207;
   reg _413208_413208 ; 
   reg __413208_413208;
   reg _413209_413209 ; 
   reg __413209_413209;
   reg _413210_413210 ; 
   reg __413210_413210;
   reg _413211_413211 ; 
   reg __413211_413211;
   reg _413212_413212 ; 
   reg __413212_413212;
   reg _413213_413213 ; 
   reg __413213_413213;
   reg _413214_413214 ; 
   reg __413214_413214;
   reg _413215_413215 ; 
   reg __413215_413215;
   reg _413216_413216 ; 
   reg __413216_413216;
   reg _413217_413217 ; 
   reg __413217_413217;
   reg _413218_413218 ; 
   reg __413218_413218;
   reg _413219_413219 ; 
   reg __413219_413219;
   reg _413220_413220 ; 
   reg __413220_413220;
   reg _413221_413221 ; 
   reg __413221_413221;
   reg _413222_413222 ; 
   reg __413222_413222;
   reg _413223_413223 ; 
   reg __413223_413223;
   reg _413224_413224 ; 
   reg __413224_413224;
   reg _413225_413225 ; 
   reg __413225_413225;
   reg _413226_413226 ; 
   reg __413226_413226;
   reg _413227_413227 ; 
   reg __413227_413227;
   reg _413228_413228 ; 
   reg __413228_413228;
   reg _413229_413229 ; 
   reg __413229_413229;
   reg _413230_413230 ; 
   reg __413230_413230;
   reg _413231_413231 ; 
   reg __413231_413231;
   reg _413232_413232 ; 
   reg __413232_413232;
   reg _413233_413233 ; 
   reg __413233_413233;
   reg _413234_413234 ; 
   reg __413234_413234;
   reg _413235_413235 ; 
   reg __413235_413235;
   reg _413236_413236 ; 
   reg __413236_413236;
   reg _413237_413237 ; 
   reg __413237_413237;
   reg _413238_413238 ; 
   reg __413238_413238;
   reg _413239_413239 ; 
   reg __413239_413239;
   reg _413240_413240 ; 
   reg __413240_413240;
   reg _413241_413241 ; 
   reg __413241_413241;
   reg _413242_413242 ; 
   reg __413242_413242;
   reg _413243_413243 ; 
   reg __413243_413243;
   reg _413244_413244 ; 
   reg __413244_413244;
   reg _413245_413245 ; 
   reg __413245_413245;
   reg _413246_413246 ; 
   reg __413246_413246;
   reg _413247_413247 ; 
   reg __413247_413247;
   reg _413248_413248 ; 
   reg __413248_413248;
   reg _413249_413249 ; 
   reg __413249_413249;
   reg _413250_413250 ; 
   reg __413250_413250;
   reg _413251_413251 ; 
   reg __413251_413251;
   reg _413252_413252 ; 
   reg __413252_413252;
   reg _413253_413253 ; 
   reg __413253_413253;
   reg _413254_413254 ; 
   reg __413254_413254;
   reg _413255_413255 ; 
   reg __413255_413255;
   reg _413256_413256 ; 
   reg __413256_413256;
   reg _413257_413257 ; 
   reg __413257_413257;
   reg _413258_413258 ; 
   reg __413258_413258;
   reg _413259_413259 ; 
   reg __413259_413259;
   reg _413260_413260 ; 
   reg __413260_413260;
   reg _413261_413261 ; 
   reg __413261_413261;
   reg _413262_413262 ; 
   reg __413262_413262;
   reg _413263_413263 ; 
   reg __413263_413263;
   reg _413264_413264 ; 
   reg __413264_413264;
   reg _413265_413265 ; 
   reg __413265_413265;
   reg _413266_413266 ; 
   reg __413266_413266;
   reg _413267_413267 ; 
   reg __413267_413267;
   reg _413268_413268 ; 
   reg __413268_413268;
   reg _413269_413269 ; 
   reg __413269_413269;
   reg _413270_413270 ; 
   reg __413270_413270;
   reg _413271_413271 ; 
   reg __413271_413271;
   reg _413272_413272 ; 
   reg __413272_413272;
   reg _413273_413273 ; 
   reg __413273_413273;
   reg _413274_413274 ; 
   reg __413274_413274;
   reg _413275_413275 ; 
   reg __413275_413275;
   reg _413276_413276 ; 
   reg __413276_413276;
   reg _413277_413277 ; 
   reg __413277_413277;
   reg _413278_413278 ; 
   reg __413278_413278;
   reg _413279_413279 ; 
   reg __413279_413279;
   reg _413280_413280 ; 
   reg __413280_413280;
   reg _413281_413281 ; 
   reg __413281_413281;
   reg _413282_413282 ; 
   reg __413282_413282;
   reg _413283_413283 ; 
   reg __413283_413283;
   reg _413284_413284 ; 
   reg __413284_413284;
   reg _413285_413285 ; 
   reg __413285_413285;
   reg _413286_413286 ; 
   reg __413286_413286;
   reg _413287_413287 ; 
   reg __413287_413287;
   reg _413288_413288 ; 
   reg __413288_413288;
   reg _413289_413289 ; 
   reg __413289_413289;
   reg _413290_413290 ; 
   reg __413290_413290;
   reg _413291_413291 ; 
   reg __413291_413291;
   reg _413292_413292 ; 
   reg __413292_413292;
   reg _413293_413293 ; 
   reg __413293_413293;
   reg _413294_413294 ; 
   reg __413294_413294;
   reg _413295_413295 ; 
   reg __413295_413295;
   reg _413296_413296 ; 
   reg __413296_413296;
   reg _413297_413297 ; 
   reg __413297_413297;
   reg _413298_413298 ; 
   reg __413298_413298;
   reg _413299_413299 ; 
   reg __413299_413299;
   reg _413300_413300 ; 
   reg __413300_413300;
   reg _413301_413301 ; 
   reg __413301_413301;
   reg _413302_413302 ; 
   reg __413302_413302;
   reg _413303_413303 ; 
   reg __413303_413303;
   reg _413304_413304 ; 
   reg __413304_413304;
   reg _413305_413305 ; 
   reg __413305_413305;
   reg _413306_413306 ; 
   reg __413306_413306;
   reg _413307_413307 ; 
   reg __413307_413307;
   reg _413308_413308 ; 
   reg __413308_413308;
   reg _413309_413309 ; 
   reg __413309_413309;
   reg _413310_413310 ; 
   reg __413310_413310;
   reg _413311_413311 ; 
   reg __413311_413311;
   reg _413312_413312 ; 
   reg __413312_413312;
   reg _413313_413313 ; 
   reg __413313_413313;
   reg _413314_413314 ; 
   reg __413314_413314;
   reg _413315_413315 ; 
   reg __413315_413315;
   reg _413316_413316 ; 
   reg __413316_413316;
   reg _413317_413317 ; 
   reg __413317_413317;
   reg _413318_413318 ; 
   reg __413318_413318;
   reg _413319_413319 ; 
   reg __413319_413319;
   reg _413320_413320 ; 
   reg __413320_413320;
   reg _413321_413321 ; 
   reg __413321_413321;
   reg _413322_413322 ; 
   reg __413322_413322;
   reg _413323_413323 ; 
   reg __413323_413323;
   reg _413324_413324 ; 
   reg __413324_413324;
   reg _413325_413325 ; 
   reg __413325_413325;
   reg _413326_413326 ; 
   reg __413326_413326;
   reg _413327_413327 ; 
   reg __413327_413327;
   reg _413328_413328 ; 
   reg __413328_413328;
   reg _413329_413329 ; 
   reg __413329_413329;
   reg _413330_413330 ; 
   reg __413330_413330;
   reg _413331_413331 ; 
   reg __413331_413331;
   reg _413332_413332 ; 
   reg __413332_413332;
   reg _413333_413333 ; 
   reg __413333_413333;
   reg _413334_413334 ; 
   reg __413334_413334;
   reg _413335_413335 ; 
   reg __413335_413335;
   reg _413336_413336 ; 
   reg __413336_413336;
   reg _413337_413337 ; 
   reg __413337_413337;
   reg _413338_413338 ; 
   reg __413338_413338;
   reg _413339_413339 ; 
   reg __413339_413339;
   reg _413340_413340 ; 
   reg __413340_413340;
   reg _413341_413341 ; 
   reg __413341_413341;
   reg _413342_413342 ; 
   reg __413342_413342;
   reg _413343_413343 ; 
   reg __413343_413343;
   reg _413344_413344 ; 
   reg __413344_413344;
   reg _413345_413345 ; 
   reg __413345_413345;
   reg _413346_413346 ; 
   reg __413346_413346;
   reg _413347_413347 ; 
   reg __413347_413347;
   reg _413348_413348 ; 
   reg __413348_413348;
   reg _413349_413349 ; 
   reg __413349_413349;
   reg _413350_413350 ; 
   reg __413350_413350;
   reg _413351_413351 ; 
   reg __413351_413351;
   reg _413352_413352 ; 
   reg __413352_413352;
   reg _413353_413353 ; 
   reg __413353_413353;
   reg _413354_413354 ; 
   reg __413354_413354;
   reg _413355_413355 ; 
   reg __413355_413355;
   reg _413356_413356 ; 
   reg __413356_413356;
   reg _413357_413357 ; 
   reg __413357_413357;
   reg _413358_413358 ; 
   reg __413358_413358;
   reg _413359_413359 ; 
   reg __413359_413359;
   reg _413360_413360 ; 
   reg __413360_413360;
   reg _413361_413361 ; 
   reg __413361_413361;
   reg _413362_413362 ; 
   reg __413362_413362;
   reg _413363_413363 ; 
   reg __413363_413363;
   reg _413364_413364 ; 
   reg __413364_413364;
   reg _413365_413365 ; 
   reg __413365_413365;
   reg _413366_413366 ; 
   reg __413366_413366;
   reg _413367_413367 ; 
   reg __413367_413367;
   reg _413368_413368 ; 
   reg __413368_413368;
   reg _413369_413369 ; 
   reg __413369_413369;
   reg _413370_413370 ; 
   reg __413370_413370;
   reg _413371_413371 ; 
   reg __413371_413371;
   reg _413372_413372 ; 
   reg __413372_413372;
   reg _413373_413373 ; 
   reg __413373_413373;
   reg _413374_413374 ; 
   reg __413374_413374;
   reg _413375_413375 ; 
   reg __413375_413375;
   reg _413376_413376 ; 
   reg __413376_413376;
   reg _413377_413377 ; 
   reg __413377_413377;
   reg _413378_413378 ; 
   reg __413378_413378;
   reg _413379_413379 ; 
   reg __413379_413379;
   reg _413380_413380 ; 
   reg __413380_413380;
   reg _413381_413381 ; 
   reg __413381_413381;
   reg _413382_413382 ; 
   reg __413382_413382;
   reg _413383_413383 ; 
   reg __413383_413383;
   reg _413384_413384 ; 
   reg __413384_413384;
   reg _413385_413385 ; 
   reg __413385_413385;
   reg _413386_413386 ; 
   reg __413386_413386;
   reg _413387_413387 ; 
   reg __413387_413387;
   reg _413388_413388 ; 
   reg __413388_413388;
   reg _413389_413389 ; 
   reg __413389_413389;
   reg _413390_413390 ; 
   reg __413390_413390;
   reg _413391_413391 ; 
   reg __413391_413391;
   reg _413392_413392 ; 
   reg __413392_413392;
   reg _413393_413393 ; 
   reg __413393_413393;
   reg _413394_413394 ; 
   reg __413394_413394;
   reg _413395_413395 ; 
   reg __413395_413395;
   reg _413396_413396 ; 
   reg __413396_413396;
   reg _413397_413397 ; 
   reg __413397_413397;
   reg _413398_413398 ; 
   reg __413398_413398;
   reg _413399_413399 ; 
   reg __413399_413399;
   reg _413400_413400 ; 
   reg __413400_413400;
   reg _413401_413401 ; 
   reg __413401_413401;
   reg _413402_413402 ; 
   reg __413402_413402;
   reg _413403_413403 ; 
   reg __413403_413403;
   reg _413404_413404 ; 
   reg __413404_413404;
   reg _413405_413405 ; 
   reg __413405_413405;
   reg _413406_413406 ; 
   reg __413406_413406;
   reg _413407_413407 ; 
   reg __413407_413407;
   reg _413408_413408 ; 
   reg __413408_413408;
   reg _413409_413409 ; 
   reg __413409_413409;
   reg _413410_413410 ; 
   reg __413410_413410;
   reg _413411_413411 ; 
   reg __413411_413411;
   reg _413412_413412 ; 
   reg __413412_413412;
   reg _413413_413413 ; 
   reg __413413_413413;
   reg _413414_413414 ; 
   reg __413414_413414;
   reg _413415_413415 ; 
   reg __413415_413415;
   reg _413416_413416 ; 
   reg __413416_413416;
   reg _413417_413417 ; 
   reg __413417_413417;
   reg _413418_413418 ; 
   reg __413418_413418;
   reg _413419_413419 ; 
   reg __413419_413419;
   reg _413420_413420 ; 
   reg __413420_413420;
   reg _413421_413421 ; 
   reg __413421_413421;
   reg _413422_413422 ; 
   reg __413422_413422;
   reg _413423_413423 ; 
   reg __413423_413423;
   reg _413424_413424 ; 
   reg __413424_413424;
   reg _413425_413425 ; 
   reg __413425_413425;
   reg _413426_413426 ; 
   reg __413426_413426;
   reg _413427_413427 ; 
   reg __413427_413427;
   reg _413428_413428 ; 
   reg __413428_413428;
   reg _413429_413429 ; 
   reg __413429_413429;
   reg _413430_413430 ; 
   reg __413430_413430;
   reg _413431_413431 ; 
   reg __413431_413431;
   reg _413432_413432 ; 
   reg __413432_413432;
   reg _413433_413433 ; 
   reg __413433_413433;
   reg _413434_413434 ; 
   reg __413434_413434;
   reg _413435_413435 ; 
   reg __413435_413435;
   reg _413436_413436 ; 
   reg __413436_413436;
   reg _413437_413437 ; 
   reg __413437_413437;
   reg _413438_413438 ; 
   reg __413438_413438;
   reg _413439_413439 ; 
   reg __413439_413439;
   reg _413440_413440 ; 
   reg __413440_413440;
   reg _413441_413441 ; 
   reg __413441_413441;
   reg _413442_413442 ; 
   reg __413442_413442;
   reg _413443_413443 ; 
   reg __413443_413443;
   reg _413444_413444 ; 
   reg __413444_413444;
   reg _413445_413445 ; 
   reg __413445_413445;
   reg _413446_413446 ; 
   reg __413446_413446;
   reg _413447_413447 ; 
   reg __413447_413447;
   reg _413448_413448 ; 
   reg __413448_413448;
   reg _413449_413449 ; 
   reg __413449_413449;
   reg _413450_413450 ; 
   reg __413450_413450;
   reg _413451_413451 ; 
   reg __413451_413451;
   reg _413452_413452 ; 
   reg __413452_413452;
   reg _413453_413453 ; 
   reg __413453_413453;
   reg _413454_413454 ; 
   reg __413454_413454;
   reg _413455_413455 ; 
   reg __413455_413455;
   reg _413456_413456 ; 
   reg __413456_413456;
   reg _413457_413457 ; 
   reg __413457_413457;
   reg _413458_413458 ; 
   reg __413458_413458;
   reg _413459_413459 ; 
   reg __413459_413459;
   reg _413460_413460 ; 
   reg __413460_413460;
   reg _413461_413461 ; 
   reg __413461_413461;
   reg _413462_413462 ; 
   reg __413462_413462;
   reg _413463_413463 ; 
   reg __413463_413463;
   reg _413464_413464 ; 
   reg __413464_413464;
   reg _413465_413465 ; 
   reg __413465_413465;
   reg _413466_413466 ; 
   reg __413466_413466;
   reg _413467_413467 ; 
   reg __413467_413467;
   reg _413468_413468 ; 
   reg __413468_413468;
   reg _413469_413469 ; 
   reg __413469_413469;
   reg _413470_413470 ; 
   reg __413470_413470;
   reg _413471_413471 ; 
   reg __413471_413471;
   reg _413472_413472 ; 
   reg __413472_413472;
   reg _413473_413473 ; 
   reg __413473_413473;
   reg _413474_413474 ; 
   reg __413474_413474;
   reg _413475_413475 ; 
   reg __413475_413475;
   reg _413476_413476 ; 
   reg __413476_413476;
   reg _413477_413477 ; 
   reg __413477_413477;
   reg _413478_413478 ; 
   reg __413478_413478;
   reg _413479_413479 ; 
   reg __413479_413479;
   reg _413480_413480 ; 
   reg __413480_413480;
   reg _413481_413481 ; 
   reg __413481_413481;
   reg _413482_413482 ; 
   reg __413482_413482;
   reg _413483_413483 ; 
   reg __413483_413483;
   reg _413484_413484 ; 
   reg __413484_413484;
   reg _413485_413485 ; 
   reg __413485_413485;
   reg _413486_413486 ; 
   reg __413486_413486;
   reg _413487_413487 ; 
   reg __413487_413487;
   reg _413488_413488 ; 
   reg __413488_413488;
   reg _413489_413489 ; 
   reg __413489_413489;
   reg _413490_413490 ; 
   reg __413490_413490;
   reg _413491_413491 ; 
   reg __413491_413491;
   reg _413492_413492 ; 
   reg __413492_413492;
   reg _413493_413493 ; 
   reg __413493_413493;
   reg _413494_413494 ; 
   reg __413494_413494;
   reg _413495_413495 ; 
   reg __413495_413495;
   reg _413496_413496 ; 
   reg __413496_413496;
   reg _413497_413497 ; 
   reg __413497_413497;
   reg _413498_413498 ; 
   reg __413498_413498;
   reg _413499_413499 ; 
   reg __413499_413499;
   reg _413500_413500 ; 
   reg __413500_413500;
   reg _413501_413501 ; 
   reg __413501_413501;
   reg _413502_413502 ; 
   reg __413502_413502;
   reg _413503_413503 ; 
   reg __413503_413503;
   reg _413504_413504 ; 
   reg __413504_413504;
   reg _413505_413505 ; 
   reg __413505_413505;
   reg _413506_413506 ; 
   reg __413506_413506;
   reg _413507_413507 ; 
   reg __413507_413507;
   reg _413508_413508 ; 
   reg __413508_413508;
   reg _413509_413509 ; 
   reg __413509_413509;
   reg _413510_413510 ; 
   reg __413510_413510;
   reg _413511_413511 ; 
   reg __413511_413511;
   reg _413512_413512 ; 
   reg __413512_413512;
   reg _413513_413513 ; 
   reg __413513_413513;
   reg _413514_413514 ; 
   reg __413514_413514;
   reg _413515_413515 ; 
   reg __413515_413515;
   reg _413516_413516 ; 
   reg __413516_413516;
   reg _413517_413517 ; 
   reg __413517_413517;
   reg _413518_413518 ; 
   reg __413518_413518;
   reg _413519_413519 ; 
   reg __413519_413519;
   reg _413520_413520 ; 
   reg __413520_413520;
   reg _413521_413521 ; 
   reg __413521_413521;
   reg _413522_413522 ; 
   reg __413522_413522;
   reg _413523_413523 ; 
   reg __413523_413523;
   reg _413524_413524 ; 
   reg __413524_413524;
   reg _413525_413525 ; 
   reg __413525_413525;
   reg _413526_413526 ; 
   reg __413526_413526;
   reg _413527_413527 ; 
   reg __413527_413527;
   reg _413528_413528 ; 
   reg __413528_413528;
   reg _413529_413529 ; 
   reg __413529_413529;
   reg _413530_413530 ; 
   reg __413530_413530;
   reg _413531_413531 ; 
   reg __413531_413531;
   reg _413532_413532 ; 
   reg __413532_413532;
   reg _413533_413533 ; 
   reg __413533_413533;
   reg _413534_413534 ; 
   reg __413534_413534;
   reg _413535_413535 ; 
   reg __413535_413535;
   reg _413536_413536 ; 
   reg __413536_413536;
   reg _413537_413537 ; 
   reg __413537_413537;
   reg _413538_413538 ; 
   reg __413538_413538;
   reg _413539_413539 ; 
   reg __413539_413539;
   reg _413540_413540 ; 
   reg __413540_413540;
   reg _413541_413541 ; 
   reg __413541_413541;
   reg _413542_413542 ; 
   reg __413542_413542;
   reg _413543_413543 ; 
   reg __413543_413543;
   reg _413544_413544 ; 
   reg __413544_413544;
   reg _413545_413545 ; 
   reg __413545_413545;
   reg _413546_413546 ; 
   reg __413546_413546;
   reg _413547_413547 ; 
   reg __413547_413547;
   reg _413548_413548 ; 
   reg __413548_413548;
   reg _413549_413549 ; 
   reg __413549_413549;
   reg _413550_413550 ; 
   reg __413550_413550;
   reg _413551_413551 ; 
   reg __413551_413551;
   reg _413552_413552 ; 
   reg __413552_413552;
   reg _413553_413553 ; 
   reg __413553_413553;
   reg _413554_413554 ; 
   reg __413554_413554;
   reg _413555_413555 ; 
   reg __413555_413555;
   reg _413556_413556 ; 
   reg __413556_413556;
   reg _413557_413557 ; 
   reg __413557_413557;
   reg _413558_413558 ; 
   reg __413558_413558;
   reg _413559_413559 ; 
   reg __413559_413559;
   reg _413560_413560 ; 
   reg __413560_413560;
   reg _413561_413561 ; 
   reg __413561_413561;
   reg _413562_413562 ; 
   reg __413562_413562;
   reg _413563_413563 ; 
   reg __413563_413563;
   reg _413564_413564 ; 
   reg __413564_413564;
   reg _413565_413565 ; 
   reg __413565_413565;
   reg _413566_413566 ; 
   reg __413566_413566;
   reg _413567_413567 ; 
   reg __413567_413567;
   reg _413568_413568 ; 
   reg __413568_413568;
   reg _413569_413569 ; 
   reg __413569_413569;
   reg _413570_413570 ; 
   reg __413570_413570;
   reg _413571_413571 ; 
   reg __413571_413571;
   reg _413572_413572 ; 
   reg __413572_413572;
   reg _413573_413573 ; 
   reg __413573_413573;
   reg _413574_413574 ; 
   reg __413574_413574;
   reg _413575_413575 ; 
   reg __413575_413575;
   reg _413576_413576 ; 
   reg __413576_413576;
   reg _413577_413577 ; 
   reg __413577_413577;
   reg _413578_413578 ; 
   reg __413578_413578;
   reg _413579_413579 ; 
   reg __413579_413579;
   reg _413580_413580 ; 
   reg __413580_413580;
   reg _413581_413581 ; 
   reg __413581_413581;
   reg _413582_413582 ; 
   reg __413582_413582;
   reg _413583_413583 ; 
   reg __413583_413583;
   reg _413584_413584 ; 
   reg __413584_413584;
   reg _413585_413585 ; 
   reg __413585_413585;
   reg _413586_413586 ; 
   reg __413586_413586;
   reg _413587_413587 ; 
   reg __413587_413587;
   reg _413588_413588 ; 
   reg __413588_413588;
   reg _413589_413589 ; 
   reg __413589_413589;
   reg _413590_413590 ; 
   reg __413590_413590;
   reg _413591_413591 ; 
   reg __413591_413591;
   reg _413592_413592 ; 
   reg __413592_413592;
   reg _413593_413593 ; 
   reg __413593_413593;
   reg _413594_413594 ; 
   reg __413594_413594;
   reg _413595_413595 ; 
   reg __413595_413595;
   reg _413596_413596 ; 
   reg __413596_413596;
   reg _413597_413597 ; 
   reg __413597_413597;
   reg _413598_413598 ; 
   reg __413598_413598;
   reg _413599_413599 ; 
   reg __413599_413599;
   reg _413600_413600 ; 
   reg __413600_413600;
   reg _413601_413601 ; 
   reg __413601_413601;
   reg _413602_413602 ; 
   reg __413602_413602;
   reg _413603_413603 ; 
   reg __413603_413603;
   reg _413604_413604 ; 
   reg __413604_413604;
   reg _413605_413605 ; 
   reg __413605_413605;
   reg _413606_413606 ; 
   reg __413606_413606;
   reg _413607_413607 ; 
   reg __413607_413607;
   reg _413608_413608 ; 
   reg __413608_413608;
   reg _413609_413609 ; 
   reg __413609_413609;
   reg _413610_413610 ; 
   reg __413610_413610;
   reg _413611_413611 ; 
   reg __413611_413611;
   reg _413612_413612 ; 
   reg __413612_413612;
   reg _413613_413613 ; 
   reg __413613_413613;
   reg _413614_413614 ; 
   reg __413614_413614;
   reg _413615_413615 ; 
   reg __413615_413615;
   reg _413616_413616 ; 
   reg __413616_413616;
   reg _413617_413617 ; 
   reg __413617_413617;
   reg _413618_413618 ; 
   reg __413618_413618;
   reg _413619_413619 ; 
   reg __413619_413619;
   reg _413620_413620 ; 
   reg __413620_413620;
   reg _413621_413621 ; 
   reg __413621_413621;
   reg _413622_413622 ; 
   reg __413622_413622;
   reg _413623_413623 ; 
   reg __413623_413623;
   reg _413624_413624 ; 
   reg __413624_413624;
   reg _413625_413625 ; 
   reg __413625_413625;
   reg _413626_413626 ; 
   reg __413626_413626;
   reg _413627_413627 ; 
   reg __413627_413627;
   reg _413628_413628 ; 
   reg __413628_413628;
   reg _413629_413629 ; 
   reg __413629_413629;
   reg _413630_413630 ; 
   reg __413630_413630;
   reg _413631_413631 ; 
   reg __413631_413631;
   reg _413632_413632 ; 
   reg __413632_413632;
   reg _413633_413633 ; 
   reg __413633_413633;
   reg _413634_413634 ; 
   reg __413634_413634;
   reg _413635_413635 ; 
   reg __413635_413635;
   reg _413636_413636 ; 
   reg __413636_413636;
   reg _413637_413637 ; 
   reg __413637_413637;
   reg _413638_413638 ; 
   reg __413638_413638;
   reg _413639_413639 ; 
   reg __413639_413639;
   reg _413640_413640 ; 
   reg __413640_413640;
   reg _413641_413641 ; 
   reg __413641_413641;
   reg _413642_413642 ; 
   reg __413642_413642;
   reg _413643_413643 ; 
   reg __413643_413643;
   reg _413644_413644 ; 
   reg __413644_413644;
   reg _413645_413645 ; 
   reg __413645_413645;
   reg _413646_413646 ; 
   reg __413646_413646;
   reg _413647_413647 ; 
   reg __413647_413647;
   reg _413648_413648 ; 
   reg __413648_413648;
   reg _413649_413649 ; 
   reg __413649_413649;
   reg _413650_413650 ; 
   reg __413650_413650;
   reg _413651_413651 ; 
   reg __413651_413651;
   reg _413652_413652 ; 
   reg __413652_413652;
   reg _413653_413653 ; 
   reg __413653_413653;
   reg _413654_413654 ; 
   reg __413654_413654;
   reg _413655_413655 ; 
   reg __413655_413655;
   reg _413656_413656 ; 
   reg __413656_413656;
   reg _413657_413657 ; 
   reg __413657_413657;
   reg _413658_413658 ; 
   reg __413658_413658;
   reg _413659_413659 ; 
   reg __413659_413659;
   reg _413660_413660 ; 
   reg __413660_413660;
   reg _413661_413661 ; 
   reg __413661_413661;
   reg _413662_413662 ; 
   reg __413662_413662;
   reg _413663_413663 ; 
   reg __413663_413663;
   reg _413664_413664 ; 
   reg __413664_413664;
   reg _413665_413665 ; 
   reg __413665_413665;
   reg _413666_413666 ; 
   reg __413666_413666;
   reg _413667_413667 ; 
   reg __413667_413667;
   reg _413668_413668 ; 
   reg __413668_413668;
   reg _413669_413669 ; 
   reg __413669_413669;
   reg _413670_413670 ; 
   reg __413670_413670;
   reg _413671_413671 ; 
   reg __413671_413671;
   reg _413672_413672 ; 
   reg __413672_413672;
   reg _413673_413673 ; 
   reg __413673_413673;
   reg _413674_413674 ; 
   reg __413674_413674;
   reg _413675_413675 ; 
   reg __413675_413675;
   reg _413676_413676 ; 
   reg __413676_413676;
   reg _413677_413677 ; 
   reg __413677_413677;
   reg _413678_413678 ; 
   reg __413678_413678;
   reg _413679_413679 ; 
   reg __413679_413679;
   reg _413680_413680 ; 
   reg __413680_413680;
   reg _413681_413681 ; 
   reg __413681_413681;
   reg _413682_413682 ; 
   reg __413682_413682;
   reg _413683_413683 ; 
   reg __413683_413683;
   reg _413684_413684 ; 
   reg __413684_413684;
   reg _413685_413685 ; 
   reg __413685_413685;
   reg _413686_413686 ; 
   reg __413686_413686;
   reg _413687_413687 ; 
   reg __413687_413687;
   reg _413688_413688 ; 
   reg __413688_413688;
   reg _413689_413689 ; 
   reg __413689_413689;
   reg _413690_413690 ; 
   reg __413690_413690;
   reg _413691_413691 ; 
   reg __413691_413691;
   reg _413692_413692 ; 
   reg __413692_413692;
   reg _413693_413693 ; 
   reg __413693_413693;
   reg _413694_413694 ; 
   reg __413694_413694;
   reg _413695_413695 ; 
   reg __413695_413695;
   reg _413696_413696 ; 
   reg __413696_413696;
   reg _413697_413697 ; 
   reg __413697_413697;
   reg _413698_413698 ; 
   reg __413698_413698;
   reg _413699_413699 ; 
   reg __413699_413699;
   reg _413700_413700 ; 
   reg __413700_413700;
   reg _413701_413701 ; 
   reg __413701_413701;
   reg _413702_413702 ; 
   reg __413702_413702;
   reg _413703_413703 ; 
   reg __413703_413703;
   reg _413704_413704 ; 
   reg __413704_413704;
   reg _413705_413705 ; 
   reg __413705_413705;
   reg _413706_413706 ; 
   reg __413706_413706;
   reg _413707_413707 ; 
   reg __413707_413707;
   reg _413708_413708 ; 
   reg __413708_413708;
   reg _413709_413709 ; 
   reg __413709_413709;
   reg _413710_413710 ; 
   reg __413710_413710;
   reg _413711_413711 ; 
   reg __413711_413711;
   reg _413712_413712 ; 
   reg __413712_413712;
   reg _413713_413713 ; 
   reg __413713_413713;
   reg _413714_413714 ; 
   reg __413714_413714;
   reg _413715_413715 ; 
   reg __413715_413715;
   reg _413716_413716 ; 
   reg __413716_413716;
   reg _413717_413717 ; 
   reg __413717_413717;
   reg _413718_413718 ; 
   reg __413718_413718;
   reg _413719_413719 ; 
   reg __413719_413719;
   reg _413720_413720 ; 
   reg __413720_413720;
   reg _413721_413721 ; 
   reg __413721_413721;
   reg _413722_413722 ; 
   reg __413722_413722;
   reg _413723_413723 ; 
   reg __413723_413723;
   reg _413724_413724 ; 
   reg __413724_413724;
   reg _413725_413725 ; 
   reg __413725_413725;
   reg _413726_413726 ; 
   reg __413726_413726;
   reg _413727_413727 ; 
   reg __413727_413727;
   reg _413728_413728 ; 
   reg __413728_413728;
   reg _413729_413729 ; 
   reg __413729_413729;
   reg _413730_413730 ; 
   reg __413730_413730;
   reg _413731_413731 ; 
   reg __413731_413731;
   reg _413732_413732 ; 
   reg __413732_413732;
   reg _413733_413733 ; 
   reg __413733_413733;
   reg _413734_413734 ; 
   reg __413734_413734;
   reg _413735_413735 ; 
   reg __413735_413735;
   reg _413736_413736 ; 
   reg __413736_413736;
   reg _413737_413737 ; 
   reg __413737_413737;
   reg _413738_413738 ; 
   reg __413738_413738;
   reg _413739_413739 ; 
   reg __413739_413739;
   reg _413740_413740 ; 
   reg __413740_413740;
   reg _413741_413741 ; 
   reg __413741_413741;
   reg _413742_413742 ; 
   reg __413742_413742;
   reg _413743_413743 ; 
   reg __413743_413743;
   reg _413744_413744 ; 
   reg __413744_413744;
   reg _413745_413745 ; 
   reg __413745_413745;
   reg _413746_413746 ; 
   reg __413746_413746;
   reg _413747_413747 ; 
   reg __413747_413747;
   reg _413748_413748 ; 
   reg __413748_413748;
   reg _413749_413749 ; 
   reg __413749_413749;
   reg _413750_413750 ; 
   reg __413750_413750;
   reg _413751_413751 ; 
   reg __413751_413751;
   reg _413752_413752 ; 
   reg __413752_413752;
   reg _413753_413753 ; 
   reg __413753_413753;
   reg _413754_413754 ; 
   reg __413754_413754;
   reg _413755_413755 ; 
   reg __413755_413755;
   reg _413756_413756 ; 
   reg __413756_413756;
   reg _413757_413757 ; 
   reg __413757_413757;
   reg _413758_413758 ; 
   reg __413758_413758;
   reg _413759_413759 ; 
   reg __413759_413759;
   reg _413760_413760 ; 
   reg __413760_413760;
   reg _413761_413761 ; 
   reg __413761_413761;
   reg _413762_413762 ; 
   reg __413762_413762;
   reg _413763_413763 ; 
   reg __413763_413763;
   reg _413764_413764 ; 
   reg __413764_413764;
   reg _413765_413765 ; 
   reg __413765_413765;
   reg _413766_413766 ; 
   reg __413766_413766;
   reg _413767_413767 ; 
   reg __413767_413767;
   reg _413768_413768 ; 
   reg __413768_413768;
   reg _413769_413769 ; 
   reg __413769_413769;
   reg _413770_413770 ; 
   reg __413770_413770;
   reg _413771_413771 ; 
   reg __413771_413771;
   reg _413772_413772 ; 
   reg __413772_413772;
   reg _413773_413773 ; 
   reg __413773_413773;
   reg _413774_413774 ; 
   reg __413774_413774;
   reg _413775_413775 ; 
   reg __413775_413775;
   reg _413776_413776 ; 
   reg __413776_413776;
   reg _413777_413777 ; 
   reg __413777_413777;
   reg _413778_413778 ; 
   reg __413778_413778;
   reg _413779_413779 ; 
   reg __413779_413779;
   reg _413780_413780 ; 
   reg __413780_413780;
   reg _413781_413781 ; 
   reg __413781_413781;
   reg _413782_413782 ; 
   reg __413782_413782;
   reg _413783_413783 ; 
   reg __413783_413783;
   reg _413784_413784 ; 
   reg __413784_413784;
   reg _413785_413785 ; 
   reg __413785_413785;
   reg _413786_413786 ; 
   reg __413786_413786;
   reg _413787_413787 ; 
   reg __413787_413787;
   reg _413788_413788 ; 
   reg __413788_413788;
   reg _413789_413789 ; 
   reg __413789_413789;
   reg _413790_413790 ; 
   reg __413790_413790;
   reg _413791_413791 ; 
   reg __413791_413791;
   reg _413792_413792 ; 
   reg __413792_413792;
   reg _413793_413793 ; 
   reg __413793_413793;
   reg _413794_413794 ; 
   reg __413794_413794;
   reg _413795_413795 ; 
   reg __413795_413795;
   reg _413796_413796 ; 
   reg __413796_413796;
   reg _413797_413797 ; 
   reg __413797_413797;
   reg _413798_413798 ; 
   reg __413798_413798;
   reg _413799_413799 ; 
   reg __413799_413799;
   reg _413800_413800 ; 
   reg __413800_413800;
   reg _413801_413801 ; 
   reg __413801_413801;
   reg _413802_413802 ; 
   reg __413802_413802;
   reg _413803_413803 ; 
   reg __413803_413803;
   reg _413804_413804 ; 
   reg __413804_413804;
   reg _413805_413805 ; 
   reg __413805_413805;
   reg _413806_413806 ; 
   reg __413806_413806;
   reg _413807_413807 ; 
   reg __413807_413807;
   reg _413808_413808 ; 
   reg __413808_413808;
   reg _413809_413809 ; 
   reg __413809_413809;
   reg _413810_413810 ; 
   reg __413810_413810;
   reg _413811_413811 ; 
   reg __413811_413811;
   reg _413812_413812 ; 
   reg __413812_413812;
   reg _413813_413813 ; 
   reg __413813_413813;
   reg _413814_413814 ; 
   reg __413814_413814;
   reg _413815_413815 ; 
   reg __413815_413815;
   reg _413816_413816 ; 
   reg __413816_413816;
   reg _413817_413817 ; 
   reg __413817_413817;
   reg _413818_413818 ; 
   reg __413818_413818;
   reg _413819_413819 ; 
   reg __413819_413819;
   reg _413820_413820 ; 
   reg __413820_413820;
   reg _413821_413821 ; 
   reg __413821_413821;
   reg _413822_413822 ; 
   reg __413822_413822;
   reg _413823_413823 ; 
   reg __413823_413823;
   reg _413824_413824 ; 
   reg __413824_413824;
   reg _413825_413825 ; 
   reg __413825_413825;
   reg _413826_413826 ; 
   reg __413826_413826;
   reg _413827_413827 ; 
   reg __413827_413827;
   reg _413828_413828 ; 
   reg __413828_413828;
   reg _413829_413829 ; 
   reg __413829_413829;
   reg _413830_413830 ; 
   reg __413830_413830;
   reg _413831_413831 ; 
   reg __413831_413831;
   reg _413832_413832 ; 
   reg __413832_413832;
   reg _413833_413833 ; 
   reg __413833_413833;
   reg _413834_413834 ; 
   reg __413834_413834;
   reg _413835_413835 ; 
   reg __413835_413835;
   reg _413836_413836 ; 
   reg __413836_413836;
   reg _413837_413837 ; 
   reg __413837_413837;
   reg _413838_413838 ; 
   reg __413838_413838;
   reg _413839_413839 ; 
   reg __413839_413839;
   reg _413840_413840 ; 
   reg __413840_413840;
   reg _413841_413841 ; 
   reg __413841_413841;
   reg _413842_413842 ; 
   reg __413842_413842;
   reg _413843_413843 ; 
   reg __413843_413843;
   reg _413844_413844 ; 
   reg __413844_413844;
   reg _413845_413845 ; 
   reg __413845_413845;
   reg _413846_413846 ; 
   reg __413846_413846;
   reg _413847_413847 ; 
   reg __413847_413847;
   reg _413848_413848 ; 
   reg __413848_413848;
   reg _413849_413849 ; 
   reg __413849_413849;
   reg _413850_413850 ; 
   reg __413850_413850;
   reg _413851_413851 ; 
   reg __413851_413851;
   reg _413852_413852 ; 
   reg __413852_413852;
   reg _413853_413853 ; 
   reg __413853_413853;
   reg _413854_413854 ; 
   reg __413854_413854;
   reg _413855_413855 ; 
   reg __413855_413855;
   reg _413856_413856 ; 
   reg __413856_413856;
   reg _413857_413857 ; 
   reg __413857_413857;
   reg _413858_413858 ; 
   reg __413858_413858;
   reg _413859_413859 ; 
   reg __413859_413859;
   reg _413860_413860 ; 
   reg __413860_413860;
   reg _413861_413861 ; 
   reg __413861_413861;
   reg _413862_413862 ; 
   reg __413862_413862;
   reg _413863_413863 ; 
   reg __413863_413863;
   reg _413864_413864 ; 
   reg __413864_413864;
   reg _413865_413865 ; 
   reg __413865_413865;
   reg _413866_413866 ; 
   reg __413866_413866;
   reg _413867_413867 ; 
   reg __413867_413867;
   reg _413868_413868 ; 
   reg __413868_413868;
   reg _413869_413869 ; 
   reg __413869_413869;
   reg _413870_413870 ; 
   reg __413870_413870;
   reg _413871_413871 ; 
   reg __413871_413871;
   reg _413872_413872 ; 
   reg __413872_413872;
   reg _413873_413873 ; 
   reg __413873_413873;
   reg _413874_413874 ; 
   reg __413874_413874;
   reg _413875_413875 ; 
   reg __413875_413875;
   reg _413876_413876 ; 
   reg __413876_413876;
   reg _413877_413877 ; 
   reg __413877_413877;
   reg _413878_413878 ; 
   reg __413878_413878;
   reg _413879_413879 ; 
   reg __413879_413879;
   reg _413880_413880 ; 
   reg __413880_413880;
   reg _413881_413881 ; 
   reg __413881_413881;
   reg _413882_413882 ; 
   reg __413882_413882;
   reg _413883_413883 ; 
   reg __413883_413883;
   reg _413884_413884 ; 
   reg __413884_413884;
   reg _413885_413885 ; 
   reg __413885_413885;
   reg _413886_413886 ; 
   reg __413886_413886;
   reg _413887_413887 ; 
   reg __413887_413887;
   reg _413888_413888 ; 
   reg __413888_413888;
   reg _413889_413889 ; 
   reg __413889_413889;
   reg _413890_413890 ; 
   reg __413890_413890;
   reg _413891_413891 ; 
   reg __413891_413891;
   reg _413892_413892 ; 
   reg __413892_413892;
   reg _413893_413893 ; 
   reg __413893_413893;
   reg _413894_413894 ; 
   reg __413894_413894;
   reg _413895_413895 ; 
   reg __413895_413895;
   reg _413896_413896 ; 
   reg __413896_413896;
   reg _413897_413897 ; 
   reg __413897_413897;
   reg _413898_413898 ; 
   reg __413898_413898;
   reg _413899_413899 ; 
   reg __413899_413899;
   reg _413900_413900 ; 
   reg __413900_413900;
   reg _413901_413901 ; 
   reg __413901_413901;
   reg _413902_413902 ; 
   reg __413902_413902;
   reg _413903_413903 ; 
   reg __413903_413903;
   reg _413904_413904 ; 
   reg __413904_413904;
   reg _413905_413905 ; 
   reg __413905_413905;
   reg _413906_413906 ; 
   reg __413906_413906;
   reg _413907_413907 ; 
   reg __413907_413907;
   reg _413908_413908 ; 
   reg __413908_413908;
   reg _413909_413909 ; 
   reg __413909_413909;
   reg _413910_413910 ; 
   reg __413910_413910;
   reg _413911_413911 ; 
   reg __413911_413911;
   reg _413912_413912 ; 
   reg __413912_413912;
   reg _413913_413913 ; 
   reg __413913_413913;
   reg _413914_413914 ; 
   reg __413914_413914;
   reg _413915_413915 ; 
   reg __413915_413915;
   reg _413916_413916 ; 
   reg __413916_413916;
   reg _413917_413917 ; 
   reg __413917_413917;
   reg _413918_413918 ; 
   reg __413918_413918;
   reg _413919_413919 ; 
   reg __413919_413919;
   reg _413920_413920 ; 
   reg __413920_413920;
   reg _413921_413921 ; 
   reg __413921_413921;
   reg _413922_413922 ; 
   reg __413922_413922;
   reg _413923_413923 ; 
   reg __413923_413923;
   reg _413924_413924 ; 
   reg __413924_413924;
   reg _413925_413925 ; 
   reg __413925_413925;
   reg _413926_413926 ; 
   reg __413926_413926;
   reg _413927_413927 ; 
   reg __413927_413927;
   reg _413928_413928 ; 
   reg __413928_413928;
   reg _413929_413929 ; 
   reg __413929_413929;
   reg _413930_413930 ; 
   reg __413930_413930;
   reg _413931_413931 ; 
   reg __413931_413931;
   reg _413932_413932 ; 
   reg __413932_413932;
   reg _413933_413933 ; 
   reg __413933_413933;
   reg _413934_413934 ; 
   reg __413934_413934;
   reg _413935_413935 ; 
   reg __413935_413935;
   reg _413936_413936 ; 
   reg __413936_413936;
   reg _413937_413937 ; 
   reg __413937_413937;
   reg _413938_413938 ; 
   reg __413938_413938;
   reg _413939_413939 ; 
   reg __413939_413939;
   reg _413940_413940 ; 
   reg __413940_413940;
   reg _413941_413941 ; 
   reg __413941_413941;
   reg _413942_413942 ; 
   reg __413942_413942;
   reg _413943_413943 ; 
   reg __413943_413943;
   reg _413944_413944 ; 
   reg __413944_413944;
   reg _413945_413945 ; 
   reg __413945_413945;
   reg _413946_413946 ; 
   reg __413946_413946;
   reg _413947_413947 ; 
   reg __413947_413947;
   reg _413948_413948 ; 
   reg __413948_413948;
   reg _413949_413949 ; 
   reg __413949_413949;
   reg _413950_413950 ; 
   reg __413950_413950;
   reg _413951_413951 ; 
   reg __413951_413951;
   reg _413952_413952 ; 
   reg __413952_413952;
   reg _413953_413953 ; 
   reg __413953_413953;
   reg _413954_413954 ; 
   reg __413954_413954;
   reg _413955_413955 ; 
   reg __413955_413955;
   reg _413956_413956 ; 
   reg __413956_413956;
   reg _413957_413957 ; 
   reg __413957_413957;
   reg _413958_413958 ; 
   reg __413958_413958;
   reg _413959_413959 ; 
   reg __413959_413959;
   reg _413960_413960 ; 
   reg __413960_413960;
   reg _413961_413961 ; 
   reg __413961_413961;
   reg _413962_413962 ; 
   reg __413962_413962;
   reg _413963_413963 ; 
   reg __413963_413963;
   reg _413964_413964 ; 
   reg __413964_413964;
   reg _413965_413965 ; 
   reg __413965_413965;
   reg _413966_413966 ; 
   reg __413966_413966;
   reg _413967_413967 ; 
   reg __413967_413967;
   reg _413968_413968 ; 
   reg __413968_413968;
   reg _413969_413969 ; 
   reg __413969_413969;
   reg _413970_413970 ; 
   reg __413970_413970;
   reg _413971_413971 ; 
   reg __413971_413971;
   reg _413972_413972 ; 
   reg __413972_413972;
   reg _413973_413973 ; 
   reg __413973_413973;
   reg _413974_413974 ; 
   reg __413974_413974;
   reg _413975_413975 ; 
   reg __413975_413975;
   reg _413976_413976 ; 
   reg __413976_413976;
   reg _413977_413977 ; 
   reg __413977_413977;
   reg _413978_413978 ; 
   reg __413978_413978;
   reg _413979_413979 ; 
   reg __413979_413979;
   reg _413980_413980 ; 
   reg __413980_413980;
   reg _413981_413981 ; 
   reg __413981_413981;
   reg _413982_413982 ; 
   reg __413982_413982;
   reg _413983_413983 ; 
   reg __413983_413983;
   reg _413984_413984 ; 
   reg __413984_413984;
   reg _413985_413985 ; 
   reg __413985_413985;
   reg _413986_413986 ; 
   reg __413986_413986;
   reg _413987_413987 ; 
   reg __413987_413987;
   reg _413988_413988 ; 
   reg __413988_413988;
   reg _413989_413989 ; 
   reg __413989_413989;
   reg _413990_413990 ; 
   reg __413990_413990;
   reg _413991_413991 ; 
   reg __413991_413991;
   reg _413992_413992 ; 
   reg __413992_413992;
   reg _413993_413993 ; 
   reg __413993_413993;
   reg _413994_413994 ; 
   reg __413994_413994;
   reg _413995_413995 ; 
   reg __413995_413995;
   reg _413996_413996 ; 
   reg __413996_413996;
   reg _413997_413997 ; 
   reg __413997_413997;
   reg _413998_413998 ; 
   reg __413998_413998;
   reg _413999_413999 ; 
   reg __413999_413999;
   reg _414000_414000 ; 
   reg __414000_414000;
   reg _414001_414001 ; 
   reg __414001_414001;
   reg _414002_414002 ; 
   reg __414002_414002;
   reg _414003_414003 ; 
   reg __414003_414003;
   reg _414004_414004 ; 
   reg __414004_414004;
   reg _414005_414005 ; 
   reg __414005_414005;
   reg _414006_414006 ; 
   reg __414006_414006;
   reg _414007_414007 ; 
   reg __414007_414007;
   reg _414008_414008 ; 
   reg __414008_414008;
   reg _414009_414009 ; 
   reg __414009_414009;
   reg _414010_414010 ; 
   reg __414010_414010;
   reg _414011_414011 ; 
   reg __414011_414011;
   reg _414012_414012 ; 
   reg __414012_414012;
   reg _414013_414013 ; 
   reg __414013_414013;
   reg _414014_414014 ; 
   reg __414014_414014;
   reg _414015_414015 ; 
   reg __414015_414015;
   reg _414016_414016 ; 
   reg __414016_414016;
   reg _414017_414017 ; 
   reg __414017_414017;
   reg _414018_414018 ; 
   reg __414018_414018;
   reg _414019_414019 ; 
   reg __414019_414019;
   reg _414020_414020 ; 
   reg __414020_414020;
   reg _414021_414021 ; 
   reg __414021_414021;
   reg _414022_414022 ; 
   reg __414022_414022;
   reg _414023_414023 ; 
   reg __414023_414023;
   reg _414024_414024 ; 
   reg __414024_414024;
   reg _414025_414025 ; 
   reg __414025_414025;
   reg _414026_414026 ; 
   reg __414026_414026;
   reg _414027_414027 ; 
   reg __414027_414027;
   reg _414028_414028 ; 
   reg __414028_414028;
   reg _414029_414029 ; 
   reg __414029_414029;
   reg _414030_414030 ; 
   reg __414030_414030;
   reg _414031_414031 ; 
   reg __414031_414031;
   reg _414032_414032 ; 
   reg __414032_414032;
   reg _414033_414033 ; 
   reg __414033_414033;
   reg _414034_414034 ; 
   reg __414034_414034;
   reg _414035_414035 ; 
   reg __414035_414035;
   reg _414036_414036 ; 
   reg __414036_414036;
   reg _414037_414037 ; 
   reg __414037_414037;
   reg _414038_414038 ; 
   reg __414038_414038;
   reg _414039_414039 ; 
   reg __414039_414039;
   reg _414040_414040 ; 
   reg __414040_414040;
   reg _414041_414041 ; 
   reg __414041_414041;
   reg _414042_414042 ; 
   reg __414042_414042;
   reg _414043_414043 ; 
   reg __414043_414043;
   reg _414044_414044 ; 
   reg __414044_414044;
   reg _414045_414045 ; 
   reg __414045_414045;
   reg _414046_414046 ; 
   reg __414046_414046;
   reg _414047_414047 ; 
   reg __414047_414047;
   reg _414048_414048 ; 
   reg __414048_414048;
   reg _414049_414049 ; 
   reg __414049_414049;
   reg _414050_414050 ; 
   reg __414050_414050;
   reg _414051_414051 ; 
   reg __414051_414051;
   reg _414052_414052 ; 
   reg __414052_414052;
   reg _414053_414053 ; 
   reg __414053_414053;
   reg _414054_414054 ; 
   reg __414054_414054;
   reg _414055_414055 ; 
   reg __414055_414055;
   reg _414056_414056 ; 
   reg __414056_414056;
   reg _414057_414057 ; 
   reg __414057_414057;
   reg _414058_414058 ; 
   reg __414058_414058;
   reg _414059_414059 ; 
   reg __414059_414059;
   reg _414060_414060 ; 
   reg __414060_414060;
   reg _414061_414061 ; 
   reg __414061_414061;
   reg _414062_414062 ; 
   reg __414062_414062;
   reg _414063_414063 ; 
   reg __414063_414063;
   reg _414064_414064 ; 
   reg __414064_414064;
   reg _414065_414065 ; 
   reg __414065_414065;
   reg _414066_414066 ; 
   reg __414066_414066;
   reg _414067_414067 ; 
   reg __414067_414067;
   reg _414068_414068 ; 
   reg __414068_414068;
   reg _414069_414069 ; 
   reg __414069_414069;
   reg _414070_414070 ; 
   reg __414070_414070;
   reg _414071_414071 ; 
   reg __414071_414071;
   reg _414072_414072 ; 
   reg __414072_414072;
   reg _414073_414073 ; 
   reg __414073_414073;
   reg _414074_414074 ; 
   reg __414074_414074;
   reg _414075_414075 ; 
   reg __414075_414075;
   reg _414076_414076 ; 
   reg __414076_414076;
   reg _414077_414077 ; 
   reg __414077_414077;
   reg _414078_414078 ; 
   reg __414078_414078;
   reg _414079_414079 ; 
   reg __414079_414079;
   reg _414080_414080 ; 
   reg __414080_414080;
   reg _414081_414081 ; 
   reg __414081_414081;
   reg _414082_414082 ; 
   reg __414082_414082;
   reg _414083_414083 ; 
   reg __414083_414083;
   reg _414084_414084 ; 
   reg __414084_414084;
   reg _414085_414085 ; 
   reg __414085_414085;
   reg _414086_414086 ; 
   reg __414086_414086;
   reg _414087_414087 ; 
   reg __414087_414087;
   reg _414088_414088 ; 
   reg __414088_414088;
   reg _414089_414089 ; 
   reg __414089_414089;
   reg _414090_414090 ; 
   reg __414090_414090;
   reg _414091_414091 ; 
   reg __414091_414091;
   reg _414092_414092 ; 
   reg __414092_414092;
   reg _414093_414093 ; 
   reg __414093_414093;
   reg _414094_414094 ; 
   reg __414094_414094;
   reg _414095_414095 ; 
   reg __414095_414095;
   reg _414096_414096 ; 
   reg __414096_414096;
   reg _414097_414097 ; 
   reg __414097_414097;
   reg _414098_414098 ; 
   reg __414098_414098;
   reg _414099_414099 ; 
   reg __414099_414099;
   reg _414100_414100 ; 
   reg __414100_414100;
   reg _414101_414101 ; 
   reg __414101_414101;
   reg _414102_414102 ; 
   reg __414102_414102;
   reg _414103_414103 ; 
   reg __414103_414103;
   reg _414104_414104 ; 
   reg __414104_414104;
   reg _414105_414105 ; 
   reg __414105_414105;
   reg _414106_414106 ; 
   reg __414106_414106;
   reg _414107_414107 ; 
   reg __414107_414107;
   reg _414108_414108 ; 
   reg __414108_414108;
   reg _414109_414109 ; 
   reg __414109_414109;
   reg _414110_414110 ; 
   reg __414110_414110;
   reg _414111_414111 ; 
   reg __414111_414111;
   reg _414112_414112 ; 
   reg __414112_414112;
   reg _414113_414113 ; 
   reg __414113_414113;
   reg _414114_414114 ; 
   reg __414114_414114;
   reg _414115_414115 ; 
   reg __414115_414115;
   reg _414116_414116 ; 
   reg __414116_414116;
   reg _414117_414117 ; 
   reg __414117_414117;
   reg _414118_414118 ; 
   reg __414118_414118;
   reg _414119_414119 ; 
   reg __414119_414119;
   reg _414120_414120 ; 
   reg __414120_414120;
   reg _414121_414121 ; 
   reg __414121_414121;
   reg _414122_414122 ; 
   reg __414122_414122;
   reg _414123_414123 ; 
   reg __414123_414123;
   reg _414124_414124 ; 
   reg __414124_414124;
   reg _414125_414125 ; 
   reg __414125_414125;
   reg _414126_414126 ; 
   reg __414126_414126;
   reg _414127_414127 ; 
   reg __414127_414127;
   reg _414128_414128 ; 
   reg __414128_414128;
   reg _414129_414129 ; 
   reg __414129_414129;
   reg _414130_414130 ; 
   reg __414130_414130;
   reg _414131_414131 ; 
   reg __414131_414131;
   reg _414132_414132 ; 
   reg __414132_414132;
   reg _414133_414133 ; 
   reg __414133_414133;
   reg _414134_414134 ; 
   reg __414134_414134;
   reg _414135_414135 ; 
   reg __414135_414135;
   reg _414136_414136 ; 
   reg __414136_414136;
   reg _414137_414137 ; 
   reg __414137_414137;
   reg _414138_414138 ; 
   reg __414138_414138;
   reg _414139_414139 ; 
   reg __414139_414139;
   reg _414140_414140 ; 
   reg __414140_414140;
   reg _414141_414141 ; 
   reg __414141_414141;
   reg _414142_414142 ; 
   reg __414142_414142;
   reg _414143_414143 ; 
   reg __414143_414143;
   reg _414144_414144 ; 
   reg __414144_414144;
   reg _414145_414145 ; 
   reg __414145_414145;
   reg _414146_414146 ; 
   reg __414146_414146;
   reg _414147_414147 ; 
   reg __414147_414147;
   reg _414148_414148 ; 
   reg __414148_414148;
   reg _414149_414149 ; 
   reg __414149_414149;
   reg _414150_414150 ; 
   reg __414150_414150;
   reg _414151_414151 ; 
   reg __414151_414151;
   reg _414152_414152 ; 
   reg __414152_414152;
   reg _414153_414153 ; 
   reg __414153_414153;
   reg _414154_414154 ; 
   reg __414154_414154;
   reg _414155_414155 ; 
   reg __414155_414155;
   reg _414156_414156 ; 
   reg __414156_414156;
   reg _414157_414157 ; 
   reg __414157_414157;
   reg _414158_414158 ; 
   reg __414158_414158;
   reg _414159_414159 ; 
   reg __414159_414159;
   reg _414160_414160 ; 
   reg __414160_414160;
   reg _414161_414161 ; 
   reg __414161_414161;
   reg _414162_414162 ; 
   reg __414162_414162;
   reg _414163_414163 ; 
   reg __414163_414163;
   reg _414164_414164 ; 
   reg __414164_414164;
   reg _414165_414165 ; 
   reg __414165_414165;
   reg _414166_414166 ; 
   reg __414166_414166;
   reg _414167_414167 ; 
   reg __414167_414167;
   reg _414168_414168 ; 
   reg __414168_414168;
   reg _414169_414169 ; 
   reg __414169_414169;
   reg _414170_414170 ; 
   reg __414170_414170;
   reg _414171_414171 ; 
   reg __414171_414171;
   reg _414172_414172 ; 
   reg __414172_414172;
   reg _414173_414173 ; 
   reg __414173_414173;
   reg _414174_414174 ; 
   reg __414174_414174;
   reg _414175_414175 ; 
   reg __414175_414175;
   reg _414176_414176 ; 
   reg __414176_414176;
   reg _414177_414177 ; 
   reg __414177_414177;
   reg _414178_414178 ; 
   reg __414178_414178;
   reg _414179_414179 ; 
   reg __414179_414179;
   reg _414180_414180 ; 
   reg __414180_414180;
   reg _414181_414181 ; 
   reg __414181_414181;
   reg _414182_414182 ; 
   reg __414182_414182;
   reg _414183_414183 ; 
   reg __414183_414183;
   reg _414184_414184 ; 
   reg __414184_414184;
   reg _414185_414185 ; 
   reg __414185_414185;
   reg _414186_414186 ; 
   reg __414186_414186;
   reg _414187_414187 ; 
   reg __414187_414187;
   reg _414188_414188 ; 
   reg __414188_414188;
   reg _414189_414189 ; 
   reg __414189_414189;
   reg _414190_414190 ; 
   reg __414190_414190;
   reg _414191_414191 ; 
   reg __414191_414191;
   reg _414192_414192 ; 
   reg __414192_414192;
   reg _414193_414193 ; 
   reg __414193_414193;
   reg _414194_414194 ; 
   reg __414194_414194;
   reg _414195_414195 ; 
   reg __414195_414195;
   reg _414196_414196 ; 
   reg __414196_414196;
   reg _414197_414197 ; 
   reg __414197_414197;
   reg _414198_414198 ; 
   reg __414198_414198;
   reg _414199_414199 ; 
   reg __414199_414199;
   reg _414200_414200 ; 
   reg __414200_414200;
   reg _414201_414201 ; 
   reg __414201_414201;
   reg _414202_414202 ; 
   reg __414202_414202;
   reg _414203_414203 ; 
   reg __414203_414203;
   reg _414204_414204 ; 
   reg __414204_414204;
   reg _414205_414205 ; 
   reg __414205_414205;
   reg _414206_414206 ; 
   reg __414206_414206;
   reg _414207_414207 ; 
   reg __414207_414207;
   reg _414208_414208 ; 
   reg __414208_414208;
   reg _414209_414209 ; 
   reg __414209_414209;
   reg _414210_414210 ; 
   reg __414210_414210;
   reg _414211_414211 ; 
   reg __414211_414211;
   reg _414212_414212 ; 
   reg __414212_414212;
   reg _414213_414213 ; 
   reg __414213_414213;
   reg _414214_414214 ; 
   reg __414214_414214;
   reg _414215_414215 ; 
   reg __414215_414215;
   reg _414216_414216 ; 
   reg __414216_414216;
   reg _414217_414217 ; 
   reg __414217_414217;
   reg _414218_414218 ; 
   reg __414218_414218;
   reg _414219_414219 ; 
   reg __414219_414219;
   reg _414220_414220 ; 
   reg __414220_414220;
   reg _414221_414221 ; 
   reg __414221_414221;
   reg _414222_414222 ; 
   reg __414222_414222;
   reg _414223_414223 ; 
   reg __414223_414223;
   reg _414224_414224 ; 
   reg __414224_414224;
   reg _414225_414225 ; 
   reg __414225_414225;
   reg _414226_414226 ; 
   reg __414226_414226;
   reg _414227_414227 ; 
   reg __414227_414227;
   reg _414228_414228 ; 
   reg __414228_414228;
   reg _414229_414229 ; 
   reg __414229_414229;
   reg _414230_414230 ; 
   reg __414230_414230;
   reg _414231_414231 ; 
   reg __414231_414231;
   reg _414232_414232 ; 
   reg __414232_414232;
   reg _414233_414233 ; 
   reg __414233_414233;
   reg _414234_414234 ; 
   reg __414234_414234;
   reg _414235_414235 ; 
   reg __414235_414235;
   reg _414236_414236 ; 
   reg __414236_414236;
   reg _414237_414237 ; 
   reg __414237_414237;
   reg _414238_414238 ; 
   reg __414238_414238;
   reg _414239_414239 ; 
   reg __414239_414239;
   reg _414240_414240 ; 
   reg __414240_414240;
   reg _414241_414241 ; 
   reg __414241_414241;
   reg _414242_414242 ; 
   reg __414242_414242;
   reg _414243_414243 ; 
   reg __414243_414243;
   reg _414244_414244 ; 
   reg __414244_414244;
   reg _414245_414245 ; 
   reg __414245_414245;
   reg _414246_414246 ; 
   reg __414246_414246;
   reg _414247_414247 ; 
   reg __414247_414247;
   reg _414248_414248 ; 
   reg __414248_414248;
   reg _414249_414249 ; 
   reg __414249_414249;
   reg _414250_414250 ; 
   reg __414250_414250;
   reg _414251_414251 ; 
   reg __414251_414251;
   reg _414252_414252 ; 
   reg __414252_414252;
   reg _414253_414253 ; 
   reg __414253_414253;
   reg _414254_414254 ; 
   reg __414254_414254;
   reg _414255_414255 ; 
   reg __414255_414255;
   reg _414256_414256 ; 
   reg __414256_414256;
   reg _414257_414257 ; 
   reg __414257_414257;
   reg _414258_414258 ; 
   reg __414258_414258;
   reg _414259_414259 ; 
   reg __414259_414259;
   reg _414260_414260 ; 
   reg __414260_414260;
   reg _414261_414261 ; 
   reg __414261_414261;
   reg _414262_414262 ; 
   reg __414262_414262;
   reg _414263_414263 ; 
   reg __414263_414263;
   reg _414264_414264 ; 
   reg __414264_414264;
   reg _414265_414265 ; 
   reg __414265_414265;
   reg _414266_414266 ; 
   reg __414266_414266;
   reg _414267_414267 ; 
   reg __414267_414267;
   reg _414268_414268 ; 
   reg __414268_414268;
   reg _414269_414269 ; 
   reg __414269_414269;
   reg _414270_414270 ; 
   reg __414270_414270;
   reg _414271_414271 ; 
   reg __414271_414271;
   reg _414272_414272 ; 
   reg __414272_414272;
   reg _414273_414273 ; 
   reg __414273_414273;
   reg _414274_414274 ; 
   reg __414274_414274;
   reg _414275_414275 ; 
   reg __414275_414275;
   reg _414276_414276 ; 
   reg __414276_414276;
   reg _414277_414277 ; 
   reg __414277_414277;
   reg _414278_414278 ; 
   reg __414278_414278;
   reg _414279_414279 ; 
   reg __414279_414279;
   reg _414280_414280 ; 
   reg __414280_414280;
   reg _414281_414281 ; 
   reg __414281_414281;
   reg _414282_414282 ; 
   reg __414282_414282;
   reg _414283_414283 ; 
   reg __414283_414283;
   reg _414284_414284 ; 
   reg __414284_414284;
   reg _414285_414285 ; 
   reg __414285_414285;
   reg _414286_414286 ; 
   reg __414286_414286;
   reg _414287_414287 ; 
   reg __414287_414287;
   reg _414288_414288 ; 
   reg __414288_414288;
   reg _414289_414289 ; 
   reg __414289_414289;
   reg _414290_414290 ; 
   reg __414290_414290;
   reg _414291_414291 ; 
   reg __414291_414291;
   reg _414292_414292 ; 
   reg __414292_414292;
   reg _414293_414293 ; 
   reg __414293_414293;
   reg _414294_414294 ; 
   reg __414294_414294;
   reg _414295_414295 ; 
   reg __414295_414295;
   reg _414296_414296 ; 
   reg __414296_414296;
   reg _414297_414297 ; 
   reg __414297_414297;
   reg _414298_414298 ; 
   reg __414298_414298;
   reg _414299_414299 ; 
   reg __414299_414299;
   reg _414300_414300 ; 
   reg __414300_414300;
   reg _414301_414301 ; 
   reg __414301_414301;
   reg _414302_414302 ; 
   reg __414302_414302;
   reg _414303_414303 ; 
   reg __414303_414303;
   reg _414304_414304 ; 
   reg __414304_414304;
   reg _414305_414305 ; 
   reg __414305_414305;
   reg _414306_414306 ; 
   reg __414306_414306;
   reg _414307_414307 ; 
   reg __414307_414307;
   reg _414308_414308 ; 
   reg __414308_414308;
   reg _414309_414309 ; 
   reg __414309_414309;
   reg _414310_414310 ; 
   reg __414310_414310;
   reg _414311_414311 ; 
   reg __414311_414311;
   reg _414312_414312 ; 
   reg __414312_414312;
   reg _414313_414313 ; 
   reg __414313_414313;
   reg _414314_414314 ; 
   reg __414314_414314;
   reg _414315_414315 ; 
   reg __414315_414315;
   reg _414316_414316 ; 
   reg __414316_414316;
   reg _414317_414317 ; 
   reg __414317_414317;
   reg _414318_414318 ; 
   reg __414318_414318;
   reg _414319_414319 ; 
   reg __414319_414319;
   reg _414320_414320 ; 
   reg __414320_414320;
   reg _414321_414321 ; 
   reg __414321_414321;
   reg _414322_414322 ; 
   reg __414322_414322;
   reg _414323_414323 ; 
   reg __414323_414323;
   reg _414324_414324 ; 
   reg __414324_414324;
   reg _414325_414325 ; 
   reg __414325_414325;
   reg _414326_414326 ; 
   reg __414326_414326;
   reg _414327_414327 ; 
   reg __414327_414327;
   reg _414328_414328 ; 
   reg __414328_414328;
   reg _414329_414329 ; 
   reg __414329_414329;
   reg _414330_414330 ; 
   reg __414330_414330;
   reg _414331_414331 ; 
   reg __414331_414331;
   reg _414332_414332 ; 
   reg __414332_414332;
   reg _414333_414333 ; 
   reg __414333_414333;
   reg _414334_414334 ; 
   reg __414334_414334;
   reg _414335_414335 ; 
   reg __414335_414335;
   reg _414336_414336 ; 
   reg __414336_414336;
   reg _414337_414337 ; 
   reg __414337_414337;
   reg _414338_414338 ; 
   reg __414338_414338;
   reg _414339_414339 ; 
   reg __414339_414339;
   reg _414340_414340 ; 
   reg __414340_414340;
   reg _414341_414341 ; 
   reg __414341_414341;
   reg _414342_414342 ; 
   reg __414342_414342;
   reg _414343_414343 ; 
   reg __414343_414343;
   reg _414344_414344 ; 
   reg __414344_414344;
   reg _414345_414345 ; 
   reg __414345_414345;
   reg _414346_414346 ; 
   reg __414346_414346;
   reg _414347_414347 ; 
   reg __414347_414347;
   reg _414348_414348 ; 
   reg __414348_414348;
   reg _414349_414349 ; 
   reg __414349_414349;
   reg _414350_414350 ; 
   reg __414350_414350;
   reg _414351_414351 ; 
   reg __414351_414351;
   reg _414352_414352 ; 
   reg __414352_414352;
   reg _414353_414353 ; 
   reg __414353_414353;
   reg _414354_414354 ; 
   reg __414354_414354;
   reg _414355_414355 ; 
   reg __414355_414355;
   reg _414356_414356 ; 
   reg __414356_414356;
   reg _414357_414357 ; 
   reg __414357_414357;
   reg _414358_414358 ; 
   reg __414358_414358;
   reg _414359_414359 ; 
   reg __414359_414359;
   reg _414360_414360 ; 
   reg __414360_414360;
   reg _414361_414361 ; 
   reg __414361_414361;
   reg _414362_414362 ; 
   reg __414362_414362;
   reg _414363_414363 ; 
   reg __414363_414363;
   reg _414364_414364 ; 
   reg __414364_414364;
   reg _414365_414365 ; 
   reg __414365_414365;
   reg _414366_414366 ; 
   reg __414366_414366;
   reg _414367_414367 ; 
   reg __414367_414367;
   reg _414368_414368 ; 
   reg __414368_414368;
   reg _414369_414369 ; 
   reg __414369_414369;
   reg _414370_414370 ; 
   reg __414370_414370;
   reg _414371_414371 ; 
   reg __414371_414371;
   reg _414372_414372 ; 
   reg __414372_414372;
   reg _414373_414373 ; 
   reg __414373_414373;
   reg _414374_414374 ; 
   reg __414374_414374;
   reg _414375_414375 ; 
   reg __414375_414375;
   reg _414376_414376 ; 
   reg __414376_414376;
   reg _414377_414377 ; 
   reg __414377_414377;
   reg _414378_414378 ; 
   reg __414378_414378;
   reg _414379_414379 ; 
   reg __414379_414379;
   reg _414380_414380 ; 
   reg __414380_414380;
   reg _414381_414381 ; 
   reg __414381_414381;
   reg _414382_414382 ; 
   reg __414382_414382;
   reg _414383_414383 ; 
   reg __414383_414383;
   reg _414384_414384 ; 
   reg __414384_414384;
   reg _414385_414385 ; 
   reg __414385_414385;
   reg _414386_414386 ; 
   reg __414386_414386;
   reg _414387_414387 ; 
   reg __414387_414387;
   reg _414388_414388 ; 
   reg __414388_414388;
   reg _414389_414389 ; 
   reg __414389_414389;
   reg _414390_414390 ; 
   reg __414390_414390;
   reg _414391_414391 ; 
   reg __414391_414391;
   reg _414392_414392 ; 
   reg __414392_414392;
   reg _414393_414393 ; 
   reg __414393_414393;
   reg _414394_414394 ; 
   reg __414394_414394;
   reg _414395_414395 ; 
   reg __414395_414395;
   reg _414396_414396 ; 
   reg __414396_414396;
   reg _414397_414397 ; 
   reg __414397_414397;
   reg _414398_414398 ; 
   reg __414398_414398;
   reg _414399_414399 ; 
   reg __414399_414399;
   reg _414400_414400 ; 
   reg __414400_414400;
   reg _414401_414401 ; 
   reg __414401_414401;
   reg _414402_414402 ; 
   reg __414402_414402;
   reg _414403_414403 ; 
   reg __414403_414403;
   reg _414404_414404 ; 
   reg __414404_414404;
   reg _414405_414405 ; 
   reg __414405_414405;
   reg _414406_414406 ; 
   reg __414406_414406;
   reg _414407_414407 ; 
   reg __414407_414407;
   reg _414408_414408 ; 
   reg __414408_414408;
   reg _414409_414409 ; 
   reg __414409_414409;
   reg _414410_414410 ; 
   reg __414410_414410;
   reg _414411_414411 ; 
   reg __414411_414411;
   reg _414412_414412 ; 
   reg __414412_414412;
   reg _414413_414413 ; 
   reg __414413_414413;
   reg _414414_414414 ; 
   reg __414414_414414;
   reg _414415_414415 ; 
   reg __414415_414415;
   reg _414416_414416 ; 
   reg __414416_414416;
   reg _414417_414417 ; 
   reg __414417_414417;
   reg _414418_414418 ; 
   reg __414418_414418;
   reg _414419_414419 ; 
   reg __414419_414419;
   reg _414420_414420 ; 
   reg __414420_414420;
   reg _414421_414421 ; 
   reg __414421_414421;
   reg _414422_414422 ; 
   reg __414422_414422;
   reg _414423_414423 ; 
   reg __414423_414423;
   reg _414424_414424 ; 
   reg __414424_414424;
   reg _414425_414425 ; 
   reg __414425_414425;
   reg _414426_414426 ; 
   reg __414426_414426;
   reg _414427_414427 ; 
   reg __414427_414427;
   reg _414428_414428 ; 
   reg __414428_414428;
   reg _414429_414429 ; 
   reg __414429_414429;
   reg _414430_414430 ; 
   reg __414430_414430;
   reg _414431_414431 ; 
   reg __414431_414431;
   reg _414432_414432 ; 
   reg __414432_414432;
   reg _414433_414433 ; 
   reg __414433_414433;
   reg _414434_414434 ; 
   reg __414434_414434;
   reg _414435_414435 ; 
   reg __414435_414435;
   reg _414436_414436 ; 
   reg __414436_414436;
   reg _414437_414437 ; 
   reg __414437_414437;
   reg _414438_414438 ; 
   reg __414438_414438;
   reg _414439_414439 ; 
   reg __414439_414439;
   reg _414440_414440 ; 
   reg __414440_414440;
   reg _414441_414441 ; 
   reg __414441_414441;
   reg _414442_414442 ; 
   reg __414442_414442;
   reg _414443_414443 ; 
   reg __414443_414443;
   reg _414444_414444 ; 
   reg __414444_414444;
   reg _414445_414445 ; 
   reg __414445_414445;
   reg _414446_414446 ; 
   reg __414446_414446;
   reg _414447_414447 ; 
   reg __414447_414447;
   reg _414448_414448 ; 
   reg __414448_414448;
   reg _414449_414449 ; 
   reg __414449_414449;
   reg _414450_414450 ; 
   reg __414450_414450;
   reg _414451_414451 ; 
   reg __414451_414451;
   reg _414452_414452 ; 
   reg __414452_414452;
   reg _414453_414453 ; 
   reg __414453_414453;
   reg _414454_414454 ; 
   reg __414454_414454;
   reg _414455_414455 ; 
   reg __414455_414455;
   reg _414456_414456 ; 
   reg __414456_414456;
   reg _414457_414457 ; 
   reg __414457_414457;
   reg _414458_414458 ; 
   reg __414458_414458;
   reg _414459_414459 ; 
   reg __414459_414459;
   reg _414460_414460 ; 
   reg __414460_414460;
   reg _414461_414461 ; 
   reg __414461_414461;
   reg _414462_414462 ; 
   reg __414462_414462;
   reg _414463_414463 ; 
   reg __414463_414463;
   reg _414464_414464 ; 
   reg __414464_414464;
   reg _414465_414465 ; 
   reg __414465_414465;
   reg _414466_414466 ; 
   reg __414466_414466;
   reg _414467_414467 ; 
   reg __414467_414467;
   reg _414468_414468 ; 
   reg __414468_414468;
   reg _414469_414469 ; 
   reg __414469_414469;
   reg _414470_414470 ; 
   reg __414470_414470;
   reg _414471_414471 ; 
   reg __414471_414471;
   reg _414472_414472 ; 
   reg __414472_414472;
   reg _414473_414473 ; 
   reg __414473_414473;
   reg _414474_414474 ; 
   reg __414474_414474;
   reg _414475_414475 ; 
   reg __414475_414475;
   reg _414476_414476 ; 
   reg __414476_414476;
   reg _414477_414477 ; 
   reg __414477_414477;
   reg _414478_414478 ; 
   reg __414478_414478;
   reg _414479_414479 ; 
   reg __414479_414479;
   reg _414480_414480 ; 
   reg __414480_414480;
   reg _414481_414481 ; 
   reg __414481_414481;
   reg _414482_414482 ; 
   reg __414482_414482;
   reg _414483_414483 ; 
   reg __414483_414483;
   reg _414484_414484 ; 
   reg __414484_414484;
   reg _414485_414485 ; 
   reg __414485_414485;
   reg _414486_414486 ; 
   reg __414486_414486;
   reg _414487_414487 ; 
   reg __414487_414487;
   reg _414488_414488 ; 
   reg __414488_414488;
   reg _414489_414489 ; 
   reg __414489_414489;
   reg _414490_414490 ; 
   reg __414490_414490;
   reg _414491_414491 ; 
   reg __414491_414491;
   reg _414492_414492 ; 
   reg __414492_414492;
   reg _414493_414493 ; 
   reg __414493_414493;
   reg _414494_414494 ; 
   reg __414494_414494;
   reg _414495_414495 ; 
   reg __414495_414495;
   reg _414496_414496 ; 
   reg __414496_414496;
   reg _414497_414497 ; 
   reg __414497_414497;
   reg _414498_414498 ; 
   reg __414498_414498;
   reg _414499_414499 ; 
   reg __414499_414499;
   reg _414500_414500 ; 
   reg __414500_414500;
   reg _414501_414501 ; 
   reg __414501_414501;
   reg _414502_414502 ; 
   reg __414502_414502;
   reg _414503_414503 ; 
   reg __414503_414503;
   reg _414504_414504 ; 
   reg __414504_414504;
   reg _414505_414505 ; 
   reg __414505_414505;
   reg _414506_414506 ; 
   reg __414506_414506;
   reg _414507_414507 ; 
   reg __414507_414507;
   reg _414508_414508 ; 
   reg __414508_414508;
   reg _414509_414509 ; 
   reg __414509_414509;
   reg _414510_414510 ; 
   reg __414510_414510;
   reg _414511_414511 ; 
   reg __414511_414511;
   reg _414512_414512 ; 
   reg __414512_414512;
   reg _414513_414513 ; 
   reg __414513_414513;
   reg _414514_414514 ; 
   reg __414514_414514;
   reg _414515_414515 ; 
   reg __414515_414515;
   reg _414516_414516 ; 
   reg __414516_414516;
   reg _414517_414517 ; 
   reg __414517_414517;
   reg _414518_414518 ; 
   reg __414518_414518;
   reg _414519_414519 ; 
   reg __414519_414519;
   reg _414520_414520 ; 
   reg __414520_414520;
   reg _414521_414521 ; 
   reg __414521_414521;
   reg _414522_414522 ; 
   reg __414522_414522;
   reg _414523_414523 ; 
   reg __414523_414523;
   reg _414524_414524 ; 
   reg __414524_414524;
   reg _414525_414525 ; 
   reg __414525_414525;
   reg _414526_414526 ; 
   reg __414526_414526;
   reg _414527_414527 ; 
   reg __414527_414527;
   reg _414528_414528 ; 
   reg __414528_414528;
   reg _414529_414529 ; 
   reg __414529_414529;
   reg _414530_414530 ; 
   reg __414530_414530;
   reg _414531_414531 ; 
   reg __414531_414531;
   reg _414532_414532 ; 
   reg __414532_414532;
   reg _414533_414533 ; 
   reg __414533_414533;
   reg _414534_414534 ; 
   reg __414534_414534;
   reg _414535_414535 ; 
   reg __414535_414535;
   reg _414536_414536 ; 
   reg __414536_414536;
   reg _414537_414537 ; 
   reg __414537_414537;
   reg _414538_414538 ; 
   reg __414538_414538;
   reg _414539_414539 ; 
   reg __414539_414539;
   reg _414540_414540 ; 
   reg __414540_414540;
   reg _414541_414541 ; 
   reg __414541_414541;
   reg _414542_414542 ; 
   reg __414542_414542;
   reg _414543_414543 ; 
   reg __414543_414543;
   reg _414544_414544 ; 
   reg __414544_414544;
   reg _414545_414545 ; 
   reg __414545_414545;
   reg _414546_414546 ; 
   reg __414546_414546;
   reg _414547_414547 ; 
   reg __414547_414547;
   reg _414548_414548 ; 
   reg __414548_414548;
   reg _414549_414549 ; 
   reg __414549_414549;
   reg _414550_414550 ; 
   reg __414550_414550;
   reg _414551_414551 ; 
   reg __414551_414551;
   reg _414552_414552 ; 
   reg __414552_414552;
   reg _414553_414553 ; 
   reg __414553_414553;
   reg _414554_414554 ; 
   reg __414554_414554;
   reg _414555_414555 ; 
   reg __414555_414555;
   reg _414556_414556 ; 
   reg __414556_414556;
   reg _414557_414557 ; 
   reg __414557_414557;
   reg _414558_414558 ; 
   reg __414558_414558;
   reg _414559_414559 ; 
   reg __414559_414559;
   reg _414560_414560 ; 
   reg __414560_414560;
   reg _414561_414561 ; 
   reg __414561_414561;
   reg _414562_414562 ; 
   reg __414562_414562;
   reg _414563_414563 ; 
   reg __414563_414563;
   reg _414564_414564 ; 
   reg __414564_414564;
   reg _414565_414565 ; 
   reg __414565_414565;
   reg _414566_414566 ; 
   reg __414566_414566;
   reg _414567_414567 ; 
   reg __414567_414567;
   reg _414568_414568 ; 
   reg __414568_414568;
   reg _414569_414569 ; 
   reg __414569_414569;
   reg _414570_414570 ; 
   reg __414570_414570;
   reg _414571_414571 ; 
   reg __414571_414571;
   reg _414572_414572 ; 
   reg __414572_414572;
   reg _414573_414573 ; 
   reg __414573_414573;
   reg _414574_414574 ; 
   reg __414574_414574;
   reg _414575_414575 ; 
   reg __414575_414575;
   reg _414576_414576 ; 
   reg __414576_414576;
   reg _414577_414577 ; 
   reg __414577_414577;
   reg _414578_414578 ; 
   reg __414578_414578;
   reg _414579_414579 ; 
   reg __414579_414579;
   reg _414580_414580 ; 
   reg __414580_414580;
   reg _414581_414581 ; 
   reg __414581_414581;
   reg _414582_414582 ; 
   reg __414582_414582;
   reg _414583_414583 ; 
   reg __414583_414583;
   reg _414584_414584 ; 
   reg __414584_414584;
   reg _414585_414585 ; 
   reg __414585_414585;
   reg _414586_414586 ; 
   reg __414586_414586;
   reg _414587_414587 ; 
   reg __414587_414587;
   reg _414588_414588 ; 
   reg __414588_414588;
   reg _414589_414589 ; 
   reg __414589_414589;
   reg _414590_414590 ; 
   reg __414590_414590;
   reg _414591_414591 ; 
   reg __414591_414591;
   reg _414592_414592 ; 
   reg __414592_414592;
   reg _414593_414593 ; 
   reg __414593_414593;
   reg _414594_414594 ; 
   reg __414594_414594;
   reg _414595_414595 ; 
   reg __414595_414595;
   reg _414596_414596 ; 
   reg __414596_414596;
   reg _414597_414597 ; 
   reg __414597_414597;
   reg _414598_414598 ; 
   reg __414598_414598;
   reg _414599_414599 ; 
   reg __414599_414599;
   reg _414600_414600 ; 
   reg __414600_414600;
   reg _414601_414601 ; 
   reg __414601_414601;
   reg _414602_414602 ; 
   reg __414602_414602;
   reg _414603_414603 ; 
   reg __414603_414603;
   reg _414604_414604 ; 
   reg __414604_414604;
   reg _414605_414605 ; 
   reg __414605_414605;
   reg _414606_414606 ; 
   reg __414606_414606;
   reg _414607_414607 ; 
   reg __414607_414607;
   reg _414608_414608 ; 
   reg __414608_414608;
   reg _414609_414609 ; 
   reg __414609_414609;
   reg _414610_414610 ; 
   reg __414610_414610;
   reg _414611_414611 ; 
   reg __414611_414611;
   reg _414612_414612 ; 
   reg __414612_414612;
   reg _414613_414613 ; 
   reg __414613_414613;
   reg _414614_414614 ; 
   reg __414614_414614;
   reg _414615_414615 ; 
   reg __414615_414615;
   reg _414616_414616 ; 
   reg __414616_414616;
   reg _414617_414617 ; 
   reg __414617_414617;
   reg _414618_414618 ; 
   reg __414618_414618;
   reg _414619_414619 ; 
   reg __414619_414619;
   reg _414620_414620 ; 
   reg __414620_414620;
   reg _414621_414621 ; 
   reg __414621_414621;
   reg _414622_414622 ; 
   reg __414622_414622;
   reg _414623_414623 ; 
   reg __414623_414623;
   reg _414624_414624 ; 
   reg __414624_414624;
   reg _414625_414625 ; 
   reg __414625_414625;
   reg _414626_414626 ; 
   reg __414626_414626;
   reg _414627_414627 ; 
   reg __414627_414627;
   reg _414628_414628 ; 
   reg __414628_414628;
   reg _414629_414629 ; 
   reg __414629_414629;
   reg _414630_414630 ; 
   reg __414630_414630;
   reg _414631_414631 ; 
   reg __414631_414631;
   reg _414632_414632 ; 
   reg __414632_414632;
   reg _414633_414633 ; 
   reg __414633_414633;
   reg _414634_414634 ; 
   reg __414634_414634;
   reg _414635_414635 ; 
   reg __414635_414635;
   reg _414636_414636 ; 
   reg __414636_414636;
   reg _414637_414637 ; 
   reg __414637_414637;
   reg _414638_414638 ; 
   reg __414638_414638;
   reg _414639_414639 ; 
   reg __414639_414639;
   reg _414640_414640 ; 
   reg __414640_414640;
   reg _414641_414641 ; 
   reg __414641_414641;
   reg _414642_414642 ; 
   reg __414642_414642;
   reg _414643_414643 ; 
   reg __414643_414643;
   reg _414644_414644 ; 
   reg __414644_414644;
   reg _414645_414645 ; 
   reg __414645_414645;
   reg _414646_414646 ; 
   reg __414646_414646;
   reg _414647_414647 ; 
   reg __414647_414647;
   reg _414648_414648 ; 
   reg __414648_414648;
   reg _414649_414649 ; 
   reg __414649_414649;
   reg _414650_414650 ; 
   reg __414650_414650;
   reg _414651_414651 ; 
   reg __414651_414651;
   reg _414652_414652 ; 
   reg __414652_414652;
   reg _414653_414653 ; 
   reg __414653_414653;
   reg _414654_414654 ; 
   reg __414654_414654;
   reg _414655_414655 ; 
   reg __414655_414655;
   reg _414656_414656 ; 
   reg __414656_414656;
   reg _414657_414657 ; 
   reg __414657_414657;
   reg _414658_414658 ; 
   reg __414658_414658;
   reg _414659_414659 ; 
   reg __414659_414659;
   reg _414660_414660 ; 
   reg __414660_414660;
   reg _414661_414661 ; 
   reg __414661_414661;
   reg _414662_414662 ; 
   reg __414662_414662;
   reg _414663_414663 ; 
   reg __414663_414663;
   reg _414664_414664 ; 
   reg __414664_414664;
   reg _414665_414665 ; 
   reg __414665_414665;
   reg _414666_414666 ; 
   reg __414666_414666;
   reg _414667_414667 ; 
   reg __414667_414667;
   reg _414668_414668 ; 
   reg __414668_414668;
   reg _414669_414669 ; 
   reg __414669_414669;
   reg _414670_414670 ; 
   reg __414670_414670;
   reg _414671_414671 ; 
   reg __414671_414671;
   reg _414672_414672 ; 
   reg __414672_414672;
   reg _414673_414673 ; 
   reg __414673_414673;
   reg _414674_414674 ; 
   reg __414674_414674;
   reg _414675_414675 ; 
   reg __414675_414675;
   reg _414676_414676 ; 
   reg __414676_414676;
   reg _414677_414677 ; 
   reg __414677_414677;
   reg _414678_414678 ; 
   reg __414678_414678;
   reg _414679_414679 ; 
   reg __414679_414679;
   reg _414680_414680 ; 
   reg __414680_414680;
   reg _414681_414681 ; 
   reg __414681_414681;
   reg _414682_414682 ; 
   reg __414682_414682;
   reg _414683_414683 ; 
   reg __414683_414683;
   reg _414684_414684 ; 
   reg __414684_414684;
   reg _414685_414685 ; 
   reg __414685_414685;
   reg _414686_414686 ; 
   reg __414686_414686;
   reg _414687_414687 ; 
   reg __414687_414687;
   reg _414688_414688 ; 
   reg __414688_414688;
   reg _414689_414689 ; 
   reg __414689_414689;
   reg _414690_414690 ; 
   reg __414690_414690;
   reg _414691_414691 ; 
   reg __414691_414691;
   reg _414692_414692 ; 
   reg __414692_414692;
   reg _414693_414693 ; 
   reg __414693_414693;
   reg _414694_414694 ; 
   reg __414694_414694;
   reg _414695_414695 ; 
   reg __414695_414695;
   reg _414696_414696 ; 
   reg __414696_414696;
   reg _414697_414697 ; 
   reg __414697_414697;
   reg _414698_414698 ; 
   reg __414698_414698;
   reg _414699_414699 ; 
   reg __414699_414699;
   reg _414700_414700 ; 
   reg __414700_414700;
   reg _414701_414701 ; 
   reg __414701_414701;
   reg _414702_414702 ; 
   reg __414702_414702;
   reg _414703_414703 ; 
   reg __414703_414703;
   reg _414704_414704 ; 
   reg __414704_414704;
   reg _414705_414705 ; 
   reg __414705_414705;
   reg _414706_414706 ; 
   reg __414706_414706;
   reg _414707_414707 ; 
   reg __414707_414707;
   reg _414708_414708 ; 
   reg __414708_414708;
   reg _414709_414709 ; 
   reg __414709_414709;
   reg _414710_414710 ; 
   reg __414710_414710;
   reg _414711_414711 ; 
   reg __414711_414711;
   reg _414712_414712 ; 
   reg __414712_414712;
   reg _414713_414713 ; 
   reg __414713_414713;
   reg _414714_414714 ; 
   reg __414714_414714;
   reg _414715_414715 ; 
   reg __414715_414715;
   reg _414716_414716 ; 
   reg __414716_414716;
   reg _414717_414717 ; 
   reg __414717_414717;
   reg _414718_414718 ; 
   reg __414718_414718;
   reg _414719_414719 ; 
   reg __414719_414719;
   reg _414720_414720 ; 
   reg __414720_414720;
   reg _414721_414721 ; 
   reg __414721_414721;
   reg _414722_414722 ; 
   reg __414722_414722;
   reg _414723_414723 ; 
   reg __414723_414723;
   reg _414724_414724 ; 
   reg __414724_414724;
   reg _414725_414725 ; 
   reg __414725_414725;
   reg _414726_414726 ; 
   reg __414726_414726;
   reg _414727_414727 ; 
   reg __414727_414727;
   reg _414728_414728 ; 
   reg __414728_414728;
   reg _414729_414729 ; 
   reg __414729_414729;
   reg _414730_414730 ; 
   reg __414730_414730;
   reg _414731_414731 ; 
   reg __414731_414731;
   reg _414732_414732 ; 
   reg __414732_414732;
   reg _414733_414733 ; 
   reg __414733_414733;
   reg _414734_414734 ; 
   reg __414734_414734;
   reg _414735_414735 ; 
   reg __414735_414735;
   reg _414736_414736 ; 
   reg __414736_414736;
   reg _414737_414737 ; 
   reg __414737_414737;
   reg _414738_414738 ; 
   reg __414738_414738;
   reg _414739_414739 ; 
   reg __414739_414739;
   reg _414740_414740 ; 
   reg __414740_414740;
   reg _414741_414741 ; 
   reg __414741_414741;
   reg _414742_414742 ; 
   reg __414742_414742;
   reg _414743_414743 ; 
   reg __414743_414743;
   reg _414744_414744 ; 
   reg __414744_414744;
   reg _414745_414745 ; 
   reg __414745_414745;
   reg _414746_414746 ; 
   reg __414746_414746;
   reg _414747_414747 ; 
   reg __414747_414747;
   reg _414748_414748 ; 
   reg __414748_414748;
   reg _414749_414749 ; 
   reg __414749_414749;
   reg _414750_414750 ; 
   reg __414750_414750;
   reg _414751_414751 ; 
   reg __414751_414751;
   reg _414752_414752 ; 
   reg __414752_414752;
   reg _414753_414753 ; 
   reg __414753_414753;
   reg _414754_414754 ; 
   reg __414754_414754;
   reg _414755_414755 ; 
   reg __414755_414755;
   reg _414756_414756 ; 
   reg __414756_414756;
   reg _414757_414757 ; 
   reg __414757_414757;
   reg _414758_414758 ; 
   reg __414758_414758;
   reg _414759_414759 ; 
   reg __414759_414759;
   reg _414760_414760 ; 
   reg __414760_414760;
   reg _414761_414761 ; 
   reg __414761_414761;
   reg _414762_414762 ; 
   reg __414762_414762;
   reg _414763_414763 ; 
   reg __414763_414763;
   reg _414764_414764 ; 
   reg __414764_414764;
   reg _414765_414765 ; 
   reg __414765_414765;
   reg _414766_414766 ; 
   reg __414766_414766;
   reg _414767_414767 ; 
   reg __414767_414767;
   reg _414768_414768 ; 
   reg __414768_414768;
   reg _414769_414769 ; 
   reg __414769_414769;
   reg _414770_414770 ; 
   reg __414770_414770;
   reg _414771_414771 ; 
   reg __414771_414771;
   reg _414772_414772 ; 
   reg __414772_414772;
   reg _414773_414773 ; 
   reg __414773_414773;
   reg _414774_414774 ; 
   reg __414774_414774;
   reg _414775_414775 ; 
   reg __414775_414775;
   reg _414776_414776 ; 
   reg __414776_414776;
   reg _414777_414777 ; 
   reg __414777_414777;
   reg _414778_414778 ; 
   reg __414778_414778;
   reg _414779_414779 ; 
   reg __414779_414779;
   reg _414780_414780 ; 
   reg __414780_414780;
   reg _414781_414781 ; 
   reg __414781_414781;
   reg _414782_414782 ; 
   reg __414782_414782;
   reg _414783_414783 ; 
   reg __414783_414783;
   reg _414784_414784 ; 
   reg __414784_414784;
   reg _414785_414785 ; 
   reg __414785_414785;
   reg _414786_414786 ; 
   reg __414786_414786;
   reg _414787_414787 ; 
   reg __414787_414787;
   reg _414788_414788 ; 
   reg __414788_414788;
   reg _414789_414789 ; 
   reg __414789_414789;
   reg _414790_414790 ; 
   reg __414790_414790;
   reg _414791_414791 ; 
   reg __414791_414791;
   reg _414792_414792 ; 
   reg __414792_414792;
   reg _414793_414793 ; 
   reg __414793_414793;
   reg _414794_414794 ; 
   reg __414794_414794;
   reg _414795_414795 ; 
   reg __414795_414795;
   reg _414796_414796 ; 
   reg __414796_414796;
   reg _414797_414797 ; 
   reg __414797_414797;
   reg _414798_414798 ; 
   reg __414798_414798;
   reg _414799_414799 ; 
   reg __414799_414799;
   reg _414800_414800 ; 
   reg __414800_414800;
   reg _414801_414801 ; 
   reg __414801_414801;
   reg _414802_414802 ; 
   reg __414802_414802;
   reg _414803_414803 ; 
   reg __414803_414803;
   reg _414804_414804 ; 
   reg __414804_414804;
   reg _414805_414805 ; 
   reg __414805_414805;
   reg _414806_414806 ; 
   reg __414806_414806;
   reg _414807_414807 ; 
   reg __414807_414807;
   reg _414808_414808 ; 
   reg __414808_414808;
   reg _414809_414809 ; 
   reg __414809_414809;
   reg _414810_414810 ; 
   reg __414810_414810;
   reg _414811_414811 ; 
   reg __414811_414811;
   reg _414812_414812 ; 
   reg __414812_414812;
   reg _414813_414813 ; 
   reg __414813_414813;
   reg _414814_414814 ; 
   reg __414814_414814;
   reg _414815_414815 ; 
   reg __414815_414815;
   reg _414816_414816 ; 
   reg __414816_414816;
   reg _414817_414817 ; 
   reg __414817_414817;
   reg _414818_414818 ; 
   reg __414818_414818;
   reg _414819_414819 ; 
   reg __414819_414819;
   reg _414820_414820 ; 
   reg __414820_414820;
   reg _414821_414821 ; 
   reg __414821_414821;
   reg _414822_414822 ; 
   reg __414822_414822;
   reg _414823_414823 ; 
   reg __414823_414823;
   reg _414824_414824 ; 
   reg __414824_414824;
   reg _414825_414825 ; 
   reg __414825_414825;
   reg _414826_414826 ; 
   reg __414826_414826;
   reg _414827_414827 ; 
   reg __414827_414827;
   reg _414828_414828 ; 
   reg __414828_414828;
   reg _414829_414829 ; 
   reg __414829_414829;
   reg _414830_414830 ; 
   reg __414830_414830;
   reg _414831_414831 ; 
   reg __414831_414831;
   reg _414832_414832 ; 
   reg __414832_414832;
   reg _414833_414833 ; 
   reg __414833_414833;
   reg _414834_414834 ; 
   reg __414834_414834;
   reg _414835_414835 ; 
   reg __414835_414835;
   reg _414836_414836 ; 
   reg __414836_414836;
   reg _414837_414837 ; 
   reg __414837_414837;
   reg _414838_414838 ; 
   reg __414838_414838;
   reg _414839_414839 ; 
   reg __414839_414839;
   reg _414840_414840 ; 
   reg __414840_414840;
   reg _414841_414841 ; 
   reg __414841_414841;
   reg _414842_414842 ; 
   reg __414842_414842;
   reg _414843_414843 ; 
   reg __414843_414843;
   reg _414844_414844 ; 
   reg __414844_414844;
   reg _414845_414845 ; 
   reg __414845_414845;
   reg _414846_414846 ; 
   reg __414846_414846;
   reg _414847_414847 ; 
   reg __414847_414847;
   reg _414848_414848 ; 
   reg __414848_414848;
   reg _414849_414849 ; 
   reg __414849_414849;
   reg _414850_414850 ; 
   reg __414850_414850;
   reg _414851_414851 ; 
   reg __414851_414851;
   reg _414852_414852 ; 
   reg __414852_414852;
   reg _414853_414853 ; 
   reg __414853_414853;
   reg _414854_414854 ; 
   reg __414854_414854;
   reg _414855_414855 ; 
   reg __414855_414855;
   reg _414856_414856 ; 
   reg __414856_414856;
   reg _414857_414857 ; 
   reg __414857_414857;
   reg _414858_414858 ; 
   reg __414858_414858;
   reg _414859_414859 ; 
   reg __414859_414859;
   reg _414860_414860 ; 
   reg __414860_414860;
   reg _414861_414861 ; 
   reg __414861_414861;
   reg _414862_414862 ; 
   reg __414862_414862;
   reg _414863_414863 ; 
   reg __414863_414863;
   reg _414864_414864 ; 
   reg __414864_414864;
   reg _414865_414865 ; 
   reg __414865_414865;
   reg _414866_414866 ; 
   reg __414866_414866;
   reg _414867_414867 ; 
   reg __414867_414867;
   reg _414868_414868 ; 
   reg __414868_414868;
   reg _414869_414869 ; 
   reg __414869_414869;
   reg _414870_414870 ; 
   reg __414870_414870;
   reg _414871_414871 ; 
   reg __414871_414871;
   reg _414872_414872 ; 
   reg __414872_414872;
   reg _414873_414873 ; 
   reg __414873_414873;
   reg _414874_414874 ; 
   reg __414874_414874;
   reg _414875_414875 ; 
   reg __414875_414875;
   reg _414876_414876 ; 
   reg __414876_414876;
   reg _414877_414877 ; 
   reg __414877_414877;
   reg _414878_414878 ; 
   reg __414878_414878;
   reg _414879_414879 ; 
   reg __414879_414879;
   reg _414880_414880 ; 
   reg __414880_414880;
   reg _414881_414881 ; 
   reg __414881_414881;
   reg _414882_414882 ; 
   reg __414882_414882;
   reg _414883_414883 ; 
   reg __414883_414883;
   reg _414884_414884 ; 
   reg __414884_414884;
   reg _414885_414885 ; 
   reg __414885_414885;
   reg _414886_414886 ; 
   reg __414886_414886;
   reg _414887_414887 ; 
   reg __414887_414887;
   reg _414888_414888 ; 
   reg __414888_414888;
   reg _414889_414889 ; 
   reg __414889_414889;
   reg _414890_414890 ; 
   reg __414890_414890;
   reg _414891_414891 ; 
   reg __414891_414891;
   reg _414892_414892 ; 
   reg __414892_414892;
   reg _414893_414893 ; 
   reg __414893_414893;
   reg _414894_414894 ; 
   reg __414894_414894;
   reg _414895_414895 ; 
   reg __414895_414895;
   reg _414896_414896 ; 
   reg __414896_414896;
   reg _414897_414897 ; 
   reg __414897_414897;
   reg _414898_414898 ; 
   reg __414898_414898;
   reg _414899_414899 ; 
   reg __414899_414899;
   reg _414900_414900 ; 
   reg __414900_414900;
   reg _414901_414901 ; 
   reg __414901_414901;
   reg _414902_414902 ; 
   reg __414902_414902;
   reg _414903_414903 ; 
   reg __414903_414903;
   reg _414904_414904 ; 
   reg __414904_414904;
   reg _414905_414905 ; 
   reg __414905_414905;
   reg _414906_414906 ; 
   reg __414906_414906;
   reg _414907_414907 ; 
   reg __414907_414907;
   reg _414908_414908 ; 
   reg __414908_414908;
   reg _414909_414909 ; 
   reg __414909_414909;
   reg _414910_414910 ; 
   reg __414910_414910;
   reg _414911_414911 ; 
   reg __414911_414911;
   reg _414912_414912 ; 
   reg __414912_414912;
   reg _414913_414913 ; 
   reg __414913_414913;
   reg _414914_414914 ; 
   reg __414914_414914;
   reg _414915_414915 ; 
   reg __414915_414915;
   reg _414916_414916 ; 
   reg __414916_414916;
   reg _414917_414917 ; 
   reg __414917_414917;
   reg _414918_414918 ; 
   reg __414918_414918;
   reg _414919_414919 ; 
   reg __414919_414919;
   reg _414920_414920 ; 
   reg __414920_414920;
   reg _414921_414921 ; 
   reg __414921_414921;
   reg _414922_414922 ; 
   reg __414922_414922;
   reg _414923_414923 ; 
   reg __414923_414923;
   reg _414924_414924 ; 
   reg __414924_414924;
   reg _414925_414925 ; 
   reg __414925_414925;
   reg _414926_414926 ; 
   reg __414926_414926;
   reg _414927_414927 ; 
   reg __414927_414927;
   reg _414928_414928 ; 
   reg __414928_414928;
   reg _414929_414929 ; 
   reg __414929_414929;
   reg _414930_414930 ; 
   reg __414930_414930;
   reg _414931_414931 ; 
   reg __414931_414931;
   reg _414932_414932 ; 
   reg __414932_414932;
   reg _414933_414933 ; 
   reg __414933_414933;
   reg _414934_414934 ; 
   reg __414934_414934;
   reg _414935_414935 ; 
   reg __414935_414935;
   reg _414936_414936 ; 
   reg __414936_414936;
   reg _414937_414937 ; 
   reg __414937_414937;
   reg _414938_414938 ; 
   reg __414938_414938;
   reg _414939_414939 ; 
   reg __414939_414939;
   reg _414940_414940 ; 
   reg __414940_414940;
   reg _414941_414941 ; 
   reg __414941_414941;
   reg _414942_414942 ; 
   reg __414942_414942;
   reg _414943_414943 ; 
   reg __414943_414943;
   reg _414944_414944 ; 
   reg __414944_414944;
   reg _414945_414945 ; 
   reg __414945_414945;
   reg _414946_414946 ; 
   reg __414946_414946;
   reg _414947_414947 ; 
   reg __414947_414947;
   reg _414948_414948 ; 
   reg __414948_414948;
   reg _414949_414949 ; 
   reg __414949_414949;
   reg _414950_414950 ; 
   reg __414950_414950;
   reg _414951_414951 ; 
   reg __414951_414951;
   reg _414952_414952 ; 
   reg __414952_414952;
   reg _414953_414953 ; 
   reg __414953_414953;
   reg _414954_414954 ; 
   reg __414954_414954;
   reg _414955_414955 ; 
   reg __414955_414955;
   reg _414956_414956 ; 
   reg __414956_414956;
   reg _414957_414957 ; 
   reg __414957_414957;
   reg _414958_414958 ; 
   reg __414958_414958;
   reg _414959_414959 ; 
   reg __414959_414959;
   reg _414960_414960 ; 
   reg __414960_414960;
   reg _414961_414961 ; 
   reg __414961_414961;
   reg _414962_414962 ; 
   reg __414962_414962;
   reg _414963_414963 ; 
   reg __414963_414963;
   reg _414964_414964 ; 
   reg __414964_414964;
   reg _414965_414965 ; 
   reg __414965_414965;
   reg _414966_414966 ; 
   reg __414966_414966;
   reg _414967_414967 ; 
   reg __414967_414967;
   reg _414968_414968 ; 
   reg __414968_414968;
   reg _414969_414969 ; 
   reg __414969_414969;
   reg _414970_414970 ; 
   reg __414970_414970;
   reg _414971_414971 ; 
   reg __414971_414971;
   reg _414972_414972 ; 
   reg __414972_414972;
   reg _414973_414973 ; 
   reg __414973_414973;
   reg _414974_414974 ; 
   reg __414974_414974;
   reg _414975_414975 ; 
   reg __414975_414975;
   reg _414976_414976 ; 
   reg __414976_414976;
   reg _414977_414977 ; 
   reg __414977_414977;
   reg _414978_414978 ; 
   reg __414978_414978;
   reg _414979_414979 ; 
   reg __414979_414979;
   reg _414980_414980 ; 
   reg __414980_414980;
   reg _414981_414981 ; 
   reg __414981_414981;
   reg _414982_414982 ; 
   reg __414982_414982;
   reg _414983_414983 ; 
   reg __414983_414983;
   reg _414984_414984 ; 
   reg __414984_414984;
   reg _414985_414985 ; 
   reg __414985_414985;
   reg _414986_414986 ; 
   reg __414986_414986;
   reg _414987_414987 ; 
   reg __414987_414987;
   reg _414988_414988 ; 
   reg __414988_414988;
   reg _414989_414989 ; 
   reg __414989_414989;
   reg _414990_414990 ; 
   reg __414990_414990;
   reg _414991_414991 ; 
   reg __414991_414991;
   reg _414992_414992 ; 
   reg __414992_414992;
   reg _414993_414993 ; 
   reg __414993_414993;
   reg _414994_414994 ; 
   reg __414994_414994;
   reg _414995_414995 ; 
   reg __414995_414995;
   reg _414996_414996 ; 
   reg __414996_414996;
   reg _414997_414997 ; 
   reg __414997_414997;
   reg _414998_414998 ; 
   reg __414998_414998;
   reg _414999_414999 ; 
   reg __414999_414999;
   reg _415000_415000 ; 
   reg __415000_415000;
   reg _415001_415001 ; 
   reg __415001_415001;
   reg _415002_415002 ; 
   reg __415002_415002;
   reg _415003_415003 ; 
   reg __415003_415003;
   reg _415004_415004 ; 
   reg __415004_415004;
   reg _415005_415005 ; 
   reg __415005_415005;
   reg _415006_415006 ; 
   reg __415006_415006;
   reg _415007_415007 ; 
   reg __415007_415007;
   reg _415008_415008 ; 
   reg __415008_415008;
   reg _415009_415009 ; 
   reg __415009_415009;
   reg _415010_415010 ; 
   reg __415010_415010;
   reg _415011_415011 ; 
   reg __415011_415011;
   reg _415012_415012 ; 
   reg __415012_415012;
   reg _415013_415013 ; 
   reg __415013_415013;
   reg _415014_415014 ; 
   reg __415014_415014;
   reg _415015_415015 ; 
   reg __415015_415015;
   reg _415016_415016 ; 
   reg __415016_415016;
   reg _415017_415017 ; 
   reg __415017_415017;
   reg _415018_415018 ; 
   reg __415018_415018;
   reg _415019_415019 ; 
   reg __415019_415019;
   reg _415020_415020 ; 
   reg __415020_415020;
   reg _415021_415021 ; 
   reg __415021_415021;
   reg _415022_415022 ; 
   reg __415022_415022;
   reg _415023_415023 ; 
   reg __415023_415023;
   reg _415024_415024 ; 
   reg __415024_415024;
   reg _415025_415025 ; 
   reg __415025_415025;
   reg _415026_415026 ; 
   reg __415026_415026;
   reg _415027_415027 ; 
   reg __415027_415027;
   reg _415028_415028 ; 
   reg __415028_415028;
   reg _415029_415029 ; 
   reg __415029_415029;
   reg _415030_415030 ; 
   reg __415030_415030;
   reg _415031_415031 ; 
   reg __415031_415031;
   reg _415032_415032 ; 
   reg __415032_415032;
   reg _415033_415033 ; 
   reg __415033_415033;
   reg _415034_415034 ; 
   reg __415034_415034;
   reg _415035_415035 ; 
   reg __415035_415035;
   reg _415036_415036 ; 
   reg __415036_415036;
   reg _415037_415037 ; 
   reg __415037_415037;
   reg _415038_415038 ; 
   reg __415038_415038;
   reg _415039_415039 ; 
   reg __415039_415039;
   reg _415040_415040 ; 
   reg __415040_415040;
   reg _415041_415041 ; 
   reg __415041_415041;
   reg _415042_415042 ; 
   reg __415042_415042;
   reg _415043_415043 ; 
   reg __415043_415043;
   reg _415044_415044 ; 
   reg __415044_415044;
   reg _415045_415045 ; 
   reg __415045_415045;
   reg _415046_415046 ; 
   reg __415046_415046;
   reg _415047_415047 ; 
   reg __415047_415047;
   reg _415048_415048 ; 
   reg __415048_415048;
   reg _415049_415049 ; 
   reg __415049_415049;
   reg _415050_415050 ; 
   reg __415050_415050;
   reg _415051_415051 ; 
   reg __415051_415051;
   reg _415052_415052 ; 
   reg __415052_415052;
   reg _415053_415053 ; 
   reg __415053_415053;
   reg _415054_415054 ; 
   reg __415054_415054;
   reg _415055_415055 ; 
   reg __415055_415055;
   reg _415056_415056 ; 
   reg __415056_415056;
   reg _415057_415057 ; 
   reg __415057_415057;
   reg _415058_415058 ; 
   reg __415058_415058;
   reg _415059_415059 ; 
   reg __415059_415059;
   reg _415060_415060 ; 
   reg __415060_415060;
   reg _415061_415061 ; 
   reg __415061_415061;
   reg _415062_415062 ; 
   reg __415062_415062;
   reg _415063_415063 ; 
   reg __415063_415063;
   reg _415064_415064 ; 
   reg __415064_415064;
   reg _415065_415065 ; 
   reg __415065_415065;
   reg _415066_415066 ; 
   reg __415066_415066;
   reg _415067_415067 ; 
   reg __415067_415067;
   reg _415068_415068 ; 
   reg __415068_415068;
   reg _415069_415069 ; 
   reg __415069_415069;
   reg _415070_415070 ; 
   reg __415070_415070;
   reg _415071_415071 ; 
   reg __415071_415071;
   reg _415072_415072 ; 
   reg __415072_415072;
   reg _415073_415073 ; 
   reg __415073_415073;
   reg _415074_415074 ; 
   reg __415074_415074;
   reg _415075_415075 ; 
   reg __415075_415075;
   reg _415076_415076 ; 
   reg __415076_415076;
   reg _415077_415077 ; 
   reg __415077_415077;
   reg _415078_415078 ; 
   reg __415078_415078;
   reg _415079_415079 ; 
   reg __415079_415079;
   reg _415080_415080 ; 
   reg __415080_415080;
   reg _415081_415081 ; 
   reg __415081_415081;
   reg _415082_415082 ; 
   reg __415082_415082;
   reg _415083_415083 ; 
   reg __415083_415083;
   reg _415084_415084 ; 
   reg __415084_415084;
   reg _415085_415085 ; 
   reg __415085_415085;
   reg _415086_415086 ; 
   reg __415086_415086;
   reg _415087_415087 ; 
   reg __415087_415087;
   reg _415088_415088 ; 
   reg __415088_415088;
   reg _415089_415089 ; 
   reg __415089_415089;
   reg _415090_415090 ; 
   reg __415090_415090;
   reg _415091_415091 ; 
   reg __415091_415091;
   reg _415092_415092 ; 
   reg __415092_415092;
   reg _415093_415093 ; 
   reg __415093_415093;
   reg _415094_415094 ; 
   reg __415094_415094;
   reg _415095_415095 ; 
   reg __415095_415095;
   reg _415096_415096 ; 
   reg __415096_415096;
   reg _415097_415097 ; 
   reg __415097_415097;
   reg _415098_415098 ; 
   reg __415098_415098;
   reg _415099_415099 ; 
   reg __415099_415099;
   reg _415100_415100 ; 
   reg __415100_415100;
   reg _415101_415101 ; 
   reg __415101_415101;
   reg _415102_415102 ; 
   reg __415102_415102;
   reg _415103_415103 ; 
   reg __415103_415103;
   reg _415104_415104 ; 
   reg __415104_415104;
   reg _415105_415105 ; 
   reg __415105_415105;
   reg _415106_415106 ; 
   reg __415106_415106;
   reg _415107_415107 ; 
   reg __415107_415107;
   reg _415108_415108 ; 
   reg __415108_415108;
   reg _415109_415109 ; 
   reg __415109_415109;
   reg _415110_415110 ; 
   reg __415110_415110;
   reg _415111_415111 ; 
   reg __415111_415111;
   reg _415112_415112 ; 
   reg __415112_415112;
   reg _415113_415113 ; 
   reg __415113_415113;
   reg _415114_415114 ; 
   reg __415114_415114;
   reg _415115_415115 ; 
   reg __415115_415115;
   reg _415116_415116 ; 
   reg __415116_415116;
   reg _415117_415117 ; 
   reg __415117_415117;
   reg _415118_415118 ; 
   reg __415118_415118;
   reg _415119_415119 ; 
   reg __415119_415119;
   reg _415120_415120 ; 
   reg __415120_415120;
   reg _415121_415121 ; 
   reg __415121_415121;
   reg _415122_415122 ; 
   reg __415122_415122;
   reg _415123_415123 ; 
   reg __415123_415123;
   reg _415124_415124 ; 
   reg __415124_415124;
   reg _415125_415125 ; 
   reg __415125_415125;
   reg _415126_415126 ; 
   reg __415126_415126;
   reg _415127_415127 ; 
   reg __415127_415127;
   reg _415128_415128 ; 
   reg __415128_415128;
   reg _415129_415129 ; 
   reg __415129_415129;
   reg _415130_415130 ; 
   reg __415130_415130;
   reg _415131_415131 ; 
   reg __415131_415131;
   reg _415132_415132 ; 
   reg __415132_415132;
   reg _415133_415133 ; 
   reg __415133_415133;
   reg _415134_415134 ; 
   reg __415134_415134;
   reg _415135_415135 ; 
   reg __415135_415135;
   reg _415136_415136 ; 
   reg __415136_415136;
   reg _415137_415137 ; 
   reg __415137_415137;
   reg _415138_415138 ; 
   reg __415138_415138;
   reg _415139_415139 ; 
   reg __415139_415139;
   reg _415140_415140 ; 
   reg __415140_415140;
   reg _415141_415141 ; 
   reg __415141_415141;
   reg _415142_415142 ; 
   reg __415142_415142;
   reg _415143_415143 ; 
   reg __415143_415143;
   reg _415144_415144 ; 
   reg __415144_415144;
   reg _415145_415145 ; 
   reg __415145_415145;
   reg _415146_415146 ; 
   reg __415146_415146;
   reg _415147_415147 ; 
   reg __415147_415147;
   reg _415148_415148 ; 
   reg __415148_415148;
   reg _415149_415149 ; 
   reg __415149_415149;
   reg _415150_415150 ; 
   reg __415150_415150;
   reg _415151_415151 ; 
   reg __415151_415151;
   reg _415152_415152 ; 
   reg __415152_415152;
   reg _415153_415153 ; 
   reg __415153_415153;
   reg _415154_415154 ; 
   reg __415154_415154;
   reg _415155_415155 ; 
   reg __415155_415155;
   reg _415156_415156 ; 
   reg __415156_415156;
   reg _415157_415157 ; 
   reg __415157_415157;
   reg _415158_415158 ; 
   reg __415158_415158;
   reg _415159_415159 ; 
   reg __415159_415159;
   reg _415160_415160 ; 
   reg __415160_415160;
   reg _415161_415161 ; 
   reg __415161_415161;
   reg _415162_415162 ; 
   reg __415162_415162;
   reg _415163_415163 ; 
   reg __415163_415163;
   reg _415164_415164 ; 
   reg __415164_415164;
   reg _415165_415165 ; 
   reg __415165_415165;
   reg _415166_415166 ; 
   reg __415166_415166;
   reg _415167_415167 ; 
   reg __415167_415167;
   reg _415168_415168 ; 
   reg __415168_415168;
   reg _415169_415169 ; 
   reg __415169_415169;
   reg _415170_415170 ; 
   reg __415170_415170;
   reg _415171_415171 ; 
   reg __415171_415171;
   reg _415172_415172 ; 
   reg __415172_415172;
   reg _415173_415173 ; 
   reg __415173_415173;
   reg _415174_415174 ; 
   reg __415174_415174;
   reg _415175_415175 ; 
   reg __415175_415175;
   reg _415176_415176 ; 
   reg __415176_415176;
   reg _415177_415177 ; 
   reg __415177_415177;
   reg _415178_415178 ; 
   reg __415178_415178;
   reg _415179_415179 ; 
   reg __415179_415179;
   reg _415180_415180 ; 
   reg __415180_415180;
   reg _415181_415181 ; 
   reg __415181_415181;
   reg _415182_415182 ; 
   reg __415182_415182;
   reg _415183_415183 ; 
   reg __415183_415183;
   reg _415184_415184 ; 
   reg __415184_415184;
   reg _415185_415185 ; 
   reg __415185_415185;
   reg _415186_415186 ; 
   reg __415186_415186;
   reg _415187_415187 ; 
   reg __415187_415187;
   reg _415188_415188 ; 
   reg __415188_415188;
   reg _415189_415189 ; 
   reg __415189_415189;
   reg _415190_415190 ; 
   reg __415190_415190;
   reg _415191_415191 ; 
   reg __415191_415191;
   reg _415192_415192 ; 
   reg __415192_415192;
   reg _415193_415193 ; 
   reg __415193_415193;
   reg _415194_415194 ; 
   reg __415194_415194;
   reg _415195_415195 ; 
   reg __415195_415195;
   reg _415196_415196 ; 
   reg __415196_415196;
   reg _415197_415197 ; 
   reg __415197_415197;
   reg _415198_415198 ; 
   reg __415198_415198;
   reg _415199_415199 ; 
   reg __415199_415199;
   reg _415200_415200 ; 
   reg __415200_415200;
   reg _415201_415201 ; 
   reg __415201_415201;
   reg _415202_415202 ; 
   reg __415202_415202;
   reg _415203_415203 ; 
   reg __415203_415203;
   reg _415204_415204 ; 
   reg __415204_415204;
   reg _415205_415205 ; 
   reg __415205_415205;
   reg _415206_415206 ; 
   reg __415206_415206;
   reg _415207_415207 ; 
   reg __415207_415207;
   reg _415208_415208 ; 
   reg __415208_415208;
   reg _415209_415209 ; 
   reg __415209_415209;
   reg _415210_415210 ; 
   reg __415210_415210;
   reg _415211_415211 ; 
   reg __415211_415211;
   reg _415212_415212 ; 
   reg __415212_415212;
   reg _415213_415213 ; 
   reg __415213_415213;
   reg _415214_415214 ; 
   reg __415214_415214;
   reg _415215_415215 ; 
   reg __415215_415215;
   reg _415216_415216 ; 
   reg __415216_415216;
   reg _415217_415217 ; 
   reg __415217_415217;
   reg _415218_415218 ; 
   reg __415218_415218;
   reg _415219_415219 ; 
   reg __415219_415219;
   reg _415220_415220 ; 
   reg __415220_415220;
   reg _415221_415221 ; 
   reg __415221_415221;
   reg _415222_415222 ; 
   reg __415222_415222;
   reg _415223_415223 ; 
   reg __415223_415223;
   reg _415224_415224 ; 
   reg __415224_415224;
   reg _415225_415225 ; 
   reg __415225_415225;
   reg _415226_415226 ; 
   reg __415226_415226;
   reg _415227_415227 ; 
   reg __415227_415227;
   reg _415228_415228 ; 
   reg __415228_415228;
   reg _415229_415229 ; 
   reg __415229_415229;
   reg _415230_415230 ; 
   reg __415230_415230;
   reg _415231_415231 ; 
   reg __415231_415231;
   reg _415232_415232 ; 
   reg __415232_415232;
   reg _415233_415233 ; 
   reg __415233_415233;
   reg _415234_415234 ; 
   reg __415234_415234;
   reg _415235_415235 ; 
   reg __415235_415235;
   reg _415236_415236 ; 
   reg __415236_415236;
   reg _415237_415237 ; 
   reg __415237_415237;
   reg _415238_415238 ; 
   reg __415238_415238;
   reg _415239_415239 ; 
   reg __415239_415239;
   reg _415240_415240 ; 
   reg __415240_415240;
   reg _415241_415241 ; 
   reg __415241_415241;
   reg _415242_415242 ; 
   reg __415242_415242;
   reg _415243_415243 ; 
   reg __415243_415243;
   reg _415244_415244 ; 
   reg __415244_415244;
   reg _415245_415245 ; 
   reg __415245_415245;
   reg _415246_415246 ; 
   reg __415246_415246;
   reg _415247_415247 ; 
   reg __415247_415247;
   reg _415248_415248 ; 
   reg __415248_415248;
   reg _415249_415249 ; 
   reg __415249_415249;
   reg _415250_415250 ; 
   reg __415250_415250;
   reg _415251_415251 ; 
   reg __415251_415251;
   reg _415252_415252 ; 
   reg __415252_415252;
   reg _415253_415253 ; 
   reg __415253_415253;
   reg _415254_415254 ; 
   reg __415254_415254;
   reg _415255_415255 ; 
   reg __415255_415255;
   reg _415256_415256 ; 
   reg __415256_415256;
   reg _415257_415257 ; 
   reg __415257_415257;
   reg _415258_415258 ; 
   reg __415258_415258;
   reg _415259_415259 ; 
   reg __415259_415259;
   reg _415260_415260 ; 
   reg __415260_415260;
   reg _415261_415261 ; 
   reg __415261_415261;
   reg _415262_415262 ; 
   reg __415262_415262;
   reg _415263_415263 ; 
   reg __415263_415263;
   reg _415264_415264 ; 
   reg __415264_415264;
   reg _415265_415265 ; 
   reg __415265_415265;
   reg _415266_415266 ; 
   reg __415266_415266;
   reg _415267_415267 ; 
   reg __415267_415267;
   reg _415268_415268 ; 
   reg __415268_415268;
   reg _415269_415269 ; 
   reg __415269_415269;
   reg _415270_415270 ; 
   reg __415270_415270;
   reg _415271_415271 ; 
   reg __415271_415271;
   reg _415272_415272 ; 
   reg __415272_415272;
   reg _415273_415273 ; 
   reg __415273_415273;
   reg _415274_415274 ; 
   reg __415274_415274;
   reg _415275_415275 ; 
   reg __415275_415275;
   reg _415276_415276 ; 
   reg __415276_415276;
   reg _415277_415277 ; 
   reg __415277_415277;
   reg _415278_415278 ; 
   reg __415278_415278;
   reg _415279_415279 ; 
   reg __415279_415279;
   reg _415280_415280 ; 
   reg __415280_415280;
   reg _415281_415281 ; 
   reg __415281_415281;
   reg _415282_415282 ; 
   reg __415282_415282;
   reg _415283_415283 ; 
   reg __415283_415283;
   reg _415284_415284 ; 
   reg __415284_415284;
   reg _415285_415285 ; 
   reg __415285_415285;
   reg _415286_415286 ; 
   reg __415286_415286;
   reg _415287_415287 ; 
   reg __415287_415287;
   reg _415288_415288 ; 
   reg __415288_415288;
   reg _415289_415289 ; 
   reg __415289_415289;
   reg _415290_415290 ; 
   reg __415290_415290;
   reg _415291_415291 ; 
   reg __415291_415291;
   reg _415292_415292 ; 
   reg __415292_415292;
   reg _415293_415293 ; 
   reg __415293_415293;
   reg _415294_415294 ; 
   reg __415294_415294;
   reg _415295_415295 ; 
   reg __415295_415295;
   reg _415296_415296 ; 
   reg __415296_415296;
   reg _415297_415297 ; 
   reg __415297_415297;
   reg _415298_415298 ; 
   reg __415298_415298;
   reg _415299_415299 ; 
   reg __415299_415299;
   reg _415300_415300 ; 
   reg __415300_415300;
   reg _415301_415301 ; 
   reg __415301_415301;
   reg _415302_415302 ; 
   reg __415302_415302;
   reg _415303_415303 ; 
   reg __415303_415303;
   reg _415304_415304 ; 
   reg __415304_415304;
   reg _415305_415305 ; 
   reg __415305_415305;
   reg _415306_415306 ; 
   reg __415306_415306;
   reg _415307_415307 ; 
   reg __415307_415307;
   reg _415308_415308 ; 
   reg __415308_415308;
   reg _415309_415309 ; 
   reg __415309_415309;
   reg _415310_415310 ; 
   reg __415310_415310;
   reg _415311_415311 ; 
   reg __415311_415311;
   reg _415312_415312 ; 
   reg __415312_415312;
   reg _415313_415313 ; 
   reg __415313_415313;
   reg _415314_415314 ; 
   reg __415314_415314;
   reg _415315_415315 ; 
   reg __415315_415315;
   reg _415316_415316 ; 
   reg __415316_415316;
   reg _415317_415317 ; 
   reg __415317_415317;
   reg _415318_415318 ; 
   reg __415318_415318;
   reg _415319_415319 ; 
   reg __415319_415319;
   reg _415320_415320 ; 
   reg __415320_415320;
   reg _415321_415321 ; 
   reg __415321_415321;
   reg _415322_415322 ; 
   reg __415322_415322;
   reg _415323_415323 ; 
   reg __415323_415323;
   reg _415324_415324 ; 
   reg __415324_415324;
   reg _415325_415325 ; 
   reg __415325_415325;
   reg _415326_415326 ; 
   reg __415326_415326;
   reg _415327_415327 ; 
   reg __415327_415327;
   reg _415328_415328 ; 
   reg __415328_415328;
   reg _415329_415329 ; 
   reg __415329_415329;
   reg _415330_415330 ; 
   reg __415330_415330;
   reg _415331_415331 ; 
   reg __415331_415331;
   reg _415332_415332 ; 
   reg __415332_415332;
   reg _415333_415333 ; 
   reg __415333_415333;
   reg _415334_415334 ; 
   reg __415334_415334;
   reg _415335_415335 ; 
   reg __415335_415335;
   reg _415336_415336 ; 
   reg __415336_415336;
   reg _415337_415337 ; 
   reg __415337_415337;
   reg _415338_415338 ; 
   reg __415338_415338;
   reg _415339_415339 ; 
   reg __415339_415339;
   reg _415340_415340 ; 
   reg __415340_415340;
   reg _415341_415341 ; 
   reg __415341_415341;
   reg _415342_415342 ; 
   reg __415342_415342;
   reg _415343_415343 ; 
   reg __415343_415343;
   reg _415344_415344 ; 
   reg __415344_415344;
   reg _415345_415345 ; 
   reg __415345_415345;
   reg _415346_415346 ; 
   reg __415346_415346;
   reg _415347_415347 ; 
   reg __415347_415347;
   reg _415348_415348 ; 
   reg __415348_415348;
   reg _415349_415349 ; 
   reg __415349_415349;
   reg _415350_415350 ; 
   reg __415350_415350;
   reg _415351_415351 ; 
   reg __415351_415351;
   reg _415352_415352 ; 
   reg __415352_415352;
   reg _415353_415353 ; 
   reg __415353_415353;
   reg _415354_415354 ; 
   reg __415354_415354;
   reg _415355_415355 ; 
   reg __415355_415355;
   reg _415356_415356 ; 
   reg __415356_415356;
   reg _415357_415357 ; 
   reg __415357_415357;
   reg _415358_415358 ; 
   reg __415358_415358;
   reg _415359_415359 ; 
   reg __415359_415359;
   reg _415360_415360 ; 
   reg __415360_415360;
   reg _415361_415361 ; 
   reg __415361_415361;
   reg _415362_415362 ; 
   reg __415362_415362;
   reg _415363_415363 ; 
   reg __415363_415363;
   reg _415364_415364 ; 
   reg __415364_415364;
   reg _415365_415365 ; 
   reg __415365_415365;
   reg _415366_415366 ; 
   reg __415366_415366;
   reg _415367_415367 ; 
   reg __415367_415367;
   reg _415368_415368 ; 
   reg __415368_415368;
   reg _415369_415369 ; 
   reg __415369_415369;
   reg _415370_415370 ; 
   reg __415370_415370;
   reg _415371_415371 ; 
   reg __415371_415371;
   reg _415372_415372 ; 
   reg __415372_415372;
   reg _415373_415373 ; 
   reg __415373_415373;
   reg _415374_415374 ; 
   reg __415374_415374;
   reg _415375_415375 ; 
   reg __415375_415375;
   reg _415376_415376 ; 
   reg __415376_415376;
   reg _415377_415377 ; 
   reg __415377_415377;
   reg _415378_415378 ; 
   reg __415378_415378;
   reg _415379_415379 ; 
   reg __415379_415379;
   reg _415380_415380 ; 
   reg __415380_415380;
   reg _415381_415381 ; 
   reg __415381_415381;
   reg _415382_415382 ; 
   reg __415382_415382;
   reg _415383_415383 ; 
   reg __415383_415383;
   reg _415384_415384 ; 
   reg __415384_415384;
   reg _415385_415385 ; 
   reg __415385_415385;
   reg _415386_415386 ; 
   reg __415386_415386;
   reg _415387_415387 ; 
   reg __415387_415387;
   reg _415388_415388 ; 
   reg __415388_415388;
   reg _415389_415389 ; 
   reg __415389_415389;
   reg _415390_415390 ; 
   reg __415390_415390;
   reg _415391_415391 ; 
   reg __415391_415391;
   reg _415392_415392 ; 
   reg __415392_415392;
   reg _415393_415393 ; 
   reg __415393_415393;
   reg _415394_415394 ; 
   reg __415394_415394;
   reg _415395_415395 ; 
   reg __415395_415395;
   reg _415396_415396 ; 
   reg __415396_415396;
   reg _415397_415397 ; 
   reg __415397_415397;
   reg _415398_415398 ; 
   reg __415398_415398;
   reg _415399_415399 ; 
   reg __415399_415399;
   reg _415400_415400 ; 
   reg __415400_415400;
   reg _415401_415401 ; 
   reg __415401_415401;
   reg _415402_415402 ; 
   reg __415402_415402;
   reg _415403_415403 ; 
   reg __415403_415403;
   reg _415404_415404 ; 
   reg __415404_415404;
   reg _415405_415405 ; 
   reg __415405_415405;
   reg _415406_415406 ; 
   reg __415406_415406;
   reg _415407_415407 ; 
   reg __415407_415407;
   reg _415408_415408 ; 
   reg __415408_415408;
   reg _415409_415409 ; 
   reg __415409_415409;
   reg _415410_415410 ; 
   reg __415410_415410;
   reg _415411_415411 ; 
   reg __415411_415411;
   reg _415412_415412 ; 
   reg __415412_415412;
   reg _415413_415413 ; 
   reg __415413_415413;
   reg _415414_415414 ; 
   reg __415414_415414;
   reg _415415_415415 ; 
   reg __415415_415415;
   reg _415416_415416 ; 
   reg __415416_415416;
   reg _415417_415417 ; 
   reg __415417_415417;
   reg _415418_415418 ; 
   reg __415418_415418;
   reg _415419_415419 ; 
   reg __415419_415419;
   reg _415420_415420 ; 
   reg __415420_415420;
   reg _415421_415421 ; 
   reg __415421_415421;
   reg _415422_415422 ; 
   reg __415422_415422;
   reg _415423_415423 ; 
   reg __415423_415423;
   reg _415424_415424 ; 
   reg __415424_415424;
   reg _415425_415425 ; 
   reg __415425_415425;
   reg _415426_415426 ; 
   reg __415426_415426;
   reg _415427_415427 ; 
   reg __415427_415427;
   reg _415428_415428 ; 
   reg __415428_415428;
   reg _415429_415429 ; 
   reg __415429_415429;
   reg _415430_415430 ; 
   reg __415430_415430;
   reg _415431_415431 ; 
   reg __415431_415431;
   reg _415432_415432 ; 
   reg __415432_415432;
   reg _415433_415433 ; 
   reg __415433_415433;
   reg _415434_415434 ; 
   reg __415434_415434;
   reg _415435_415435 ; 
   reg __415435_415435;
   reg _415436_415436 ; 
   reg __415436_415436;
   reg _415437_415437 ; 
   reg __415437_415437;
   reg _415438_415438 ; 
   reg __415438_415438;
   reg _415439_415439 ; 
   reg __415439_415439;
   reg _415440_415440 ; 
   reg __415440_415440;
   reg _415441_415441 ; 
   reg __415441_415441;
   reg _415442_415442 ; 
   reg __415442_415442;
   reg _415443_415443 ; 
   reg __415443_415443;
   reg _415444_415444 ; 
   reg __415444_415444;
   reg _415445_415445 ; 
   reg __415445_415445;
   reg _415446_415446 ; 
   reg __415446_415446;
   reg _415447_415447 ; 
   reg __415447_415447;
   reg _415448_415448 ; 
   reg __415448_415448;
   reg _415449_415449 ; 
   reg __415449_415449;
   reg _415450_415450 ; 
   reg __415450_415450;
   reg _415451_415451 ; 
   reg __415451_415451;
   reg _415452_415452 ; 
   reg __415452_415452;
   reg _415453_415453 ; 
   reg __415453_415453;
   reg _415454_415454 ; 
   reg __415454_415454;
   reg _415455_415455 ; 
   reg __415455_415455;
   reg _415456_415456 ; 
   reg __415456_415456;
   reg _415457_415457 ; 
   reg __415457_415457;
   reg _415458_415458 ; 
   reg __415458_415458;
   reg _415459_415459 ; 
   reg __415459_415459;
   reg _415460_415460 ; 
   reg __415460_415460;
   reg _415461_415461 ; 
   reg __415461_415461;
   reg _415462_415462 ; 
   reg __415462_415462;
   reg _415463_415463 ; 
   reg __415463_415463;
   reg _415464_415464 ; 
   reg __415464_415464;
   reg _415465_415465 ; 
   reg __415465_415465;
   reg _415466_415466 ; 
   reg __415466_415466;
   reg _415467_415467 ; 
   reg __415467_415467;
   reg _415468_415468 ; 
   reg __415468_415468;
   reg _415469_415469 ; 
   reg __415469_415469;
   reg _415470_415470 ; 
   reg __415470_415470;
   reg _415471_415471 ; 
   reg __415471_415471;
   reg _415472_415472 ; 
   reg __415472_415472;
   reg _415473_415473 ; 
   reg __415473_415473;
   reg _415474_415474 ; 
   reg __415474_415474;
   reg _415475_415475 ; 
   reg __415475_415475;
   reg _415476_415476 ; 
   reg __415476_415476;
   reg _415477_415477 ; 
   reg __415477_415477;
   reg _415478_415478 ; 
   reg __415478_415478;
   reg _415479_415479 ; 
   reg __415479_415479;
   reg _415480_415480 ; 
   reg __415480_415480;
   reg _415481_415481 ; 
   reg __415481_415481;
   reg _415482_415482 ; 
   reg __415482_415482;
   reg _415483_415483 ; 
   reg __415483_415483;
   reg _415484_415484 ; 
   reg __415484_415484;
   reg _415485_415485 ; 
   reg __415485_415485;
   reg _415486_415486 ; 
   reg __415486_415486;
   reg _415487_415487 ; 
   reg __415487_415487;
   reg _415488_415488 ; 
   reg __415488_415488;
   reg _415489_415489 ; 
   reg __415489_415489;
   reg _415490_415490 ; 
   reg __415490_415490;
   reg _415491_415491 ; 
   reg __415491_415491;
   reg _415492_415492 ; 
   reg __415492_415492;
   reg _415493_415493 ; 
   reg __415493_415493;
   reg _415494_415494 ; 
   reg __415494_415494;
   reg _415495_415495 ; 
   reg __415495_415495;
   reg _415496_415496 ; 
   reg __415496_415496;
   reg _415497_415497 ; 
   reg __415497_415497;
   reg _415498_415498 ; 
   reg __415498_415498;
   reg _415499_415499 ; 
   reg __415499_415499;
   reg _415500_415500 ; 
   reg __415500_415500;
   reg _415501_415501 ; 
   reg __415501_415501;
   reg _415502_415502 ; 
   reg __415502_415502;
   reg _415503_415503 ; 
   reg __415503_415503;
   reg _415504_415504 ; 
   reg __415504_415504;
   reg _415505_415505 ; 
   reg __415505_415505;
   reg _415506_415506 ; 
   reg __415506_415506;
   reg _415507_415507 ; 
   reg __415507_415507;
   reg _415508_415508 ; 
   reg __415508_415508;
   reg _415509_415509 ; 
   reg __415509_415509;
   reg _415510_415510 ; 
   reg __415510_415510;
   reg _415511_415511 ; 
   reg __415511_415511;
   reg _415512_415512 ; 
   reg __415512_415512;
   reg _415513_415513 ; 
   reg __415513_415513;
   reg _415514_415514 ; 
   reg __415514_415514;
   reg _415515_415515 ; 
   reg __415515_415515;
   reg _415516_415516 ; 
   reg __415516_415516;
   reg _415517_415517 ; 
   reg __415517_415517;
   reg _415518_415518 ; 
   reg __415518_415518;
   reg _415519_415519 ; 
   reg __415519_415519;
   reg _415520_415520 ; 
   reg __415520_415520;
   reg _415521_415521 ; 
   reg __415521_415521;
   reg _415522_415522 ; 
   reg __415522_415522;
   reg _415523_415523 ; 
   reg __415523_415523;
   reg _415524_415524 ; 
   reg __415524_415524;
   reg _415525_415525 ; 
   reg __415525_415525;
   reg _415526_415526 ; 
   reg __415526_415526;
   reg _415527_415527 ; 
   reg __415527_415527;
   reg _415528_415528 ; 
   reg __415528_415528;
   reg _415529_415529 ; 
   reg __415529_415529;
   reg _415530_415530 ; 
   reg __415530_415530;
   reg _415531_415531 ; 
   reg __415531_415531;
   reg _415532_415532 ; 
   reg __415532_415532;
   reg _415533_415533 ; 
   reg __415533_415533;
   reg _415534_415534 ; 
   reg __415534_415534;
   reg _415535_415535 ; 
   reg __415535_415535;
   reg _415536_415536 ; 
   reg __415536_415536;
   reg _415537_415537 ; 
   reg __415537_415537;
   reg _415538_415538 ; 
   reg __415538_415538;
   reg _415539_415539 ; 
   reg __415539_415539;
   reg _415540_415540 ; 
   reg __415540_415540;
   reg _415541_415541 ; 
   reg __415541_415541;
   reg _415542_415542 ; 
   reg __415542_415542;
   reg _415543_415543 ; 
   reg __415543_415543;
   reg _415544_415544 ; 
   reg __415544_415544;
   reg _415545_415545 ; 
   reg __415545_415545;
   reg _415546_415546 ; 
   reg __415546_415546;
   reg _415547_415547 ; 
   reg __415547_415547;
   reg _415548_415548 ; 
   reg __415548_415548;
   reg _415549_415549 ; 
   reg __415549_415549;
   reg _415550_415550 ; 
   reg __415550_415550;
   reg _415551_415551 ; 
   reg __415551_415551;
   reg _415552_415552 ; 
   reg __415552_415552;
   reg _415553_415553 ; 
   reg __415553_415553;
   reg _415554_415554 ; 
   reg __415554_415554;
   reg _415555_415555 ; 
   reg __415555_415555;
   reg _415556_415556 ; 
   reg __415556_415556;
   reg _415557_415557 ; 
   reg __415557_415557;
   reg _415558_415558 ; 
   reg __415558_415558;
   reg _415559_415559 ; 
   reg __415559_415559;
   reg _415560_415560 ; 
   reg __415560_415560;
   reg _415561_415561 ; 
   reg __415561_415561;
   reg _415562_415562 ; 
   reg __415562_415562;
   reg _415563_415563 ; 
   reg __415563_415563;
   reg _415564_415564 ; 
   reg __415564_415564;
   reg _415565_415565 ; 
   reg __415565_415565;
   reg _415566_415566 ; 
   reg __415566_415566;
   reg _415567_415567 ; 
   reg __415567_415567;
   reg _415568_415568 ; 
   reg __415568_415568;
   reg _415569_415569 ; 
   reg __415569_415569;
   reg _415570_415570 ; 
   reg __415570_415570;
   reg _415571_415571 ; 
   reg __415571_415571;
   reg _415572_415572 ; 
   reg __415572_415572;
   reg _415573_415573 ; 
   reg __415573_415573;
   reg _415574_415574 ; 
   reg __415574_415574;
   reg _415575_415575 ; 
   reg __415575_415575;
   reg _415576_415576 ; 
   reg __415576_415576;
   reg _415577_415577 ; 
   reg __415577_415577;
   reg _415578_415578 ; 
   reg __415578_415578;
   reg _415579_415579 ; 
   reg __415579_415579;
   reg _415580_415580 ; 
   reg __415580_415580;
   reg _415581_415581 ; 
   reg __415581_415581;
   reg _415582_415582 ; 
   reg __415582_415582;
   reg _415583_415583 ; 
   reg __415583_415583;
   reg _415584_415584 ; 
   reg __415584_415584;
   reg _415585_415585 ; 
   reg __415585_415585;
   reg _415586_415586 ; 
   reg __415586_415586;
   reg _415587_415587 ; 
   reg __415587_415587;
   reg _415588_415588 ; 
   reg __415588_415588;
   reg _415589_415589 ; 
   reg __415589_415589;
   reg _415590_415590 ; 
   reg __415590_415590;
   reg _415591_415591 ; 
   reg __415591_415591;
   reg _415592_415592 ; 
   reg __415592_415592;
   reg _415593_415593 ; 
   reg __415593_415593;
   reg _415594_415594 ; 
   reg __415594_415594;
   reg _415595_415595 ; 
   reg __415595_415595;
   reg _415596_415596 ; 
   reg __415596_415596;
   reg _415597_415597 ; 
   reg __415597_415597;
   reg _415598_415598 ; 
   reg __415598_415598;
   reg _415599_415599 ; 
   reg __415599_415599;
   reg _415600_415600 ; 
   reg __415600_415600;
   reg _415601_415601 ; 
   reg __415601_415601;
   reg _415602_415602 ; 
   reg __415602_415602;
   reg _415603_415603 ; 
   reg __415603_415603;
   reg _415604_415604 ; 
   reg __415604_415604;
   reg _415605_415605 ; 
   reg __415605_415605;
   reg _415606_415606 ; 
   reg __415606_415606;
   reg _415607_415607 ; 
   reg __415607_415607;
   reg _415608_415608 ; 
   reg __415608_415608;
   reg _415609_415609 ; 
   reg __415609_415609;
   reg _415610_415610 ; 
   reg __415610_415610;
   reg _415611_415611 ; 
   reg __415611_415611;
   reg _415612_415612 ; 
   reg __415612_415612;
   reg _415613_415613 ; 
   reg __415613_415613;
   reg _415614_415614 ; 
   reg __415614_415614;
   reg _415615_415615 ; 
   reg __415615_415615;
   reg _415616_415616 ; 
   reg __415616_415616;
   reg _415617_415617 ; 
   reg __415617_415617;
   reg _415618_415618 ; 
   reg __415618_415618;
   reg _415619_415619 ; 
   reg __415619_415619;
   reg _415620_415620 ; 
   reg __415620_415620;
   reg _415621_415621 ; 
   reg __415621_415621;
   reg _415622_415622 ; 
   reg __415622_415622;
   reg _415623_415623 ; 
   reg __415623_415623;
   reg _415624_415624 ; 
   reg __415624_415624;
   reg _415625_415625 ; 
   reg __415625_415625;
   reg _415626_415626 ; 
   reg __415626_415626;
   reg _415627_415627 ; 
   reg __415627_415627;
   reg _415628_415628 ; 
   reg __415628_415628;
   reg _415629_415629 ; 
   reg __415629_415629;
   reg _415630_415630 ; 
   reg __415630_415630;
   reg _415631_415631 ; 
   reg __415631_415631;
   reg _415632_415632 ; 
   reg __415632_415632;
   reg _415633_415633 ; 
   reg __415633_415633;
   reg _415634_415634 ; 
   reg __415634_415634;
   reg _415635_415635 ; 
   reg __415635_415635;
   reg _415636_415636 ; 
   reg __415636_415636;
   reg _415637_415637 ; 
   reg __415637_415637;
   reg _415638_415638 ; 
   reg __415638_415638;
   reg _415639_415639 ; 
   reg __415639_415639;
   reg _415640_415640 ; 
   reg __415640_415640;
   reg _415641_415641 ; 
   reg __415641_415641;
   reg _415642_415642 ; 
   reg __415642_415642;
   reg _415643_415643 ; 
   reg __415643_415643;
   reg _415644_415644 ; 
   reg __415644_415644;
   reg _415645_415645 ; 
   reg __415645_415645;
   reg _415646_415646 ; 
   reg __415646_415646;
   reg _415647_415647 ; 
   reg __415647_415647;
   reg _415648_415648 ; 
   reg __415648_415648;
   reg _415649_415649 ; 
   reg __415649_415649;
   reg _415650_415650 ; 
   reg __415650_415650;
   reg _415651_415651 ; 
   reg __415651_415651;
   reg _415652_415652 ; 
   reg __415652_415652;
   reg _415653_415653 ; 
   reg __415653_415653;
   reg _415654_415654 ; 
   reg __415654_415654;
   reg _415655_415655 ; 
   reg __415655_415655;
   reg _415656_415656 ; 
   reg __415656_415656;
   reg _415657_415657 ; 
   reg __415657_415657;
   reg _415658_415658 ; 
   reg __415658_415658;
   reg _415659_415659 ; 
   reg __415659_415659;
   reg _415660_415660 ; 
   reg __415660_415660;
   reg _415661_415661 ; 
   reg __415661_415661;
   reg _415662_415662 ; 
   reg __415662_415662;
   reg _415663_415663 ; 
   reg __415663_415663;
   reg _415664_415664 ; 
   reg __415664_415664;
   reg _415665_415665 ; 
   reg __415665_415665;
   reg _415666_415666 ; 
   reg __415666_415666;
   reg _415667_415667 ; 
   reg __415667_415667;
   reg _415668_415668 ; 
   reg __415668_415668;
   reg _415669_415669 ; 
   reg __415669_415669;
   reg _415670_415670 ; 
   reg __415670_415670;
   reg _415671_415671 ; 
   reg __415671_415671;
   reg _415672_415672 ; 
   reg __415672_415672;
   reg _415673_415673 ; 
   reg __415673_415673;
   reg _415674_415674 ; 
   reg __415674_415674;
   reg _415675_415675 ; 
   reg __415675_415675;
   reg _415676_415676 ; 
   reg __415676_415676;
   reg _415677_415677 ; 
   reg __415677_415677;
   reg _415678_415678 ; 
   reg __415678_415678;
   reg _415679_415679 ; 
   reg __415679_415679;
   reg _415680_415680 ; 
   reg __415680_415680;
   reg _415681_415681 ; 
   reg __415681_415681;
   reg _415682_415682 ; 
   reg __415682_415682;
   reg _415683_415683 ; 
   reg __415683_415683;
   reg _415684_415684 ; 
   reg __415684_415684;
   reg _415685_415685 ; 
   reg __415685_415685;
   reg _415686_415686 ; 
   reg __415686_415686;
   reg _415687_415687 ; 
   reg __415687_415687;
   reg _415688_415688 ; 
   reg __415688_415688;
   reg _415689_415689 ; 
   reg __415689_415689;
   reg _415690_415690 ; 
   reg __415690_415690;
   reg _415691_415691 ; 
   reg __415691_415691;
   reg _415692_415692 ; 
   reg __415692_415692;
   reg _415693_415693 ; 
   reg __415693_415693;
   reg _415694_415694 ; 
   reg __415694_415694;
   reg _415695_415695 ; 
   reg __415695_415695;
   reg _415696_415696 ; 
   reg __415696_415696;
   reg _415697_415697 ; 
   reg __415697_415697;
   reg _415698_415698 ; 
   reg __415698_415698;
   reg _415699_415699 ; 
   reg __415699_415699;
   reg _415700_415700 ; 
   reg __415700_415700;
   reg _415701_415701 ; 
   reg __415701_415701;
   reg _415702_415702 ; 
   reg __415702_415702;
   reg _415703_415703 ; 
   reg __415703_415703;
   reg _415704_415704 ; 
   reg __415704_415704;
   reg _415705_415705 ; 
   reg __415705_415705;
   reg _415706_415706 ; 
   reg __415706_415706;
   reg _415707_415707 ; 
   reg __415707_415707;
   reg _415708_415708 ; 
   reg __415708_415708;
   reg _415709_415709 ; 
   reg __415709_415709;
   reg _415710_415710 ; 
   reg __415710_415710;
   reg _415711_415711 ; 
   reg __415711_415711;
   reg _415712_415712 ; 
   reg __415712_415712;
   reg _415713_415713 ; 
   reg __415713_415713;
   reg _415714_415714 ; 
   reg __415714_415714;
   reg _415715_415715 ; 
   reg __415715_415715;
   reg _415716_415716 ; 
   reg __415716_415716;
   reg _415717_415717 ; 
   reg __415717_415717;
   reg _415718_415718 ; 
   reg __415718_415718;
   reg _415719_415719 ; 
   reg __415719_415719;
   reg _415720_415720 ; 
   reg __415720_415720;
   reg _415721_415721 ; 
   reg __415721_415721;
   reg _415722_415722 ; 
   reg __415722_415722;
   reg _415723_415723 ; 
   reg __415723_415723;
   reg _415724_415724 ; 
   reg __415724_415724;
   reg _415725_415725 ; 
   reg __415725_415725;
   reg _415726_415726 ; 
   reg __415726_415726;
   reg _415727_415727 ; 
   reg __415727_415727;
   reg _415728_415728 ; 
   reg __415728_415728;
   reg _415729_415729 ; 
   reg __415729_415729;
   reg _415730_415730 ; 
   reg __415730_415730;
   reg _415731_415731 ; 
   reg __415731_415731;
   reg _415732_415732 ; 
   reg __415732_415732;
   reg _415733_415733 ; 
   reg __415733_415733;
   reg _415734_415734 ; 
   reg __415734_415734;
   reg _415735_415735 ; 
   reg __415735_415735;
   reg _415736_415736 ; 
   reg __415736_415736;
   reg _415737_415737 ; 
   reg __415737_415737;
   reg _415738_415738 ; 
   reg __415738_415738;
   reg _415739_415739 ; 
   reg __415739_415739;
   reg _415740_415740 ; 
   reg __415740_415740;
   reg _415741_415741 ; 
   reg __415741_415741;
   reg _415742_415742 ; 
   reg __415742_415742;
   reg _415743_415743 ; 
   reg __415743_415743;
   reg _415744_415744 ; 
   reg __415744_415744;
   reg _415745_415745 ; 
   reg __415745_415745;
   reg _415746_415746 ; 
   reg __415746_415746;
   reg _415747_415747 ; 
   reg __415747_415747;
   reg _415748_415748 ; 
   reg __415748_415748;
   reg _415749_415749 ; 
   reg __415749_415749;
   reg _415750_415750 ; 
   reg __415750_415750;
   reg _415751_415751 ; 
   reg __415751_415751;
   reg _415752_415752 ; 
   reg __415752_415752;
   reg _415753_415753 ; 
   reg __415753_415753;
   reg _415754_415754 ; 
   reg __415754_415754;
   reg _415755_415755 ; 
   reg __415755_415755;
   reg _415756_415756 ; 
   reg __415756_415756;
   reg _415757_415757 ; 
   reg __415757_415757;
   reg _415758_415758 ; 
   reg __415758_415758;
   reg _415759_415759 ; 
   reg __415759_415759;
   reg _415760_415760 ; 
   reg __415760_415760;
   reg _415761_415761 ; 
   reg __415761_415761;
   reg _415762_415762 ; 
   reg __415762_415762;
   reg _415763_415763 ; 
   reg __415763_415763;
   reg _415764_415764 ; 
   reg __415764_415764;
   reg _415765_415765 ; 
   reg __415765_415765;
   reg _415766_415766 ; 
   reg __415766_415766;
   reg _415767_415767 ; 
   reg __415767_415767;
   reg _415768_415768 ; 
   reg __415768_415768;
   reg _415769_415769 ; 
   reg __415769_415769;
   reg _415770_415770 ; 
   reg __415770_415770;
   reg _415771_415771 ; 
   reg __415771_415771;
   reg _415772_415772 ; 
   reg __415772_415772;
   reg _415773_415773 ; 
   reg __415773_415773;
   reg _415774_415774 ; 
   reg __415774_415774;
   reg _415775_415775 ; 
   reg __415775_415775;
   reg _415776_415776 ; 
   reg __415776_415776;
   reg _415777_415777 ; 
   reg __415777_415777;
   reg _415778_415778 ; 
   reg __415778_415778;
   reg _415779_415779 ; 
   reg __415779_415779;
   reg _415780_415780 ; 
   reg __415780_415780;
   reg _415781_415781 ; 
   reg __415781_415781;
   reg _415782_415782 ; 
   reg __415782_415782;
   reg _415783_415783 ; 
   reg __415783_415783;
   reg _415784_415784 ; 
   reg __415784_415784;
   reg _415785_415785 ; 
   reg __415785_415785;
   reg _415786_415786 ; 
   reg __415786_415786;
   reg _415787_415787 ; 
   reg __415787_415787;
   reg _415788_415788 ; 
   reg __415788_415788;
   reg _415789_415789 ; 
   reg __415789_415789;
   reg _415790_415790 ; 
   reg __415790_415790;
   reg _415791_415791 ; 
   reg __415791_415791;
   reg _415792_415792 ; 
   reg __415792_415792;
   reg _415793_415793 ; 
   reg __415793_415793;
   reg _415794_415794 ; 
   reg __415794_415794;
   reg _415795_415795 ; 
   reg __415795_415795;
   reg _415796_415796 ; 
   reg __415796_415796;
   reg _415797_415797 ; 
   reg __415797_415797;
   reg _415798_415798 ; 
   reg __415798_415798;
   reg _415799_415799 ; 
   reg __415799_415799;
   reg _415800_415800 ; 
   reg __415800_415800;
   reg _415801_415801 ; 
   reg __415801_415801;
   reg _415802_415802 ; 
   reg __415802_415802;
   reg _415803_415803 ; 
   reg __415803_415803;
   reg _415804_415804 ; 
   reg __415804_415804;
   reg _415805_415805 ; 
   reg __415805_415805;
   reg _415806_415806 ; 
   reg __415806_415806;
   reg _415807_415807 ; 
   reg __415807_415807;
   reg _415808_415808 ; 
   reg __415808_415808;
   reg _415809_415809 ; 
   reg __415809_415809;
   reg _415810_415810 ; 
   reg __415810_415810;
   reg _415811_415811 ; 
   reg __415811_415811;
   reg _415812_415812 ; 
   reg __415812_415812;
   reg _415813_415813 ; 
   reg __415813_415813;
   reg _415814_415814 ; 
   reg __415814_415814;
   reg _415815_415815 ; 
   reg __415815_415815;
   reg _415816_415816 ; 
   reg __415816_415816;
   reg _415817_415817 ; 
   reg __415817_415817;
   reg _415818_415818 ; 
   reg __415818_415818;
   reg _415819_415819 ; 
   reg __415819_415819;
   reg _415820_415820 ; 
   reg __415820_415820;
   reg _415821_415821 ; 
   reg __415821_415821;
   reg _415822_415822 ; 
   reg __415822_415822;
   reg _415823_415823 ; 
   reg __415823_415823;
   reg _415824_415824 ; 
   reg __415824_415824;
   reg _415825_415825 ; 
   reg __415825_415825;
   reg _415826_415826 ; 
   reg __415826_415826;
   reg _415827_415827 ; 
   reg __415827_415827;
   reg _415828_415828 ; 
   reg __415828_415828;
   reg _415829_415829 ; 
   reg __415829_415829;
   reg _415830_415830 ; 
   reg __415830_415830;
   reg _415831_415831 ; 
   reg __415831_415831;
   reg _415832_415832 ; 
   reg __415832_415832;
   reg _415833_415833 ; 
   reg __415833_415833;
   reg _415834_415834 ; 
   reg __415834_415834;
   reg _415835_415835 ; 
   reg __415835_415835;
   reg _415836_415836 ; 
   reg __415836_415836;
   reg _415837_415837 ; 
   reg __415837_415837;
   reg _415838_415838 ; 
   reg __415838_415838;
   reg _415839_415839 ; 
   reg __415839_415839;
   reg _415840_415840 ; 
   reg __415840_415840;
   reg _415841_415841 ; 
   reg __415841_415841;
   reg _415842_415842 ; 
   reg __415842_415842;
   reg _415843_415843 ; 
   reg __415843_415843;
   reg _415844_415844 ; 
   reg __415844_415844;
   reg _415845_415845 ; 
   reg __415845_415845;
   reg _415846_415846 ; 
   reg __415846_415846;
   reg _415847_415847 ; 
   reg __415847_415847;
   reg _415848_415848 ; 
   reg __415848_415848;
   reg _415849_415849 ; 
   reg __415849_415849;
   reg _415850_415850 ; 
   reg __415850_415850;
   reg _415851_415851 ; 
   reg __415851_415851;
   reg _415852_415852 ; 
   reg __415852_415852;
   reg _415853_415853 ; 
   reg __415853_415853;
   reg _415854_415854 ; 
   reg __415854_415854;
   reg _415855_415855 ; 
   reg __415855_415855;
   reg _415856_415856 ; 
   reg __415856_415856;
   reg _415857_415857 ; 
   reg __415857_415857;
   reg _415858_415858 ; 
   reg __415858_415858;
   reg _415859_415859 ; 
   reg __415859_415859;
   reg _415860_415860 ; 
   reg __415860_415860;
   reg _415861_415861 ; 
   reg __415861_415861;
   reg _415862_415862 ; 
   reg __415862_415862;
   reg _415863_415863 ; 
   reg __415863_415863;
   reg _415864_415864 ; 
   reg __415864_415864;
   reg _415865_415865 ; 
   reg __415865_415865;
   reg _415866_415866 ; 
   reg __415866_415866;
   reg _415867_415867 ; 
   reg __415867_415867;
   reg _415868_415868 ; 
   reg __415868_415868;
   reg _415869_415869 ; 
   reg __415869_415869;
   reg _415870_415870 ; 
   reg __415870_415870;
   reg _415871_415871 ; 
   reg __415871_415871;
   reg _415872_415872 ; 
   reg __415872_415872;
   reg _415873_415873 ; 
   reg __415873_415873;
   reg _415874_415874 ; 
   reg __415874_415874;
   reg _415875_415875 ; 
   reg __415875_415875;
   reg _415876_415876 ; 
   reg __415876_415876;
   reg _415877_415877 ; 
   reg __415877_415877;
   reg _415878_415878 ; 
   reg __415878_415878;
   reg _415879_415879 ; 
   reg __415879_415879;
   reg _415880_415880 ; 
   reg __415880_415880;
   reg _415881_415881 ; 
   reg __415881_415881;
   reg _415882_415882 ; 
   reg __415882_415882;
   reg _415883_415883 ; 
   reg __415883_415883;
   reg _415884_415884 ; 
   reg __415884_415884;
   reg _415885_415885 ; 
   reg __415885_415885;
   reg _415886_415886 ; 
   reg __415886_415886;
   reg _415887_415887 ; 
   reg __415887_415887;
   reg _415888_415888 ; 
   reg __415888_415888;
   reg _415889_415889 ; 
   reg __415889_415889;
   reg _415890_415890 ; 
   reg __415890_415890;
   reg _415891_415891 ; 
   reg __415891_415891;
   reg _415892_415892 ; 
   reg __415892_415892;
   reg _415893_415893 ; 
   reg __415893_415893;
   reg _415894_415894 ; 
   reg __415894_415894;
   reg _415895_415895 ; 
   reg __415895_415895;
   reg _415896_415896 ; 
   reg __415896_415896;
   reg _415897_415897 ; 
   reg __415897_415897;
   reg _415898_415898 ; 
   reg __415898_415898;
   reg _415899_415899 ; 
   reg __415899_415899;
   reg _415900_415900 ; 
   reg __415900_415900;
   reg _415901_415901 ; 
   reg __415901_415901;
   reg _415902_415902 ; 
   reg __415902_415902;
   reg _415903_415903 ; 
   reg __415903_415903;
   reg _415904_415904 ; 
   reg __415904_415904;
   reg _415905_415905 ; 
   reg __415905_415905;
   reg _415906_415906 ; 
   reg __415906_415906;
   reg _415907_415907 ; 
   reg __415907_415907;
   reg _415908_415908 ; 
   reg __415908_415908;
   reg _415909_415909 ; 
   reg __415909_415909;
   reg _415910_415910 ; 
   reg __415910_415910;
   reg _415911_415911 ; 
   reg __415911_415911;
   reg _415912_415912 ; 
   reg __415912_415912;
   reg _415913_415913 ; 
   reg __415913_415913;
   reg _415914_415914 ; 
   reg __415914_415914;
   reg _415915_415915 ; 
   reg __415915_415915;
   reg _415916_415916 ; 
   reg __415916_415916;
   reg _415917_415917 ; 
   reg __415917_415917;
   reg _415918_415918 ; 
   reg __415918_415918;
   reg _415919_415919 ; 
   reg __415919_415919;
   reg _415920_415920 ; 
   reg __415920_415920;
   reg _415921_415921 ; 
   reg __415921_415921;
   reg _415922_415922 ; 
   reg __415922_415922;
   reg _415923_415923 ; 
   reg __415923_415923;
   reg _415924_415924 ; 
   reg __415924_415924;
   reg _415925_415925 ; 
   reg __415925_415925;
   reg _415926_415926 ; 
   reg __415926_415926;
   reg _415927_415927 ; 
   reg __415927_415927;
   reg _415928_415928 ; 
   reg __415928_415928;
   reg _415929_415929 ; 
   reg __415929_415929;
   reg _415930_415930 ; 
   reg __415930_415930;
   reg _415931_415931 ; 
   reg __415931_415931;
   reg _415932_415932 ; 
   reg __415932_415932;
   reg _415933_415933 ; 
   reg __415933_415933;
   reg _415934_415934 ; 
   reg __415934_415934;
   reg _415935_415935 ; 
   reg __415935_415935;
   reg _415936_415936 ; 
   reg __415936_415936;
   reg _415937_415937 ; 
   reg __415937_415937;
   reg _415938_415938 ; 
   reg __415938_415938;
   reg _415939_415939 ; 
   reg __415939_415939;
   reg _415940_415940 ; 
   reg __415940_415940;
   reg _415941_415941 ; 
   reg __415941_415941;
   reg _415942_415942 ; 
   reg __415942_415942;
   reg _415943_415943 ; 
   reg __415943_415943;
   reg _415944_415944 ; 
   reg __415944_415944;
   reg _415945_415945 ; 
   reg __415945_415945;
   reg _415946_415946 ; 
   reg __415946_415946;
   reg _415947_415947 ; 
   reg __415947_415947;
   reg _415948_415948 ; 
   reg __415948_415948;
   reg _415949_415949 ; 
   reg __415949_415949;
   reg _415950_415950 ; 
   reg __415950_415950;
   reg _415951_415951 ; 
   reg __415951_415951;
   reg _415952_415952 ; 
   reg __415952_415952;
   reg _415953_415953 ; 
   reg __415953_415953;
   reg _415954_415954 ; 
   reg __415954_415954;
   reg _415955_415955 ; 
   reg __415955_415955;
   reg _415956_415956 ; 
   reg __415956_415956;
   reg _415957_415957 ; 
   reg __415957_415957;
   reg _415958_415958 ; 
   reg __415958_415958;
   reg _415959_415959 ; 
   reg __415959_415959;
   reg _415960_415960 ; 
   reg __415960_415960;
   reg _415961_415961 ; 
   reg __415961_415961;
   reg _415962_415962 ; 
   reg __415962_415962;
   reg _415963_415963 ; 
   reg __415963_415963;
   reg _415964_415964 ; 
   reg __415964_415964;
   reg _415965_415965 ; 
   reg __415965_415965;
   reg _415966_415966 ; 
   reg __415966_415966;
   reg _415967_415967 ; 
   reg __415967_415967;
   reg _415968_415968 ; 
   reg __415968_415968;
   reg _415969_415969 ; 
   reg __415969_415969;
   reg _415970_415970 ; 
   reg __415970_415970;
   reg _415971_415971 ; 
   reg __415971_415971;
   reg _415972_415972 ; 
   reg __415972_415972;
   reg _415973_415973 ; 
   reg __415973_415973;
   reg _415974_415974 ; 
   reg __415974_415974;
   reg _415975_415975 ; 
   reg __415975_415975;
   reg _415976_415976 ; 
   reg __415976_415976;
   reg _415977_415977 ; 
   reg __415977_415977;
   reg _415978_415978 ; 
   reg __415978_415978;
   reg _415979_415979 ; 
   reg __415979_415979;
   reg _415980_415980 ; 
   reg __415980_415980;
   reg _415981_415981 ; 
   reg __415981_415981;
   reg _415982_415982 ; 
   reg __415982_415982;
   reg _415983_415983 ; 
   reg __415983_415983;
   reg _415984_415984 ; 
   reg __415984_415984;
   reg _415985_415985 ; 
   reg __415985_415985;
   reg _415986_415986 ; 
   reg __415986_415986;
   reg _415987_415987 ; 
   reg __415987_415987;
   reg _415988_415988 ; 
   reg __415988_415988;
   reg _415989_415989 ; 
   reg __415989_415989;
   reg _415990_415990 ; 
   reg __415990_415990;
   reg _415991_415991 ; 
   reg __415991_415991;
   reg _415992_415992 ; 
   reg __415992_415992;
   reg _415993_415993 ; 
   reg __415993_415993;
   reg _415994_415994 ; 
   reg __415994_415994;
   reg _415995_415995 ; 
   reg __415995_415995;
   reg _415996_415996 ; 
   reg __415996_415996;
   reg _415997_415997 ; 
   reg __415997_415997;
   reg _415998_415998 ; 
   reg __415998_415998;
   reg _415999_415999 ; 
   reg __415999_415999;
   reg _416000_416000 ; 
   reg __416000_416000;
   reg _416001_416001 ; 
   reg __416001_416001;
   reg _416002_416002 ; 
   reg __416002_416002;
   reg _416003_416003 ; 
   reg __416003_416003;
   reg _416004_416004 ; 
   reg __416004_416004;
   reg _416005_416005 ; 
   reg __416005_416005;
   reg _416006_416006 ; 
   reg __416006_416006;
   reg _416007_416007 ; 
   reg __416007_416007;
   reg _416008_416008 ; 
   reg __416008_416008;
   reg _416009_416009 ; 
   reg __416009_416009;
   reg _416010_416010 ; 
   reg __416010_416010;
   reg _416011_416011 ; 
   reg __416011_416011;
   reg _416012_416012 ; 
   reg __416012_416012;
   reg _416013_416013 ; 
   reg __416013_416013;
   reg _416014_416014 ; 
   reg __416014_416014;
   reg _416015_416015 ; 
   reg __416015_416015;
   reg _416016_416016 ; 
   reg __416016_416016;
   reg _416017_416017 ; 
   reg __416017_416017;
   reg _416018_416018 ; 
   reg __416018_416018;
   reg _416019_416019 ; 
   reg __416019_416019;
   reg _416020_416020 ; 
   reg __416020_416020;
   reg _416021_416021 ; 
   reg __416021_416021;
   reg _416022_416022 ; 
   reg __416022_416022;
   reg _416023_416023 ; 
   reg __416023_416023;
   reg _416024_416024 ; 
   reg __416024_416024;
   reg _416025_416025 ; 
   reg __416025_416025;
   reg _416026_416026 ; 
   reg __416026_416026;
   reg _416027_416027 ; 
   reg __416027_416027;
   reg _416028_416028 ; 
   reg __416028_416028;
   reg _416029_416029 ; 
   reg __416029_416029;
   reg _416030_416030 ; 
   reg __416030_416030;
   reg _416031_416031 ; 
   reg __416031_416031;
   reg _416032_416032 ; 
   reg __416032_416032;
   reg _416033_416033 ; 
   reg __416033_416033;
   reg _416034_416034 ; 
   reg __416034_416034;
   reg _416035_416035 ; 
   reg __416035_416035;
   reg _416036_416036 ; 
   reg __416036_416036;
   reg _416037_416037 ; 
   reg __416037_416037;
   reg _416038_416038 ; 
   reg __416038_416038;
   reg _416039_416039 ; 
   reg __416039_416039;
   reg _416040_416040 ; 
   reg __416040_416040;
   reg _416041_416041 ; 
   reg __416041_416041;
   reg _416042_416042 ; 
   reg __416042_416042;
   reg _416043_416043 ; 
   reg __416043_416043;
   reg _416044_416044 ; 
   reg __416044_416044;
   reg _416045_416045 ; 
   reg __416045_416045;
   reg _416046_416046 ; 
   reg __416046_416046;
   reg _416047_416047 ; 
   reg __416047_416047;
   reg _416048_416048 ; 
   reg __416048_416048;
   reg _416049_416049 ; 
   reg __416049_416049;
   reg _416050_416050 ; 
   reg __416050_416050;
   reg _416051_416051 ; 
   reg __416051_416051;
   reg _416052_416052 ; 
   reg __416052_416052;
   reg _416053_416053 ; 
   reg __416053_416053;
   reg _416054_416054 ; 
   reg __416054_416054;
   reg _416055_416055 ; 
   reg __416055_416055;
   reg _416056_416056 ; 
   reg __416056_416056;
   reg _416057_416057 ; 
   reg __416057_416057;
   reg _416058_416058 ; 
   reg __416058_416058;
   reg _416059_416059 ; 
   reg __416059_416059;
   reg _416060_416060 ; 
   reg __416060_416060;
   reg _416061_416061 ; 
   reg __416061_416061;
   reg _416062_416062 ; 
   reg __416062_416062;
   reg _416063_416063 ; 
   reg __416063_416063;
   reg _416064_416064 ; 
   reg __416064_416064;
   reg _416065_416065 ; 
   reg __416065_416065;
   reg _416066_416066 ; 
   reg __416066_416066;
   reg _416067_416067 ; 
   reg __416067_416067;
   reg _416068_416068 ; 
   reg __416068_416068;
   reg _416069_416069 ; 
   reg __416069_416069;
   reg _416070_416070 ; 
   reg __416070_416070;
   reg _416071_416071 ; 
   reg __416071_416071;
   reg _416072_416072 ; 
   reg __416072_416072;
   reg _416073_416073 ; 
   reg __416073_416073;
   reg _416074_416074 ; 
   reg __416074_416074;
   reg _416075_416075 ; 
   reg __416075_416075;
   reg _416076_416076 ; 
   reg __416076_416076;
   reg _416077_416077 ; 
   reg __416077_416077;
   reg _416078_416078 ; 
   reg __416078_416078;
   reg _416079_416079 ; 
   reg __416079_416079;
   reg _416080_416080 ; 
   reg __416080_416080;
   reg _416081_416081 ; 
   reg __416081_416081;
   reg _416082_416082 ; 
   reg __416082_416082;
   reg _416083_416083 ; 
   reg __416083_416083;
   reg _416084_416084 ; 
   reg __416084_416084;
   reg _416085_416085 ; 
   reg __416085_416085;
   reg _416086_416086 ; 
   reg __416086_416086;
   reg _416087_416087 ; 
   reg __416087_416087;
   reg _416088_416088 ; 
   reg __416088_416088;
   reg _416089_416089 ; 
   reg __416089_416089;
   reg _416090_416090 ; 
   reg __416090_416090;
   reg _416091_416091 ; 
   reg __416091_416091;
   reg _416092_416092 ; 
   reg __416092_416092;
   reg _416093_416093 ; 
   reg __416093_416093;
   reg _416094_416094 ; 
   reg __416094_416094;
   reg _416095_416095 ; 
   reg __416095_416095;
   reg _416096_416096 ; 
   reg __416096_416096;
   reg _416097_416097 ; 
   reg __416097_416097;
   reg _416098_416098 ; 
   reg __416098_416098;
   reg _416099_416099 ; 
   reg __416099_416099;
   reg _416100_416100 ; 
   reg __416100_416100;
   reg _416101_416101 ; 
   reg __416101_416101;
   reg _416102_416102 ; 
   reg __416102_416102;
   reg _416103_416103 ; 
   reg __416103_416103;
   reg _416104_416104 ; 
   reg __416104_416104;
   reg _416105_416105 ; 
   reg __416105_416105;
   reg _416106_416106 ; 
   reg __416106_416106;
   reg _416107_416107 ; 
   reg __416107_416107;
   reg _416108_416108 ; 
   reg __416108_416108;
   reg _416109_416109 ; 
   reg __416109_416109;
   reg _416110_416110 ; 
   reg __416110_416110;
   reg _416111_416111 ; 
   reg __416111_416111;
   reg _416112_416112 ; 
   reg __416112_416112;
   reg _416113_416113 ; 
   reg __416113_416113;
   reg _416114_416114 ; 
   reg __416114_416114;
   reg _416115_416115 ; 
   reg __416115_416115;
   reg _416116_416116 ; 
   reg __416116_416116;
   reg _416117_416117 ; 
   reg __416117_416117;
   reg _416118_416118 ; 
   reg __416118_416118;
   reg _416119_416119 ; 
   reg __416119_416119;
   reg _416120_416120 ; 
   reg __416120_416120;
   reg _416121_416121 ; 
   reg __416121_416121;
   reg _416122_416122 ; 
   reg __416122_416122;
   reg _416123_416123 ; 
   reg __416123_416123;
   reg _416124_416124 ; 
   reg __416124_416124;
   reg _416125_416125 ; 
   reg __416125_416125;
   reg _416126_416126 ; 
   reg __416126_416126;
   reg _416127_416127 ; 
   reg __416127_416127;
   reg _416128_416128 ; 
   reg __416128_416128;
   reg _416129_416129 ; 
   reg __416129_416129;
   reg _416130_416130 ; 
   reg __416130_416130;
   reg _416131_416131 ; 
   reg __416131_416131;
   reg _416132_416132 ; 
   reg __416132_416132;
   reg _416133_416133 ; 
   reg __416133_416133;
   reg _416134_416134 ; 
   reg __416134_416134;
   reg _416135_416135 ; 
   reg __416135_416135;
   reg _416136_416136 ; 
   reg __416136_416136;
   reg _416137_416137 ; 
   reg __416137_416137;
   reg _416138_416138 ; 
   reg __416138_416138;
   reg _416139_416139 ; 
   reg __416139_416139;
   reg _416140_416140 ; 
   reg __416140_416140;
   reg _416141_416141 ; 
   reg __416141_416141;
   reg _416142_416142 ; 
   reg __416142_416142;
   reg _416143_416143 ; 
   reg __416143_416143;
   reg _416144_416144 ; 
   reg __416144_416144;
   reg _416145_416145 ; 
   reg __416145_416145;
   reg _416146_416146 ; 
   reg __416146_416146;
   reg _416147_416147 ; 
   reg __416147_416147;
   reg _416148_416148 ; 
   reg __416148_416148;
   reg _416149_416149 ; 
   reg __416149_416149;
   reg _416150_416150 ; 
   reg __416150_416150;
   reg _416151_416151 ; 
   reg __416151_416151;
   reg _416152_416152 ; 
   reg __416152_416152;
   reg _416153_416153 ; 
   reg __416153_416153;
   reg _416154_416154 ; 
   reg __416154_416154;
   reg _416155_416155 ; 
   reg __416155_416155;
   reg _416156_416156 ; 
   reg __416156_416156;
   reg _416157_416157 ; 
   reg __416157_416157;
   reg _416158_416158 ; 
   reg __416158_416158;
   reg _416159_416159 ; 
   reg __416159_416159;
   reg _416160_416160 ; 
   reg __416160_416160;
   reg _416161_416161 ; 
   reg __416161_416161;
   reg _416162_416162 ; 
   reg __416162_416162;
   reg _416163_416163 ; 
   reg __416163_416163;
   reg _416164_416164 ; 
   reg __416164_416164;
   reg _416165_416165 ; 
   reg __416165_416165;
   reg _416166_416166 ; 
   reg __416166_416166;
   reg _416167_416167 ; 
   reg __416167_416167;
   reg _416168_416168 ; 
   reg __416168_416168;
   reg _416169_416169 ; 
   reg __416169_416169;
   reg _416170_416170 ; 
   reg __416170_416170;
   reg _416171_416171 ; 
   reg __416171_416171;
   reg _416172_416172 ; 
   reg __416172_416172;
   reg _416173_416173 ; 
   reg __416173_416173;
   reg _416174_416174 ; 
   reg __416174_416174;
   reg _416175_416175 ; 
   reg __416175_416175;
   reg _416176_416176 ; 
   reg __416176_416176;
   reg _416177_416177 ; 
   reg __416177_416177;
   reg _416178_416178 ; 
   reg __416178_416178;
   reg _416179_416179 ; 
   reg __416179_416179;
   reg _416180_416180 ; 
   reg __416180_416180;
   reg _416181_416181 ; 
   reg __416181_416181;
   reg _416182_416182 ; 
   reg __416182_416182;
   reg _416183_416183 ; 
   reg __416183_416183;
   reg _416184_416184 ; 
   reg __416184_416184;
   reg _416185_416185 ; 
   reg __416185_416185;
   reg _416186_416186 ; 
   reg __416186_416186;
   reg _416187_416187 ; 
   reg __416187_416187;
   reg _416188_416188 ; 
   reg __416188_416188;
   reg _416189_416189 ; 
   reg __416189_416189;
   reg _416190_416190 ; 
   reg __416190_416190;
   reg _416191_416191 ; 
   reg __416191_416191;
   reg _416192_416192 ; 
   reg __416192_416192;
   reg _416193_416193 ; 
   reg __416193_416193;
   reg _416194_416194 ; 
   reg __416194_416194;
   reg _416195_416195 ; 
   reg __416195_416195;
   reg _416196_416196 ; 
   reg __416196_416196;
   reg _416197_416197 ; 
   reg __416197_416197;
   reg _416198_416198 ; 
   reg __416198_416198;
   reg _416199_416199 ; 
   reg __416199_416199;
   reg _416200_416200 ; 
   reg __416200_416200;
   reg _416201_416201 ; 
   reg __416201_416201;
   reg _416202_416202 ; 
   reg __416202_416202;
   reg _416203_416203 ; 
   reg __416203_416203;
   reg _416204_416204 ; 
   reg __416204_416204;
   reg _416205_416205 ; 
   reg __416205_416205;
   reg _416206_416206 ; 
   reg __416206_416206;
   reg _416207_416207 ; 
   reg __416207_416207;
   reg _416208_416208 ; 
   reg __416208_416208;
   reg _416209_416209 ; 
   reg __416209_416209;
   reg _416210_416210 ; 
   reg __416210_416210;
   reg _416211_416211 ; 
   reg __416211_416211;
   reg _416212_416212 ; 
   reg __416212_416212;
   reg _416213_416213 ; 
   reg __416213_416213;
   reg _416214_416214 ; 
   reg __416214_416214;
   reg _416215_416215 ; 
   reg __416215_416215;
   reg _416216_416216 ; 
   reg __416216_416216;
   reg _416217_416217 ; 
   reg __416217_416217;
   reg _416218_416218 ; 
   reg __416218_416218;
   reg _416219_416219 ; 
   reg __416219_416219;
   reg _416220_416220 ; 
   reg __416220_416220;
   reg _416221_416221 ; 
   reg __416221_416221;
   reg _416222_416222 ; 
   reg __416222_416222;
   reg _416223_416223 ; 
   reg __416223_416223;
   reg _416224_416224 ; 
   reg __416224_416224;
   reg _416225_416225 ; 
   reg __416225_416225;
   reg _416226_416226 ; 
   reg __416226_416226;
   reg _416227_416227 ; 
   reg __416227_416227;
   reg _416228_416228 ; 
   reg __416228_416228;
   reg _416229_416229 ; 
   reg __416229_416229;
   reg _416230_416230 ; 
   reg __416230_416230;
   reg _416231_416231 ; 
   reg __416231_416231;
   reg _416232_416232 ; 
   reg __416232_416232;
   reg _416233_416233 ; 
   reg __416233_416233;
   reg _416234_416234 ; 
   reg __416234_416234;
   reg _416235_416235 ; 
   reg __416235_416235;
   reg _416236_416236 ; 
   reg __416236_416236;
   reg _416237_416237 ; 
   reg __416237_416237;
   reg _416238_416238 ; 
   reg __416238_416238;
   reg _416239_416239 ; 
   reg __416239_416239;
   reg _416240_416240 ; 
   reg __416240_416240;
   reg _416241_416241 ; 
   reg __416241_416241;
   reg _416242_416242 ; 
   reg __416242_416242;
   reg _416243_416243 ; 
   reg __416243_416243;
   reg _416244_416244 ; 
   reg __416244_416244;
   reg _416245_416245 ; 
   reg __416245_416245;
   reg _416246_416246 ; 
   reg __416246_416246;
   reg _416247_416247 ; 
   reg __416247_416247;
   reg _416248_416248 ; 
   reg __416248_416248;
   reg _416249_416249 ; 
   reg __416249_416249;
   reg _416250_416250 ; 
   reg __416250_416250;
   reg _416251_416251 ; 
   reg __416251_416251;
   reg _416252_416252 ; 
   reg __416252_416252;
   reg _416253_416253 ; 
   reg __416253_416253;
   reg _416254_416254 ; 
   reg __416254_416254;
   reg _416255_416255 ; 
   reg __416255_416255;
   reg _416256_416256 ; 
   reg __416256_416256;
   reg _416257_416257 ; 
   reg __416257_416257;
   reg _416258_416258 ; 
   reg __416258_416258;
   reg _416259_416259 ; 
   reg __416259_416259;
   reg _416260_416260 ; 
   reg __416260_416260;
   reg _416261_416261 ; 
   reg __416261_416261;
   reg _416262_416262 ; 
   reg __416262_416262;
   reg _416263_416263 ; 
   reg __416263_416263;
   reg _416264_416264 ; 
   reg __416264_416264;
   reg _416265_416265 ; 
   reg __416265_416265;
   reg _416266_416266 ; 
   reg __416266_416266;
   reg _416267_416267 ; 
   reg __416267_416267;
   reg _416268_416268 ; 
   reg __416268_416268;
   reg _416269_416269 ; 
   reg __416269_416269;
   reg _416270_416270 ; 
   reg __416270_416270;
   reg _416271_416271 ; 
   reg __416271_416271;
   reg _416272_416272 ; 
   reg __416272_416272;
   reg _416273_416273 ; 
   reg __416273_416273;
   reg _416274_416274 ; 
   reg __416274_416274;
   reg _416275_416275 ; 
   reg __416275_416275;
   reg _416276_416276 ; 
   reg __416276_416276;
   reg _416277_416277 ; 
   reg __416277_416277;
   reg _416278_416278 ; 
   reg __416278_416278;
   reg _416279_416279 ; 
   reg __416279_416279;
   reg _416280_416280 ; 
   reg __416280_416280;
   reg _416281_416281 ; 
   reg __416281_416281;
   reg _416282_416282 ; 
   reg __416282_416282;
   reg _416283_416283 ; 
   reg __416283_416283;
   reg _416284_416284 ; 
   reg __416284_416284;
   reg _416285_416285 ; 
   reg __416285_416285;
   reg _416286_416286 ; 
   reg __416286_416286;
   reg _416287_416287 ; 
   reg __416287_416287;
   reg _416288_416288 ; 
   reg __416288_416288;
   reg _416289_416289 ; 
   reg __416289_416289;
   reg _416290_416290 ; 
   reg __416290_416290;
   reg _416291_416291 ; 
   reg __416291_416291;
   reg _416292_416292 ; 
   reg __416292_416292;
   reg _416293_416293 ; 
   reg __416293_416293;
   reg _416294_416294 ; 
   reg __416294_416294;
   reg _416295_416295 ; 
   reg __416295_416295;
   reg _416296_416296 ; 
   reg __416296_416296;
   reg _416297_416297 ; 
   reg __416297_416297;
   reg _416298_416298 ; 
   reg __416298_416298;
   reg _416299_416299 ; 
   reg __416299_416299;
   reg _416300_416300 ; 
   reg __416300_416300;
   reg _416301_416301 ; 
   reg __416301_416301;
   reg _416302_416302 ; 
   reg __416302_416302;
   reg _416303_416303 ; 
   reg __416303_416303;
   reg _416304_416304 ; 
   reg __416304_416304;
   reg _416305_416305 ; 
   reg __416305_416305;
   reg _416306_416306 ; 
   reg __416306_416306;
   reg _416307_416307 ; 
   reg __416307_416307;
   reg _416308_416308 ; 
   reg __416308_416308;
   reg _416309_416309 ; 
   reg __416309_416309;
   reg _416310_416310 ; 
   reg __416310_416310;
   reg _416311_416311 ; 
   reg __416311_416311;
   reg _416312_416312 ; 
   reg __416312_416312;
   reg _416313_416313 ; 
   reg __416313_416313;
   reg _416314_416314 ; 
   reg __416314_416314;
   reg _416315_416315 ; 
   reg __416315_416315;
   reg _416316_416316 ; 
   reg __416316_416316;
   reg _416317_416317 ; 
   reg __416317_416317;
   reg _416318_416318 ; 
   reg __416318_416318;
   reg _416319_416319 ; 
   reg __416319_416319;
   reg _416320_416320 ; 
   reg __416320_416320;
   reg _416321_416321 ; 
   reg __416321_416321;
   reg _416322_416322 ; 
   reg __416322_416322;
   reg _416323_416323 ; 
   reg __416323_416323;
   reg _416324_416324 ; 
   reg __416324_416324;
   reg _416325_416325 ; 
   reg __416325_416325;
   reg _416326_416326 ; 
   reg __416326_416326;
   reg _416327_416327 ; 
   reg __416327_416327;
   reg _416328_416328 ; 
   reg __416328_416328;
   reg _416329_416329 ; 
   reg __416329_416329;
   reg _416330_416330 ; 
   reg __416330_416330;
   reg _416331_416331 ; 
   reg __416331_416331;
   reg _416332_416332 ; 
   reg __416332_416332;
   reg _416333_416333 ; 
   reg __416333_416333;
   reg _416334_416334 ; 
   reg __416334_416334;
   reg _416335_416335 ; 
   reg __416335_416335;
   reg _416336_416336 ; 
   reg __416336_416336;
   reg _416337_416337 ; 
   reg __416337_416337;
   reg _416338_416338 ; 
   reg __416338_416338;
   reg _416339_416339 ; 
   reg __416339_416339;
   reg _416340_416340 ; 
   reg __416340_416340;
   reg _416341_416341 ; 
   reg __416341_416341;
   reg _416342_416342 ; 
   reg __416342_416342;
   reg _416343_416343 ; 
   reg __416343_416343;
   reg _416344_416344 ; 
   reg __416344_416344;
   reg _416345_416345 ; 
   reg __416345_416345;
   reg _416346_416346 ; 
   reg __416346_416346;
   reg _416347_416347 ; 
   reg __416347_416347;
   reg _416348_416348 ; 
   reg __416348_416348;
   reg _416349_416349 ; 
   reg __416349_416349;
   reg _416350_416350 ; 
   reg __416350_416350;
   reg _416351_416351 ; 
   reg __416351_416351;
   reg _416352_416352 ; 
   reg __416352_416352;
   reg _416353_416353 ; 
   reg __416353_416353;
   reg _416354_416354 ; 
   reg __416354_416354;
   reg _416355_416355 ; 
   reg __416355_416355;
   reg _416356_416356 ; 
   reg __416356_416356;
   reg _416357_416357 ; 
   reg __416357_416357;
   reg _416358_416358 ; 
   reg __416358_416358;
   reg _416359_416359 ; 
   reg __416359_416359;
   reg _416360_416360 ; 
   reg __416360_416360;
   reg _416361_416361 ; 
   reg __416361_416361;
   reg _416362_416362 ; 
   reg __416362_416362;
   reg _416363_416363 ; 
   reg __416363_416363;
   reg _416364_416364 ; 
   reg __416364_416364;
   reg _416365_416365 ; 
   reg __416365_416365;
   reg _416366_416366 ; 
   reg __416366_416366;
   reg _416367_416367 ; 
   reg __416367_416367;
   reg _416368_416368 ; 
   reg __416368_416368;
   reg _416369_416369 ; 
   reg __416369_416369;
   reg _416370_416370 ; 
   reg __416370_416370;
   reg _416371_416371 ; 
   reg __416371_416371;
   reg _416372_416372 ; 
   reg __416372_416372;
   reg _416373_416373 ; 
   reg __416373_416373;
   reg _416374_416374 ; 
   reg __416374_416374;
   reg _416375_416375 ; 
   reg __416375_416375;
   reg _416376_416376 ; 
   reg __416376_416376;
   reg _416377_416377 ; 
   reg __416377_416377;
   reg _416378_416378 ; 
   reg __416378_416378;
   reg _416379_416379 ; 
   reg __416379_416379;
   reg _416380_416380 ; 
   reg __416380_416380;
   reg _416381_416381 ; 
   reg __416381_416381;
   reg _416382_416382 ; 
   reg __416382_416382;
   reg _416383_416383 ; 
   reg __416383_416383;
   reg _416384_416384 ; 
   reg __416384_416384;
   reg _416385_416385 ; 
   reg __416385_416385;
   reg _416386_416386 ; 
   reg __416386_416386;
   reg _416387_416387 ; 
   reg __416387_416387;
   reg _416388_416388 ; 
   reg __416388_416388;
   reg _416389_416389 ; 
   reg __416389_416389;
   reg _416390_416390 ; 
   reg __416390_416390;
   reg _416391_416391 ; 
   reg __416391_416391;
   reg _416392_416392 ; 
   reg __416392_416392;
   reg _416393_416393 ; 
   reg __416393_416393;
   reg _416394_416394 ; 
   reg __416394_416394;
   reg _416395_416395 ; 
   reg __416395_416395;
   reg _416396_416396 ; 
   reg __416396_416396;
   reg _416397_416397 ; 
   reg __416397_416397;
   reg _416398_416398 ; 
   reg __416398_416398;
   reg _416399_416399 ; 
   reg __416399_416399;
   reg _416400_416400 ; 
   reg __416400_416400;
   reg _416401_416401 ; 
   reg __416401_416401;
   reg _416402_416402 ; 
   reg __416402_416402;
   reg _416403_416403 ; 
   reg __416403_416403;
   reg _416404_416404 ; 
   reg __416404_416404;
   reg _416405_416405 ; 
   reg __416405_416405;
   reg _416406_416406 ; 
   reg __416406_416406;
   reg _416407_416407 ; 
   reg __416407_416407;
   reg _416408_416408 ; 
   reg __416408_416408;
   reg _416409_416409 ; 
   reg __416409_416409;
   reg _416410_416410 ; 
   reg __416410_416410;
   reg _416411_416411 ; 
   reg __416411_416411;
   reg _416412_416412 ; 
   reg __416412_416412;
   reg _416413_416413 ; 
   reg __416413_416413;
   reg _416414_416414 ; 
   reg __416414_416414;
   reg _416415_416415 ; 
   reg __416415_416415;
   reg _416416_416416 ; 
   reg __416416_416416;
   reg _416417_416417 ; 
   reg __416417_416417;
   reg _416418_416418 ; 
   reg __416418_416418;
   reg _416419_416419 ; 
   reg __416419_416419;
   reg _416420_416420 ; 
   reg __416420_416420;
   reg _416421_416421 ; 
   reg __416421_416421;
   reg _416422_416422 ; 
   reg __416422_416422;
   reg _416423_416423 ; 
   reg __416423_416423;
   reg _416424_416424 ; 
   reg __416424_416424;
   reg _416425_416425 ; 
   reg __416425_416425;
   reg _416426_416426 ; 
   reg __416426_416426;
   reg _416427_416427 ; 
   reg __416427_416427;
   reg _416428_416428 ; 
   reg __416428_416428;
   reg _416429_416429 ; 
   reg __416429_416429;
   reg _416430_416430 ; 
   reg __416430_416430;
   reg _416431_416431 ; 
   reg __416431_416431;
   reg _416432_416432 ; 
   reg __416432_416432;
   reg _416433_416433 ; 
   reg __416433_416433;
   reg _416434_416434 ; 
   reg __416434_416434;
   reg _416435_416435 ; 
   reg __416435_416435;
   reg _416436_416436 ; 
   reg __416436_416436;
   reg _416437_416437 ; 
   reg __416437_416437;
   reg _416438_416438 ; 
   reg __416438_416438;
   reg _416439_416439 ; 
   reg __416439_416439;
   reg _416440_416440 ; 
   reg __416440_416440;
   reg _416441_416441 ; 
   reg __416441_416441;
   reg _416442_416442 ; 
   reg __416442_416442;
   reg _416443_416443 ; 
   reg __416443_416443;
   reg _416444_416444 ; 
   reg __416444_416444;
   reg _416445_416445 ; 
   reg __416445_416445;
   reg _416446_416446 ; 
   reg __416446_416446;
   reg _416447_416447 ; 
   reg __416447_416447;
   reg _416448_416448 ; 
   reg __416448_416448;
   reg _416449_416449 ; 
   reg __416449_416449;
   reg _416450_416450 ; 
   reg __416450_416450;
   reg _416451_416451 ; 
   reg __416451_416451;
   reg _416452_416452 ; 
   reg __416452_416452;
   reg _416453_416453 ; 
   reg __416453_416453;
   reg _416454_416454 ; 
   reg __416454_416454;
   reg _416455_416455 ; 
   reg __416455_416455;
   reg _416456_416456 ; 
   reg __416456_416456;
   reg _416457_416457 ; 
   reg __416457_416457;
   reg _416458_416458 ; 
   reg __416458_416458;
   reg _416459_416459 ; 
   reg __416459_416459;
   reg _416460_416460 ; 
   reg __416460_416460;
   reg _416461_416461 ; 
   reg __416461_416461;
   reg _416462_416462 ; 
   reg __416462_416462;
   reg _416463_416463 ; 
   reg __416463_416463;
   reg _416464_416464 ; 
   reg __416464_416464;
   reg _416465_416465 ; 
   reg __416465_416465;
   reg _416466_416466 ; 
   reg __416466_416466;
   reg _416467_416467 ; 
   reg __416467_416467;
   reg _416468_416468 ; 
   reg __416468_416468;
   reg _416469_416469 ; 
   reg __416469_416469;
   reg _416470_416470 ; 
   reg __416470_416470;
   reg _416471_416471 ; 
   reg __416471_416471;
   reg _416472_416472 ; 
   reg __416472_416472;
   reg _416473_416473 ; 
   reg __416473_416473;
   reg _416474_416474 ; 
   reg __416474_416474;
   reg _416475_416475 ; 
   reg __416475_416475;
   reg _416476_416476 ; 
   reg __416476_416476;
   reg _416477_416477 ; 
   reg __416477_416477;
   reg _416478_416478 ; 
   reg __416478_416478;
   reg _416479_416479 ; 
   reg __416479_416479;
   reg _416480_416480 ; 
   reg __416480_416480;
   reg _416481_416481 ; 
   reg __416481_416481;
   reg _416482_416482 ; 
   reg __416482_416482;
   reg _416483_416483 ; 
   reg __416483_416483;
   reg _416484_416484 ; 
   reg __416484_416484;
   reg _416485_416485 ; 
   reg __416485_416485;
   reg _416486_416486 ; 
   reg __416486_416486;
   reg _416487_416487 ; 
   reg __416487_416487;
   reg _416488_416488 ; 
   reg __416488_416488;
   reg _416489_416489 ; 
   reg __416489_416489;
   reg _416490_416490 ; 
   reg __416490_416490;
   reg _416491_416491 ; 
   reg __416491_416491;
   reg _416492_416492 ; 
   reg __416492_416492;
   reg _416493_416493 ; 
   reg __416493_416493;
   reg _416494_416494 ; 
   reg __416494_416494;
   reg _416495_416495 ; 
   reg __416495_416495;
   reg _416496_416496 ; 
   reg __416496_416496;
   reg _416497_416497 ; 
   reg __416497_416497;
   reg _416498_416498 ; 
   reg __416498_416498;
   reg _416499_416499 ; 
   reg __416499_416499;
   reg _416500_416500 ; 
   reg __416500_416500;
   reg _416501_416501 ; 
   reg __416501_416501;
   reg _416502_416502 ; 
   reg __416502_416502;
   reg _416503_416503 ; 
   reg __416503_416503;
   reg _416504_416504 ; 
   reg __416504_416504;
   reg _416505_416505 ; 
   reg __416505_416505;
   reg _416506_416506 ; 
   reg __416506_416506;
   reg _416507_416507 ; 
   reg __416507_416507;
   reg _416508_416508 ; 
   reg __416508_416508;
   reg _416509_416509 ; 
   reg __416509_416509;
   reg _416510_416510 ; 
   reg __416510_416510;
   reg _416511_416511 ; 
   reg __416511_416511;
   reg _416512_416512 ; 
   reg __416512_416512;
   reg _416513_416513 ; 
   reg __416513_416513;
   reg _416514_416514 ; 
   reg __416514_416514;
   reg _416515_416515 ; 
   reg __416515_416515;
   reg _416516_416516 ; 
   reg __416516_416516;
   reg _416517_416517 ; 
   reg __416517_416517;
   reg _416518_416518 ; 
   reg __416518_416518;
   reg _416519_416519 ; 
   reg __416519_416519;
   reg _416520_416520 ; 
   reg __416520_416520;
   reg _416521_416521 ; 
   reg __416521_416521;
   reg _416522_416522 ; 
   reg __416522_416522;
   reg _416523_416523 ; 
   reg __416523_416523;
   reg _416524_416524 ; 
   reg __416524_416524;
   reg _416525_416525 ; 
   reg __416525_416525;
   reg _416526_416526 ; 
   reg __416526_416526;
   reg _416527_416527 ; 
   reg __416527_416527;
   reg _416528_416528 ; 
   reg __416528_416528;
   reg _416529_416529 ; 
   reg __416529_416529;
   reg _416530_416530 ; 
   reg __416530_416530;
   reg _416531_416531 ; 
   reg __416531_416531;
   reg _416532_416532 ; 
   reg __416532_416532;
   reg _416533_416533 ; 
   reg __416533_416533;
   reg _416534_416534 ; 
   reg __416534_416534;
   reg _416535_416535 ; 
   reg __416535_416535;
   reg _416536_416536 ; 
   reg __416536_416536;
   reg _416537_416537 ; 
   reg __416537_416537;
   reg _416538_416538 ; 
   reg __416538_416538;
   reg _416539_416539 ; 
   reg __416539_416539;
   reg _416540_416540 ; 
   reg __416540_416540;
   reg _416541_416541 ; 
   reg __416541_416541;
   reg _416542_416542 ; 
   reg __416542_416542;
   reg _416543_416543 ; 
   reg __416543_416543;
   reg _416544_416544 ; 
   reg __416544_416544;
   reg _416545_416545 ; 
   reg __416545_416545;
   reg _416546_416546 ; 
   reg __416546_416546;
   reg _416547_416547 ; 
   reg __416547_416547;
   reg _416548_416548 ; 
   reg __416548_416548;
   reg _416549_416549 ; 
   reg __416549_416549;
   reg _416550_416550 ; 
   reg __416550_416550;
   reg _416551_416551 ; 
   reg __416551_416551;
   reg _416552_416552 ; 
   reg __416552_416552;
   reg _416553_416553 ; 
   reg __416553_416553;
   reg _416554_416554 ; 
   reg __416554_416554;
   reg _416555_416555 ; 
   reg __416555_416555;
   reg _416556_416556 ; 
   reg __416556_416556;
   reg _416557_416557 ; 
   reg __416557_416557;
   reg _416558_416558 ; 
   reg __416558_416558;
   reg _416559_416559 ; 
   reg __416559_416559;
   reg _416560_416560 ; 
   reg __416560_416560;
   reg _416561_416561 ; 
   reg __416561_416561;
   reg _416562_416562 ; 
   reg __416562_416562;
   reg _416563_416563 ; 
   reg __416563_416563;
   reg _416564_416564 ; 
   reg __416564_416564;
   reg _416565_416565 ; 
   reg __416565_416565;
   reg _416566_416566 ; 
   reg __416566_416566;
   reg _416567_416567 ; 
   reg __416567_416567;
   reg _416568_416568 ; 
   reg __416568_416568;
   reg _416569_416569 ; 
   reg __416569_416569;
   reg _416570_416570 ; 
   reg __416570_416570;
   reg _416571_416571 ; 
   reg __416571_416571;
   reg _416572_416572 ; 
   reg __416572_416572;
   reg _416573_416573 ; 
   reg __416573_416573;
   reg _416574_416574 ; 
   reg __416574_416574;
   reg _416575_416575 ; 
   reg __416575_416575;
   reg _416576_416576 ; 
   reg __416576_416576;
   reg _416577_416577 ; 
   reg __416577_416577;
   reg _416578_416578 ; 
   reg __416578_416578;
   reg _416579_416579 ; 
   reg __416579_416579;
   reg _416580_416580 ; 
   reg __416580_416580;
   reg _416581_416581 ; 
   reg __416581_416581;
   reg _416582_416582 ; 
   reg __416582_416582;
   reg _416583_416583 ; 
   reg __416583_416583;
   reg _416584_416584 ; 
   reg __416584_416584;
   reg _416585_416585 ; 
   reg __416585_416585;
   reg _416586_416586 ; 
   reg __416586_416586;
   reg _416587_416587 ; 
   reg __416587_416587;
   reg _416588_416588 ; 
   reg __416588_416588;
   reg _416589_416589 ; 
   reg __416589_416589;
   reg _416590_416590 ; 
   reg __416590_416590;
   reg _416591_416591 ; 
   reg __416591_416591;
   reg _416592_416592 ; 
   reg __416592_416592;
   reg _416593_416593 ; 
   reg __416593_416593;
   reg _416594_416594 ; 
   reg __416594_416594;
   reg _416595_416595 ; 
   reg __416595_416595;
   reg _416596_416596 ; 
   reg __416596_416596;
   reg _416597_416597 ; 
   reg __416597_416597;
   reg _416598_416598 ; 
   reg __416598_416598;
   reg _416599_416599 ; 
   reg __416599_416599;
   reg _416600_416600 ; 
   reg __416600_416600;
   reg _416601_416601 ; 
   reg __416601_416601;
   reg _416602_416602 ; 
   reg __416602_416602;
   reg _416603_416603 ; 
   reg __416603_416603;
   reg _416604_416604 ; 
   reg __416604_416604;
   reg _416605_416605 ; 
   reg __416605_416605;
   reg _416606_416606 ; 
   reg __416606_416606;
   reg _416607_416607 ; 
   reg __416607_416607;
   reg _416608_416608 ; 
   reg __416608_416608;
   reg _416609_416609 ; 
   reg __416609_416609;
   reg _416610_416610 ; 
   reg __416610_416610;
   reg _416611_416611 ; 
   reg __416611_416611;
   reg _416612_416612 ; 
   reg __416612_416612;
   reg _416613_416613 ; 
   reg __416613_416613;
   reg _416614_416614 ; 
   reg __416614_416614;
   reg _416615_416615 ; 
   reg __416615_416615;
   reg _416616_416616 ; 
   reg __416616_416616;
   reg _416617_416617 ; 
   reg __416617_416617;
   reg _416618_416618 ; 
   reg __416618_416618;
   reg _416619_416619 ; 
   reg __416619_416619;
   reg _416620_416620 ; 
   reg __416620_416620;
   reg _416621_416621 ; 
   reg __416621_416621;
   reg _416622_416622 ; 
   reg __416622_416622;
   reg _416623_416623 ; 
   reg __416623_416623;
   reg _416624_416624 ; 
   reg __416624_416624;
   reg _416625_416625 ; 
   reg __416625_416625;
   reg _416626_416626 ; 
   reg __416626_416626;
   reg _416627_416627 ; 
   reg __416627_416627;
   reg _416628_416628 ; 
   reg __416628_416628;
   reg _416629_416629 ; 
   reg __416629_416629;
   reg _416630_416630 ; 
   reg __416630_416630;
   reg _416631_416631 ; 
   reg __416631_416631;
   reg _416632_416632 ; 
   reg __416632_416632;
   reg _416633_416633 ; 
   reg __416633_416633;
   reg _416634_416634 ; 
   reg __416634_416634;
   reg _416635_416635 ; 
   reg __416635_416635;
   reg _416636_416636 ; 
   reg __416636_416636;
   reg _416637_416637 ; 
   reg __416637_416637;
   reg _416638_416638 ; 
   reg __416638_416638;
   reg _416639_416639 ; 
   reg __416639_416639;
   reg _416640_416640 ; 
   reg __416640_416640;
   reg _416641_416641 ; 
   reg __416641_416641;
   reg _416642_416642 ; 
   reg __416642_416642;
   reg _416643_416643 ; 
   reg __416643_416643;
   reg _416644_416644 ; 
   reg __416644_416644;
   reg _416645_416645 ; 
   reg __416645_416645;
   reg _416646_416646 ; 
   reg __416646_416646;
   reg _416647_416647 ; 
   reg __416647_416647;
   reg _416648_416648 ; 
   reg __416648_416648;
   reg _416649_416649 ; 
   reg __416649_416649;
   reg _416650_416650 ; 
   reg __416650_416650;
   reg _416651_416651 ; 
   reg __416651_416651;
   reg _416652_416652 ; 
   reg __416652_416652;
   reg _416653_416653 ; 
   reg __416653_416653;
   reg _416654_416654 ; 
   reg __416654_416654;
   reg _416655_416655 ; 
   reg __416655_416655;
   reg _416656_416656 ; 
   reg __416656_416656;
   reg _416657_416657 ; 
   reg __416657_416657;
   reg _416658_416658 ; 
   reg __416658_416658;
   reg _416659_416659 ; 
   reg __416659_416659;
   reg _416660_416660 ; 
   reg __416660_416660;
   reg _416661_416661 ; 
   reg __416661_416661;
   reg _416662_416662 ; 
   reg __416662_416662;
   reg _416663_416663 ; 
   reg __416663_416663;
   reg _416664_416664 ; 
   reg __416664_416664;
   reg _416665_416665 ; 
   reg __416665_416665;
   reg _416666_416666 ; 
   reg __416666_416666;
   reg _416667_416667 ; 
   reg __416667_416667;
   reg _416668_416668 ; 
   reg __416668_416668;
   reg _416669_416669 ; 
   reg __416669_416669;
   reg _416670_416670 ; 
   reg __416670_416670;
   reg _416671_416671 ; 
   reg __416671_416671;
   reg _416672_416672 ; 
   reg __416672_416672;
   reg _416673_416673 ; 
   reg __416673_416673;
   reg _416674_416674 ; 
   reg __416674_416674;
   reg _416675_416675 ; 
   reg __416675_416675;
   reg _416676_416676 ; 
   reg __416676_416676;
   reg _416677_416677 ; 
   reg __416677_416677;
   reg _416678_416678 ; 
   reg __416678_416678;
   reg _416679_416679 ; 
   reg __416679_416679;
   reg _416680_416680 ; 
   reg __416680_416680;
   reg _416681_416681 ; 
   reg __416681_416681;
   reg _416682_416682 ; 
   reg __416682_416682;
   reg _416683_416683 ; 
   reg __416683_416683;
   reg _416684_416684 ; 
   reg __416684_416684;
   reg _416685_416685 ; 
   reg __416685_416685;
   reg _416686_416686 ; 
   reg __416686_416686;
   reg _416687_416687 ; 
   reg __416687_416687;
   reg _416688_416688 ; 
   reg __416688_416688;
   reg _416689_416689 ; 
   reg __416689_416689;
   reg _416690_416690 ; 
   reg __416690_416690;
   reg _416691_416691 ; 
   reg __416691_416691;
   reg _416692_416692 ; 
   reg __416692_416692;
   reg _416693_416693 ; 
   reg __416693_416693;
   reg _416694_416694 ; 
   reg __416694_416694;
   reg _416695_416695 ; 
   reg __416695_416695;
   reg _416696_416696 ; 
   reg __416696_416696;
   reg _416697_416697 ; 
   reg __416697_416697;
   reg _416698_416698 ; 
   reg __416698_416698;
   reg _416699_416699 ; 
   reg __416699_416699;
   reg _416700_416700 ; 
   reg __416700_416700;
   reg _416701_416701 ; 
   reg __416701_416701;
   reg _416702_416702 ; 
   reg __416702_416702;
   reg _416703_416703 ; 
   reg __416703_416703;
   reg _416704_416704 ; 
   reg __416704_416704;
   reg _416705_416705 ; 
   reg __416705_416705;
   reg _416706_416706 ; 
   reg __416706_416706;
   reg _416707_416707 ; 
   reg __416707_416707;
   reg _416708_416708 ; 
   reg __416708_416708;
   reg _416709_416709 ; 
   reg __416709_416709;
   reg _416710_416710 ; 
   reg __416710_416710;
   reg _416711_416711 ; 
   reg __416711_416711;
   reg _416712_416712 ; 
   reg __416712_416712;
   reg _416713_416713 ; 
   reg __416713_416713;
   reg _416714_416714 ; 
   reg __416714_416714;
   reg _416715_416715 ; 
   reg __416715_416715;
   reg _416716_416716 ; 
   reg __416716_416716;
   reg _416717_416717 ; 
   reg __416717_416717;
   reg _416718_416718 ; 
   reg __416718_416718;
   reg _416719_416719 ; 
   reg __416719_416719;
   reg _416720_416720 ; 
   reg __416720_416720;
   reg _416721_416721 ; 
   reg __416721_416721;
   reg _416722_416722 ; 
   reg __416722_416722;
   reg _416723_416723 ; 
   reg __416723_416723;
   reg _416724_416724 ; 
   reg __416724_416724;
   reg _416725_416725 ; 
   reg __416725_416725;
   reg _416726_416726 ; 
   reg __416726_416726;
   reg _416727_416727 ; 
   reg __416727_416727;
   reg _416728_416728 ; 
   reg __416728_416728;
   reg _416729_416729 ; 
   reg __416729_416729;
   reg _416730_416730 ; 
   reg __416730_416730;
   reg _416731_416731 ; 
   reg __416731_416731;
   reg _416732_416732 ; 
   reg __416732_416732;
   reg _416733_416733 ; 
   reg __416733_416733;
   reg _416734_416734 ; 
   reg __416734_416734;
   reg _416735_416735 ; 
   reg __416735_416735;
   reg _416736_416736 ; 
   reg __416736_416736;
   reg _416737_416737 ; 
   reg __416737_416737;
   reg _416738_416738 ; 
   reg __416738_416738;
   reg _416739_416739 ; 
   reg __416739_416739;
   reg _416740_416740 ; 
   reg __416740_416740;
   reg _416741_416741 ; 
   reg __416741_416741;
   reg _416742_416742 ; 
   reg __416742_416742;
   reg _416743_416743 ; 
   reg __416743_416743;
   reg _416744_416744 ; 
   reg __416744_416744;
   reg _416745_416745 ; 
   reg __416745_416745;
   reg _416746_416746 ; 
   reg __416746_416746;
   reg _416747_416747 ; 
   reg __416747_416747;
   reg _416748_416748 ; 
   reg __416748_416748;
   reg _416749_416749 ; 
   reg __416749_416749;
   reg _416750_416750 ; 
   reg __416750_416750;
   reg _416751_416751 ; 
   reg __416751_416751;
   reg _416752_416752 ; 
   reg __416752_416752;
   reg _416753_416753 ; 
   reg __416753_416753;
   reg _416754_416754 ; 
   reg __416754_416754;
   reg _416755_416755 ; 
   reg __416755_416755;
   reg _416756_416756 ; 
   reg __416756_416756;
   reg _416757_416757 ; 
   reg __416757_416757;
   reg _416758_416758 ; 
   reg __416758_416758;
   reg _416759_416759 ; 
   reg __416759_416759;
   reg _416760_416760 ; 
   reg __416760_416760;
   reg _416761_416761 ; 
   reg __416761_416761;
   reg _416762_416762 ; 
   reg __416762_416762;
   reg _416763_416763 ; 
   reg __416763_416763;
   reg _416764_416764 ; 
   reg __416764_416764;
   reg _416765_416765 ; 
   reg __416765_416765;
   reg _416766_416766 ; 
   reg __416766_416766;
   reg _416767_416767 ; 
   reg __416767_416767;
   reg _416768_416768 ; 
   reg __416768_416768;
   reg _416769_416769 ; 
   reg __416769_416769;
   reg _416770_416770 ; 
   reg __416770_416770;
   reg _416771_416771 ; 
   reg __416771_416771;
   reg _416772_416772 ; 
   reg __416772_416772;
   reg _416773_416773 ; 
   reg __416773_416773;
   reg _416774_416774 ; 
   reg __416774_416774;
   reg _416775_416775 ; 
   reg __416775_416775;
   reg _416776_416776 ; 
   reg __416776_416776;
   reg _416777_416777 ; 
   reg __416777_416777;
   reg _416778_416778 ; 
   reg __416778_416778;
   reg _416779_416779 ; 
   reg __416779_416779;
   reg _416780_416780 ; 
   reg __416780_416780;
   reg _416781_416781 ; 
   reg __416781_416781;
   reg _416782_416782 ; 
   reg __416782_416782;
   reg _416783_416783 ; 
   reg __416783_416783;
   reg _416784_416784 ; 
   reg __416784_416784;
   reg _416785_416785 ; 
   reg __416785_416785;
   reg _416786_416786 ; 
   reg __416786_416786;
   reg _416787_416787 ; 
   reg __416787_416787;
   reg _416788_416788 ; 
   reg __416788_416788;
   reg _416789_416789 ; 
   reg __416789_416789;
   reg _416790_416790 ; 
   reg __416790_416790;
   reg _416791_416791 ; 
   reg __416791_416791;
   reg _416792_416792 ; 
   reg __416792_416792;
   reg _416793_416793 ; 
   reg __416793_416793;
   reg _416794_416794 ; 
   reg __416794_416794;
   reg _416795_416795 ; 
   reg __416795_416795;
   reg _416796_416796 ; 
   reg __416796_416796;
   reg _416797_416797 ; 
   reg __416797_416797;
   reg _416798_416798 ; 
   reg __416798_416798;
   reg _416799_416799 ; 
   reg __416799_416799;
   reg _416800_416800 ; 
   reg __416800_416800;
   reg _416801_416801 ; 
   reg __416801_416801;
   reg _416802_416802 ; 
   reg __416802_416802;
   reg _416803_416803 ; 
   reg __416803_416803;
   reg _416804_416804 ; 
   reg __416804_416804;
   reg _416805_416805 ; 
   reg __416805_416805;
   reg _416806_416806 ; 
   reg __416806_416806;
   reg _416807_416807 ; 
   reg __416807_416807;
   reg _416808_416808 ; 
   reg __416808_416808;
   reg _416809_416809 ; 
   reg __416809_416809;
   reg _416810_416810 ; 
   reg __416810_416810;
   reg _416811_416811 ; 
   reg __416811_416811;
   reg _416812_416812 ; 
   reg __416812_416812;
   reg _416813_416813 ; 
   reg __416813_416813;
   reg _416814_416814 ; 
   reg __416814_416814;
   reg _416815_416815 ; 
   reg __416815_416815;
   reg _416816_416816 ; 
   reg __416816_416816;
   reg _416817_416817 ; 
   reg __416817_416817;
   reg _416818_416818 ; 
   reg __416818_416818;
   reg _416819_416819 ; 
   reg __416819_416819;
   reg _416820_416820 ; 
   reg __416820_416820;
   reg _416821_416821 ; 
   reg __416821_416821;
   reg _416822_416822 ; 
   reg __416822_416822;
   reg _416823_416823 ; 
   reg __416823_416823;
   reg _416824_416824 ; 
   reg __416824_416824;
   reg _416825_416825 ; 
   reg __416825_416825;
   reg _416826_416826 ; 
   reg __416826_416826;
   reg _416827_416827 ; 
   reg __416827_416827;
   reg _416828_416828 ; 
   reg __416828_416828;
   reg _416829_416829 ; 
   reg __416829_416829;
   reg _416830_416830 ; 
   reg __416830_416830;
   reg _416831_416831 ; 
   reg __416831_416831;
   reg _416832_416832 ; 
   reg __416832_416832;
   reg _416833_416833 ; 
   reg __416833_416833;
   reg _416834_416834 ; 
   reg __416834_416834;
   reg _416835_416835 ; 
   reg __416835_416835;
   reg _416836_416836 ; 
   reg __416836_416836;
   reg _416837_416837 ; 
   reg __416837_416837;
   reg _416838_416838 ; 
   reg __416838_416838;
   reg _416839_416839 ; 
   reg __416839_416839;
   reg _416840_416840 ; 
   reg __416840_416840;
   reg _416841_416841 ; 
   reg __416841_416841;
   reg _416842_416842 ; 
   reg __416842_416842;
   reg _416843_416843 ; 
   reg __416843_416843;
   reg _416844_416844 ; 
   reg __416844_416844;
   reg _416845_416845 ; 
   reg __416845_416845;
   reg _416846_416846 ; 
   reg __416846_416846;
   reg _416847_416847 ; 
   reg __416847_416847;
   reg _416848_416848 ; 
   reg __416848_416848;
   reg _416849_416849 ; 
   reg __416849_416849;
   reg _416850_416850 ; 
   reg __416850_416850;
   reg _416851_416851 ; 
   reg __416851_416851;
   reg _416852_416852 ; 
   reg __416852_416852;
   reg _416853_416853 ; 
   reg __416853_416853;
   reg _416854_416854 ; 
   reg __416854_416854;
   reg _416855_416855 ; 
   reg __416855_416855;
   reg _416856_416856 ; 
   reg __416856_416856;
   reg _416857_416857 ; 
   reg __416857_416857;
   reg _416858_416858 ; 
   reg __416858_416858;
   reg _416859_416859 ; 
   reg __416859_416859;
   reg _416860_416860 ; 
   reg __416860_416860;
   reg _416861_416861 ; 
   reg __416861_416861;
   reg _416862_416862 ; 
   reg __416862_416862;
   reg _416863_416863 ; 
   reg __416863_416863;
   reg _416864_416864 ; 
   reg __416864_416864;
   reg _416865_416865 ; 
   reg __416865_416865;
   reg _416866_416866 ; 
   reg __416866_416866;
   reg _416867_416867 ; 
   reg __416867_416867;
   reg _416868_416868 ; 
   reg __416868_416868;
   reg _416869_416869 ; 
   reg __416869_416869;
   reg _416870_416870 ; 
   reg __416870_416870;
   reg _416871_416871 ; 
   reg __416871_416871;
   reg _416872_416872 ; 
   reg __416872_416872;
   reg _416873_416873 ; 
   reg __416873_416873;
   reg _416874_416874 ; 
   reg __416874_416874;
   reg _416875_416875 ; 
   reg __416875_416875;
   reg _416876_416876 ; 
   reg __416876_416876;
   reg _416877_416877 ; 
   reg __416877_416877;
   reg _416878_416878 ; 
   reg __416878_416878;
   reg _416879_416879 ; 
   reg __416879_416879;
   reg _416880_416880 ; 
   reg __416880_416880;
   reg _416881_416881 ; 
   reg __416881_416881;
   reg _416882_416882 ; 
   reg __416882_416882;
   reg _416883_416883 ; 
   reg __416883_416883;
   reg _416884_416884 ; 
   reg __416884_416884;
   reg _416885_416885 ; 
   reg __416885_416885;
   reg _416886_416886 ; 
   reg __416886_416886;
   reg _416887_416887 ; 
   reg __416887_416887;
   reg _416888_416888 ; 
   reg __416888_416888;
   reg _416889_416889 ; 
   reg __416889_416889;
   reg _416890_416890 ; 
   reg __416890_416890;
   reg _416891_416891 ; 
   reg __416891_416891;
   reg _416892_416892 ; 
   reg __416892_416892;
   reg _416893_416893 ; 
   reg __416893_416893;
   reg _416894_416894 ; 
   reg __416894_416894;
   reg _416895_416895 ; 
   reg __416895_416895;
   reg _416896_416896 ; 
   reg __416896_416896;
   reg _416897_416897 ; 
   reg __416897_416897;
   reg _416898_416898 ; 
   reg __416898_416898;
   reg _416899_416899 ; 
   reg __416899_416899;
   reg _416900_416900 ; 
   reg __416900_416900;
   reg _416901_416901 ; 
   reg __416901_416901;
   reg _416902_416902 ; 
   reg __416902_416902;
   reg _416903_416903 ; 
   reg __416903_416903;
   reg _416904_416904 ; 
   reg __416904_416904;
   reg _416905_416905 ; 
   reg __416905_416905;
   reg _416906_416906 ; 
   reg __416906_416906;
   reg _416907_416907 ; 
   reg __416907_416907;
   reg _416908_416908 ; 
   reg __416908_416908;
   reg _416909_416909 ; 
   reg __416909_416909;
   reg _416910_416910 ; 
   reg __416910_416910;
   reg _416911_416911 ; 
   reg __416911_416911;
   reg _416912_416912 ; 
   reg __416912_416912;
   reg _416913_416913 ; 
   reg __416913_416913;
   reg _416914_416914 ; 
   reg __416914_416914;
   reg _416915_416915 ; 
   reg __416915_416915;
   reg _416916_416916 ; 
   reg __416916_416916;
   reg _416917_416917 ; 
   reg __416917_416917;
   reg _416918_416918 ; 
   reg __416918_416918;
   reg _416919_416919 ; 
   reg __416919_416919;
   reg _416920_416920 ; 
   reg __416920_416920;
   reg _416921_416921 ; 
   reg __416921_416921;
   reg _416922_416922 ; 
   reg __416922_416922;
   reg _416923_416923 ; 
   reg __416923_416923;
   reg _416924_416924 ; 
   reg __416924_416924;
   reg _416925_416925 ; 
   reg __416925_416925;
   reg _416926_416926 ; 
   reg __416926_416926;
   reg _416927_416927 ; 
   reg __416927_416927;
   reg _416928_416928 ; 
   reg __416928_416928;
   reg _416929_416929 ; 
   reg __416929_416929;
   reg _416930_416930 ; 
   reg __416930_416930;
   reg _416931_416931 ; 
   reg __416931_416931;
   reg _416932_416932 ; 
   reg __416932_416932;
   reg _416933_416933 ; 
   reg __416933_416933;
   reg _416934_416934 ; 
   reg __416934_416934;
   reg _416935_416935 ; 
   reg __416935_416935;
   reg _416936_416936 ; 
   reg __416936_416936;
   reg _416937_416937 ; 
   reg __416937_416937;
   reg _416938_416938 ; 
   reg __416938_416938;
   reg _416939_416939 ; 
   reg __416939_416939;
   reg _416940_416940 ; 
   reg __416940_416940;
   reg _416941_416941 ; 
   reg __416941_416941;
   reg _416942_416942 ; 
   reg __416942_416942;
   reg _416943_416943 ; 
   reg __416943_416943;
   reg _416944_416944 ; 
   reg __416944_416944;
   reg _416945_416945 ; 
   reg __416945_416945;
   reg _416946_416946 ; 
   reg __416946_416946;
   reg _416947_416947 ; 
   reg __416947_416947;
   reg _416948_416948 ; 
   reg __416948_416948;
   reg _416949_416949 ; 
   reg __416949_416949;
   reg _416950_416950 ; 
   reg __416950_416950;
   reg _416951_416951 ; 
   reg __416951_416951;
   reg _416952_416952 ; 
   reg __416952_416952;
   reg _416953_416953 ; 
   reg __416953_416953;
   reg _416954_416954 ; 
   reg __416954_416954;
   reg _416955_416955 ; 
   reg __416955_416955;
   reg _416956_416956 ; 
   reg __416956_416956;
   reg _416957_416957 ; 
   reg __416957_416957;
   reg _416958_416958 ; 
   reg __416958_416958;
   reg _416959_416959 ; 
   reg __416959_416959;
   reg _416960_416960 ; 
   reg __416960_416960;
   reg _416961_416961 ; 
   reg __416961_416961;
   reg _416962_416962 ; 
   reg __416962_416962;
   reg _416963_416963 ; 
   reg __416963_416963;
   reg _416964_416964 ; 
   reg __416964_416964;
   reg _416965_416965 ; 
   reg __416965_416965;
   reg _416966_416966 ; 
   reg __416966_416966;
   reg _416967_416967 ; 
   reg __416967_416967;
   reg _416968_416968 ; 
   reg __416968_416968;
   reg _416969_416969 ; 
   reg __416969_416969;
   reg _416970_416970 ; 
   reg __416970_416970;
   reg _416971_416971 ; 
   reg __416971_416971;
   reg _416972_416972 ; 
   reg __416972_416972;
   reg _416973_416973 ; 
   reg __416973_416973;
   reg _416974_416974 ; 
   reg __416974_416974;
   reg _416975_416975 ; 
   reg __416975_416975;
   reg _416976_416976 ; 
   reg __416976_416976;
   reg _416977_416977 ; 
   reg __416977_416977;
   reg _416978_416978 ; 
   reg __416978_416978;
   reg _416979_416979 ; 
   reg __416979_416979;
   reg _416980_416980 ; 
   reg __416980_416980;
   reg _416981_416981 ; 
   reg __416981_416981;
   reg _416982_416982 ; 
   reg __416982_416982;
   reg _416983_416983 ; 
   reg __416983_416983;
   reg _416984_416984 ; 
   reg __416984_416984;
   reg _416985_416985 ; 
   reg __416985_416985;
   reg _416986_416986 ; 
   reg __416986_416986;
   reg _416987_416987 ; 
   reg __416987_416987;
   reg _416988_416988 ; 
   reg __416988_416988;
   reg _416989_416989 ; 
   reg __416989_416989;
   reg _416990_416990 ; 
   reg __416990_416990;
   reg _416991_416991 ; 
   reg __416991_416991;
   reg _416992_416992 ; 
   reg __416992_416992;
   reg _416993_416993 ; 
   reg __416993_416993;
   reg _416994_416994 ; 
   reg __416994_416994;
   reg _416995_416995 ; 
   reg __416995_416995;
   reg _416996_416996 ; 
   reg __416996_416996;
   reg _416997_416997 ; 
   reg __416997_416997;
   reg _416998_416998 ; 
   reg __416998_416998;
   reg _416999_416999 ; 
   reg __416999_416999;
   reg _417000_417000 ; 
   reg __417000_417000;
   reg _417001_417001 ; 
   reg __417001_417001;
   reg _417002_417002 ; 
   reg __417002_417002;
   reg _417003_417003 ; 
   reg __417003_417003;
   reg _417004_417004 ; 
   reg __417004_417004;
   reg _417005_417005 ; 
   reg __417005_417005;
   reg _417006_417006 ; 
   reg __417006_417006;
   reg _417007_417007 ; 
   reg __417007_417007;
   reg _417008_417008 ; 
   reg __417008_417008;
   reg _417009_417009 ; 
   reg __417009_417009;
   reg _417010_417010 ; 
   reg __417010_417010;
   reg _417011_417011 ; 
   reg __417011_417011;
   reg _417012_417012 ; 
   reg __417012_417012;
   reg _417013_417013 ; 
   reg __417013_417013;
   reg _417014_417014 ; 
   reg __417014_417014;
   reg _417015_417015 ; 
   reg __417015_417015;
   reg _417016_417016 ; 
   reg __417016_417016;
   reg _417017_417017 ; 
   reg __417017_417017;
   reg _417018_417018 ; 
   reg __417018_417018;
   reg _417019_417019 ; 
   reg __417019_417019;
   reg _417020_417020 ; 
   reg __417020_417020;
   reg _417021_417021 ; 
   reg __417021_417021;
   reg _417022_417022 ; 
   reg __417022_417022;
   reg _417023_417023 ; 
   reg __417023_417023;
   reg _417024_417024 ; 
   reg __417024_417024;
   reg _417025_417025 ; 
   reg __417025_417025;
   reg _417026_417026 ; 
   reg __417026_417026;
   reg _417027_417027 ; 
   reg __417027_417027;
   reg _417028_417028 ; 
   reg __417028_417028;
   reg _417029_417029 ; 
   reg __417029_417029;
   reg _417030_417030 ; 
   reg __417030_417030;
   reg _417031_417031 ; 
   reg __417031_417031;
   reg _417032_417032 ; 
   reg __417032_417032;
   reg _417033_417033 ; 
   reg __417033_417033;
   reg _417034_417034 ; 
   reg __417034_417034;
   reg _417035_417035 ; 
   reg __417035_417035;
   reg _417036_417036 ; 
   reg __417036_417036;
   reg _417037_417037 ; 
   reg __417037_417037;
   reg _417038_417038 ; 
   reg __417038_417038;
   reg _417039_417039 ; 
   reg __417039_417039;
   reg _417040_417040 ; 
   reg __417040_417040;
   reg _417041_417041 ; 
   reg __417041_417041;
   reg _417042_417042 ; 
   reg __417042_417042;
   reg _417043_417043 ; 
   reg __417043_417043;
   reg _417044_417044 ; 
   reg __417044_417044;
   reg _417045_417045 ; 
   reg __417045_417045;
   reg _417046_417046 ; 
   reg __417046_417046;
   reg _417047_417047 ; 
   reg __417047_417047;
   reg _417048_417048 ; 
   reg __417048_417048;
   reg _417049_417049 ; 
   reg __417049_417049;
   reg _417050_417050 ; 
   reg __417050_417050;
   reg _417051_417051 ; 
   reg __417051_417051;
   reg _417052_417052 ; 
   reg __417052_417052;
   reg _417053_417053 ; 
   reg __417053_417053;
   reg _417054_417054 ; 
   reg __417054_417054;
   reg _417055_417055 ; 
   reg __417055_417055;
   reg _417056_417056 ; 
   reg __417056_417056;
   reg _417057_417057 ; 
   reg __417057_417057;
   reg _417058_417058 ; 
   reg __417058_417058;
   reg _417059_417059 ; 
   reg __417059_417059;
   reg _417060_417060 ; 
   reg __417060_417060;
   reg _417061_417061 ; 
   reg __417061_417061;
   reg _417062_417062 ; 
   reg __417062_417062;
   reg _417063_417063 ; 
   reg __417063_417063;
   reg _417064_417064 ; 
   reg __417064_417064;
   reg _417065_417065 ; 
   reg __417065_417065;
   reg _417066_417066 ; 
   reg __417066_417066;
   reg _417067_417067 ; 
   reg __417067_417067;
   reg _417068_417068 ; 
   reg __417068_417068;
   reg _417069_417069 ; 
   reg __417069_417069;
   reg _417070_417070 ; 
   reg __417070_417070;
   reg _417071_417071 ; 
   reg __417071_417071;
   reg _417072_417072 ; 
   reg __417072_417072;
   reg _417073_417073 ; 
   reg __417073_417073;
   reg _417074_417074 ; 
   reg __417074_417074;
   reg _417075_417075 ; 
   reg __417075_417075;
   reg _417076_417076 ; 
   reg __417076_417076;
   reg _417077_417077 ; 
   reg __417077_417077;
   reg _417078_417078 ; 
   reg __417078_417078;
   reg _417079_417079 ; 
   reg __417079_417079;
   reg _417080_417080 ; 
   reg __417080_417080;
   reg _417081_417081 ; 
   reg __417081_417081;
   reg _417082_417082 ; 
   reg __417082_417082;
   reg _417083_417083 ; 
   reg __417083_417083;
   reg _417084_417084 ; 
   reg __417084_417084;
   reg _417085_417085 ; 
   reg __417085_417085;
   reg _417086_417086 ; 
   reg __417086_417086;
   reg _417087_417087 ; 
   reg __417087_417087;
   reg _417088_417088 ; 
   reg __417088_417088;
   reg _417089_417089 ; 
   reg __417089_417089;
   reg _417090_417090 ; 
   reg __417090_417090;
   reg _417091_417091 ; 
   reg __417091_417091;
   reg _417092_417092 ; 
   reg __417092_417092;
   reg _417093_417093 ; 
   reg __417093_417093;
   reg _417094_417094 ; 
   reg __417094_417094;
   reg _417095_417095 ; 
   reg __417095_417095;
   reg _417096_417096 ; 
   reg __417096_417096;
   reg _417097_417097 ; 
   reg __417097_417097;
   reg _417098_417098 ; 
   reg __417098_417098;
   reg _417099_417099 ; 
   reg __417099_417099;
   reg _417100_417100 ; 
   reg __417100_417100;
   reg _417101_417101 ; 
   reg __417101_417101;
   reg _417102_417102 ; 
   reg __417102_417102;
   reg _417103_417103 ; 
   reg __417103_417103;
   reg _417104_417104 ; 
   reg __417104_417104;
   reg _417105_417105 ; 
   reg __417105_417105;
   reg _417106_417106 ; 
   reg __417106_417106;
   reg _417107_417107 ; 
   reg __417107_417107;
   reg _417108_417108 ; 
   reg __417108_417108;
   reg _417109_417109 ; 
   reg __417109_417109;
   reg _417110_417110 ; 
   reg __417110_417110;
   reg _417111_417111 ; 
   reg __417111_417111;
   reg _417112_417112 ; 
   reg __417112_417112;
   reg _417113_417113 ; 
   reg __417113_417113;
   reg _417114_417114 ; 
   reg __417114_417114;
   reg _417115_417115 ; 
   reg __417115_417115;
   reg _417116_417116 ; 
   reg __417116_417116;
   reg _417117_417117 ; 
   reg __417117_417117;
   reg _417118_417118 ; 
   reg __417118_417118;
   reg _417119_417119 ; 
   reg __417119_417119;
   reg _417120_417120 ; 
   reg __417120_417120;
   reg _417121_417121 ; 
   reg __417121_417121;
   reg _417122_417122 ; 
   reg __417122_417122;
   reg _417123_417123 ; 
   reg __417123_417123;
   reg _417124_417124 ; 
   reg __417124_417124;
   reg _417125_417125 ; 
   reg __417125_417125;
   reg _417126_417126 ; 
   reg __417126_417126;
   reg _417127_417127 ; 
   reg __417127_417127;
   reg _417128_417128 ; 
   reg __417128_417128;
   reg _417129_417129 ; 
   reg __417129_417129;
   reg _417130_417130 ; 
   reg __417130_417130;
   reg _417131_417131 ; 
   reg __417131_417131;
   reg _417132_417132 ; 
   reg __417132_417132;
   reg _417133_417133 ; 
   reg __417133_417133;
   reg _417134_417134 ; 
   reg __417134_417134;
   reg _417135_417135 ; 
   reg __417135_417135;
   reg _417136_417136 ; 
   reg __417136_417136;
   reg _417137_417137 ; 
   reg __417137_417137;
   reg _417138_417138 ; 
   reg __417138_417138;
   reg _417139_417139 ; 
   reg __417139_417139;
   reg _417140_417140 ; 
   reg __417140_417140;
   reg _417141_417141 ; 
   reg __417141_417141;
   reg _417142_417142 ; 
   reg __417142_417142;
   reg _417143_417143 ; 
   reg __417143_417143;
   reg _417144_417144 ; 
   reg __417144_417144;
   reg _417145_417145 ; 
   reg __417145_417145;
   reg _417146_417146 ; 
   reg __417146_417146;
   reg _417147_417147 ; 
   reg __417147_417147;
   reg _417148_417148 ; 
   reg __417148_417148;
   reg _417149_417149 ; 
   reg __417149_417149;
   reg _417150_417150 ; 
   reg __417150_417150;
   reg _417151_417151 ; 
   reg __417151_417151;
   reg _417152_417152 ; 
   reg __417152_417152;
   reg _417153_417153 ; 
   reg __417153_417153;
   reg _417154_417154 ; 
   reg __417154_417154;
   reg _417155_417155 ; 
   reg __417155_417155;
   reg _417156_417156 ; 
   reg __417156_417156;
   reg _417157_417157 ; 
   reg __417157_417157;
   reg _417158_417158 ; 
   reg __417158_417158;
   reg _417159_417159 ; 
   reg __417159_417159;
   reg _417160_417160 ; 
   reg __417160_417160;
   reg _417161_417161 ; 
   reg __417161_417161;
   reg _417162_417162 ; 
   reg __417162_417162;
   reg _417163_417163 ; 
   reg __417163_417163;
   reg _417164_417164 ; 
   reg __417164_417164;
   reg _417165_417165 ; 
   reg __417165_417165;
   reg _417166_417166 ; 
   reg __417166_417166;
   reg _417167_417167 ; 
   reg __417167_417167;
   reg _417168_417168 ; 
   reg __417168_417168;
   reg _417169_417169 ; 
   reg __417169_417169;
   reg _417170_417170 ; 
   reg __417170_417170;
   reg _417171_417171 ; 
   reg __417171_417171;
   reg _417172_417172 ; 
   reg __417172_417172;
   reg _417173_417173 ; 
   reg __417173_417173;
   reg _417174_417174 ; 
   reg __417174_417174;
   reg _417175_417175 ; 
   reg __417175_417175;
   reg _417176_417176 ; 
   reg __417176_417176;
   reg _417177_417177 ; 
   reg __417177_417177;
   reg _417178_417178 ; 
   reg __417178_417178;
   reg _417179_417179 ; 
   reg __417179_417179;
   reg _417180_417180 ; 
   reg __417180_417180;
   reg _417181_417181 ; 
   reg __417181_417181;
   reg _417182_417182 ; 
   reg __417182_417182;
   reg _417183_417183 ; 
   reg __417183_417183;
   reg _417184_417184 ; 
   reg __417184_417184;
   reg _417185_417185 ; 
   reg __417185_417185;
   reg _417186_417186 ; 
   reg __417186_417186;
   reg _417187_417187 ; 
   reg __417187_417187;
   reg _417188_417188 ; 
   reg __417188_417188;
   reg _417189_417189 ; 
   reg __417189_417189;
   reg _417190_417190 ; 
   reg __417190_417190;
   reg _417191_417191 ; 
   reg __417191_417191;
   reg _417192_417192 ; 
   reg __417192_417192;
   reg _417193_417193 ; 
   reg __417193_417193;
   reg _417194_417194 ; 
   reg __417194_417194;
   reg _417195_417195 ; 
   reg __417195_417195;
   reg _417196_417196 ; 
   reg __417196_417196;
   reg _417197_417197 ; 
   reg __417197_417197;
   reg _417198_417198 ; 
   reg __417198_417198;
   reg _417199_417199 ; 
   reg __417199_417199;
   reg _417200_417200 ; 
   reg __417200_417200;
   reg _417201_417201 ; 
   reg __417201_417201;
   reg _417202_417202 ; 
   reg __417202_417202;
   reg _417203_417203 ; 
   reg __417203_417203;
   reg _417204_417204 ; 
   reg __417204_417204;
   reg _417205_417205 ; 
   reg __417205_417205;
   reg _417206_417206 ; 
   reg __417206_417206;
   reg _417207_417207 ; 
   reg __417207_417207;
   reg _417208_417208 ; 
   reg __417208_417208;
   reg _417209_417209 ; 
   reg __417209_417209;
   reg _417210_417210 ; 
   reg __417210_417210;
   reg _417211_417211 ; 
   reg __417211_417211;
   reg _417212_417212 ; 
   reg __417212_417212;
   reg _417213_417213 ; 
   reg __417213_417213;
   reg _417214_417214 ; 
   reg __417214_417214;
   reg _417215_417215 ; 
   reg __417215_417215;
   reg _417216_417216 ; 
   reg __417216_417216;
   reg _417217_417217 ; 
   reg __417217_417217;
   reg _417218_417218 ; 
   reg __417218_417218;
   reg _417219_417219 ; 
   reg __417219_417219;
   reg _417220_417220 ; 
   reg __417220_417220;
   reg _417221_417221 ; 
   reg __417221_417221;
   reg _417222_417222 ; 
   reg __417222_417222;
   reg _417223_417223 ; 
   reg __417223_417223;
   reg _417224_417224 ; 
   reg __417224_417224;
   reg _417225_417225 ; 
   reg __417225_417225;
   reg _417226_417226 ; 
   reg __417226_417226;
   reg _417227_417227 ; 
   reg __417227_417227;
   reg _417228_417228 ; 
   reg __417228_417228;
   reg _417229_417229 ; 
   reg __417229_417229;
   reg _417230_417230 ; 
   reg __417230_417230;
   reg _417231_417231 ; 
   reg __417231_417231;
   reg _417232_417232 ; 
   reg __417232_417232;
   reg _417233_417233 ; 
   reg __417233_417233;
   reg _417234_417234 ; 
   reg __417234_417234;
   reg _417235_417235 ; 
   reg __417235_417235;
   reg _417236_417236 ; 
   reg __417236_417236;
   reg _417237_417237 ; 
   reg __417237_417237;
   reg _417238_417238 ; 
   reg __417238_417238;
   reg _417239_417239 ; 
   reg __417239_417239;
   reg _417240_417240 ; 
   reg __417240_417240;
   reg _417241_417241 ; 
   reg __417241_417241;
   reg _417242_417242 ; 
   reg __417242_417242;
   reg _417243_417243 ; 
   reg __417243_417243;
   reg _417244_417244 ; 
   reg __417244_417244;
   reg _417245_417245 ; 
   reg __417245_417245;
   reg _417246_417246 ; 
   reg __417246_417246;
   reg _417247_417247 ; 
   reg __417247_417247;
   reg _417248_417248 ; 
   reg __417248_417248;
   reg _417249_417249 ; 
   reg __417249_417249;
   reg _417250_417250 ; 
   reg __417250_417250;
   reg _417251_417251 ; 
   reg __417251_417251;
   reg _417252_417252 ; 
   reg __417252_417252;
   reg _417253_417253 ; 
   reg __417253_417253;
   reg _417254_417254 ; 
   reg __417254_417254;
   reg _417255_417255 ; 
   reg __417255_417255;
   reg _417256_417256 ; 
   reg __417256_417256;
   reg _417257_417257 ; 
   reg __417257_417257;
   reg _417258_417258 ; 
   reg __417258_417258;
   reg _417259_417259 ; 
   reg __417259_417259;
   reg _417260_417260 ; 
   reg __417260_417260;
   reg _417261_417261 ; 
   reg __417261_417261;
   reg _417262_417262 ; 
   reg __417262_417262;
   reg _417263_417263 ; 
   reg __417263_417263;
   reg _417264_417264 ; 
   reg __417264_417264;
   reg _417265_417265 ; 
   reg __417265_417265;
   reg _417266_417266 ; 
   reg __417266_417266;
   reg _417267_417267 ; 
   reg __417267_417267;
   reg _417268_417268 ; 
   reg __417268_417268;
   reg _417269_417269 ; 
   reg __417269_417269;
   reg _417270_417270 ; 
   reg __417270_417270;
   reg _417271_417271 ; 
   reg __417271_417271;
   reg _417272_417272 ; 
   reg __417272_417272;
   reg _417273_417273 ; 
   reg __417273_417273;
   reg _417274_417274 ; 
   reg __417274_417274;
   reg _417275_417275 ; 
   reg __417275_417275;
   reg _417276_417276 ; 
   reg __417276_417276;
   reg _417277_417277 ; 
   reg __417277_417277;
   reg _417278_417278 ; 
   reg __417278_417278;
   reg _417279_417279 ; 
   reg __417279_417279;
   reg _417280_417280 ; 
   reg __417280_417280;
   reg _417281_417281 ; 
   reg __417281_417281;
   reg _417282_417282 ; 
   reg __417282_417282;
   reg _417283_417283 ; 
   reg __417283_417283;
   reg _417284_417284 ; 
   reg __417284_417284;
   reg _417285_417285 ; 
   reg __417285_417285;
   reg _417286_417286 ; 
   reg __417286_417286;
   reg _417287_417287 ; 
   reg __417287_417287;
   reg _417288_417288 ; 
   reg __417288_417288;
   reg _417289_417289 ; 
   reg __417289_417289;
   reg _417290_417290 ; 
   reg __417290_417290;
   reg _417291_417291 ; 
   reg __417291_417291;
   reg _417292_417292 ; 
   reg __417292_417292;
   reg _417293_417293 ; 
   reg __417293_417293;
   reg _417294_417294 ; 
   reg __417294_417294;
   reg _417295_417295 ; 
   reg __417295_417295;
   reg _417296_417296 ; 
   reg __417296_417296;
   reg _417297_417297 ; 
   reg __417297_417297;
   reg _417298_417298 ; 
   reg __417298_417298;
   reg _417299_417299 ; 
   reg __417299_417299;
   reg _417300_417300 ; 
   reg __417300_417300;
   reg _417301_417301 ; 
   reg __417301_417301;
   reg _417302_417302 ; 
   reg __417302_417302;
   reg _417303_417303 ; 
   reg __417303_417303;
   reg _417304_417304 ; 
   reg __417304_417304;
   reg _417305_417305 ; 
   reg __417305_417305;
   reg _417306_417306 ; 
   reg __417306_417306;
   reg _417307_417307 ; 
   reg __417307_417307;
   reg _417308_417308 ; 
   reg __417308_417308;
   reg _417309_417309 ; 
   reg __417309_417309;
   reg _417310_417310 ; 
   reg __417310_417310;
   reg _417311_417311 ; 
   reg __417311_417311;
   reg _417312_417312 ; 
   reg __417312_417312;
   reg _417313_417313 ; 
   reg __417313_417313;
   reg _417314_417314 ; 
   reg __417314_417314;
   reg _417315_417315 ; 
   reg __417315_417315;
   reg _417316_417316 ; 
   reg __417316_417316;
   reg _417317_417317 ; 
   reg __417317_417317;
   reg _417318_417318 ; 
   reg __417318_417318;
   reg _417319_417319 ; 
   reg __417319_417319;
   reg _417320_417320 ; 
   reg __417320_417320;
   reg _417321_417321 ; 
   reg __417321_417321;
   reg _417322_417322 ; 
   reg __417322_417322;
   reg _417323_417323 ; 
   reg __417323_417323;
   reg _417324_417324 ; 
   reg __417324_417324;
   reg _417325_417325 ; 
   reg __417325_417325;
   reg _417326_417326 ; 
   reg __417326_417326;
   reg _417327_417327 ; 
   reg __417327_417327;
   reg _417328_417328 ; 
   reg __417328_417328;
   reg _417329_417329 ; 
   reg __417329_417329;
   reg _417330_417330 ; 
   reg __417330_417330;
   reg _417331_417331 ; 
   reg __417331_417331;
   reg _417332_417332 ; 
   reg __417332_417332;
   reg _417333_417333 ; 
   reg __417333_417333;
   reg _417334_417334 ; 
   reg __417334_417334;
   reg _417335_417335 ; 
   reg __417335_417335;
   reg _417336_417336 ; 
   reg __417336_417336;
   reg _417337_417337 ; 
   reg __417337_417337;
   reg _417338_417338 ; 
   reg __417338_417338;
   reg _417339_417339 ; 
   reg __417339_417339;
   reg _417340_417340 ; 
   reg __417340_417340;
   reg _417341_417341 ; 
   reg __417341_417341;
   reg _417342_417342 ; 
   reg __417342_417342;
   reg _417343_417343 ; 
   reg __417343_417343;
   reg _417344_417344 ; 
   reg __417344_417344;
   reg _417345_417345 ; 
   reg __417345_417345;
   reg _417346_417346 ; 
   reg __417346_417346;
   reg _417347_417347 ; 
   reg __417347_417347;
   reg _417348_417348 ; 
   reg __417348_417348;
   reg _417349_417349 ; 
   reg __417349_417349;
   reg _417350_417350 ; 
   reg __417350_417350;
   reg _417351_417351 ; 
   reg __417351_417351;
   reg _417352_417352 ; 
   reg __417352_417352;
   reg _417353_417353 ; 
   reg __417353_417353;
   reg _417354_417354 ; 
   reg __417354_417354;
   reg _417355_417355 ; 
   reg __417355_417355;
   reg _417356_417356 ; 
   reg __417356_417356;
   reg _417357_417357 ; 
   reg __417357_417357;
   reg _417358_417358 ; 
   reg __417358_417358;
   reg _417359_417359 ; 
   reg __417359_417359;
   reg _417360_417360 ; 
   reg __417360_417360;
   reg _417361_417361 ; 
   reg __417361_417361;
   reg _417362_417362 ; 
   reg __417362_417362;
   reg _417363_417363 ; 
   reg __417363_417363;
   reg _417364_417364 ; 
   reg __417364_417364;
   reg _417365_417365 ; 
   reg __417365_417365;
   reg _417366_417366 ; 
   reg __417366_417366;
   reg _417367_417367 ; 
   reg __417367_417367;
   reg _417368_417368 ; 
   reg __417368_417368;
   reg _417369_417369 ; 
   reg __417369_417369;
   reg _417370_417370 ; 
   reg __417370_417370;
   reg _417371_417371 ; 
   reg __417371_417371;
   reg _417372_417372 ; 
   reg __417372_417372;
   reg _417373_417373 ; 
   reg __417373_417373;
   reg _417374_417374 ; 
   reg __417374_417374;
   reg _417375_417375 ; 
   reg __417375_417375;
   reg _417376_417376 ; 
   reg __417376_417376;
   reg _417377_417377 ; 
   reg __417377_417377;
   reg _417378_417378 ; 
   reg __417378_417378;
   reg _417379_417379 ; 
   reg __417379_417379;
   reg _417380_417380 ; 
   reg __417380_417380;
   reg _417381_417381 ; 
   reg __417381_417381;
   reg _417382_417382 ; 
   reg __417382_417382;
   reg _417383_417383 ; 
   reg __417383_417383;
   reg _417384_417384 ; 
   reg __417384_417384;
   reg _417385_417385 ; 
   reg __417385_417385;
   reg _417386_417386 ; 
   reg __417386_417386;
   reg _417387_417387 ; 
   reg __417387_417387;
   reg _417388_417388 ; 
   reg __417388_417388;
   reg _417389_417389 ; 
   reg __417389_417389;
   reg _417390_417390 ; 
   reg __417390_417390;
   reg _417391_417391 ; 
   reg __417391_417391;
   reg _417392_417392 ; 
   reg __417392_417392;
   reg _417393_417393 ; 
   reg __417393_417393;
   reg _417394_417394 ; 
   reg __417394_417394;
   reg _417395_417395 ; 
   reg __417395_417395;
   reg _417396_417396 ; 
   reg __417396_417396;
   reg _417397_417397 ; 
   reg __417397_417397;
   reg _417398_417398 ; 
   reg __417398_417398;
   reg _417399_417399 ; 
   reg __417399_417399;
   reg _417400_417400 ; 
   reg __417400_417400;
   reg _417401_417401 ; 
   reg __417401_417401;
   reg _417402_417402 ; 
   reg __417402_417402;
   reg _417403_417403 ; 
   reg __417403_417403;
   reg _417404_417404 ; 
   reg __417404_417404;
   reg _417405_417405 ; 
   reg __417405_417405;
   reg _417406_417406 ; 
   reg __417406_417406;
   reg _417407_417407 ; 
   reg __417407_417407;
   reg _417408_417408 ; 
   reg __417408_417408;
   reg _417409_417409 ; 
   reg __417409_417409;
   reg _417410_417410 ; 
   reg __417410_417410;
   reg _417411_417411 ; 
   reg __417411_417411;
   reg _417412_417412 ; 
   reg __417412_417412;
   reg _417413_417413 ; 
   reg __417413_417413;
   reg _417414_417414 ; 
   reg __417414_417414;
   reg _417415_417415 ; 
   reg __417415_417415;
   reg _417416_417416 ; 
   reg __417416_417416;
   reg _417417_417417 ; 
   reg __417417_417417;
   reg _417418_417418 ; 
   reg __417418_417418;
   reg _417419_417419 ; 
   reg __417419_417419;
   reg _417420_417420 ; 
   reg __417420_417420;
   reg _417421_417421 ; 
   reg __417421_417421;
   reg _417422_417422 ; 
   reg __417422_417422;
   reg _417423_417423 ; 
   reg __417423_417423;
   reg _417424_417424 ; 
   reg __417424_417424;
   reg _417425_417425 ; 
   reg __417425_417425;
   reg _417426_417426 ; 
   reg __417426_417426;
   reg _417427_417427 ; 
   reg __417427_417427;
   reg _417428_417428 ; 
   reg __417428_417428;
   reg _417429_417429 ; 
   reg __417429_417429;
   reg _417430_417430 ; 
   reg __417430_417430;
   reg _417431_417431 ; 
   reg __417431_417431;
   reg _417432_417432 ; 
   reg __417432_417432;
   reg _417433_417433 ; 
   reg __417433_417433;
   reg _417434_417434 ; 
   reg __417434_417434;
   reg _417435_417435 ; 
   reg __417435_417435;
   reg _417436_417436 ; 
   reg __417436_417436;
   reg _417437_417437 ; 
   reg __417437_417437;
   reg _417438_417438 ; 
   reg __417438_417438;
   reg _417439_417439 ; 
   reg __417439_417439;
   reg _417440_417440 ; 
   reg __417440_417440;
   reg _417441_417441 ; 
   reg __417441_417441;
   reg _417442_417442 ; 
   reg __417442_417442;
   reg _417443_417443 ; 
   reg __417443_417443;
   reg _417444_417444 ; 
   reg __417444_417444;
   reg _417445_417445 ; 
   reg __417445_417445;
   reg _417446_417446 ; 
   reg __417446_417446;
   reg _417447_417447 ; 
   reg __417447_417447;
   reg _417448_417448 ; 
   reg __417448_417448;
   reg _417449_417449 ; 
   reg __417449_417449;
   reg _417450_417450 ; 
   reg __417450_417450;
   reg _417451_417451 ; 
   reg __417451_417451;
   reg _417452_417452 ; 
   reg __417452_417452;
   reg _417453_417453 ; 
   reg __417453_417453;
   reg _417454_417454 ; 
   reg __417454_417454;
   reg _417455_417455 ; 
   reg __417455_417455;
   reg _417456_417456 ; 
   reg __417456_417456;
   reg _417457_417457 ; 
   reg __417457_417457;
   reg _417458_417458 ; 
   reg __417458_417458;
   reg _417459_417459 ; 
   reg __417459_417459;
   reg _417460_417460 ; 
   reg __417460_417460;
   reg _417461_417461 ; 
   reg __417461_417461;
   reg _417462_417462 ; 
   reg __417462_417462;
   reg _417463_417463 ; 
   reg __417463_417463;
   reg _417464_417464 ; 
   reg __417464_417464;
   reg _417465_417465 ; 
   reg __417465_417465;
   reg _417466_417466 ; 
   reg __417466_417466;
   reg _417467_417467 ; 
   reg __417467_417467;
   reg _417468_417468 ; 
   reg __417468_417468;
   reg _417469_417469 ; 
   reg __417469_417469;
   reg _417470_417470 ; 
   reg __417470_417470;
   reg _417471_417471 ; 
   reg __417471_417471;
   reg _417472_417472 ; 
   reg __417472_417472;
   reg _417473_417473 ; 
   reg __417473_417473;
   reg _417474_417474 ; 
   reg __417474_417474;
   reg _417475_417475 ; 
   reg __417475_417475;
   reg _417476_417476 ; 
   reg __417476_417476;
   reg _417477_417477 ; 
   reg __417477_417477;
   reg _417478_417478 ; 
   reg __417478_417478;
   reg _417479_417479 ; 
   reg __417479_417479;
   reg _417480_417480 ; 
   reg __417480_417480;
   reg _417481_417481 ; 
   reg __417481_417481;
   reg _417482_417482 ; 
   reg __417482_417482;
   reg _417483_417483 ; 
   reg __417483_417483;
   reg _417484_417484 ; 
   reg __417484_417484;
   reg _417485_417485 ; 
   reg __417485_417485;
   reg _417486_417486 ; 
   reg __417486_417486;
   reg _417487_417487 ; 
   reg __417487_417487;
   reg _417488_417488 ; 
   reg __417488_417488;
   reg _417489_417489 ; 
   reg __417489_417489;
   reg _417490_417490 ; 
   reg __417490_417490;
   reg _417491_417491 ; 
   reg __417491_417491;
   reg _417492_417492 ; 
   reg __417492_417492;
   reg _417493_417493 ; 
   reg __417493_417493;
   reg _417494_417494 ; 
   reg __417494_417494;
   reg _417495_417495 ; 
   reg __417495_417495;
   reg _417496_417496 ; 
   reg __417496_417496;
   reg _417497_417497 ; 
   reg __417497_417497;
   reg _417498_417498 ; 
   reg __417498_417498;
   reg _417499_417499 ; 
   reg __417499_417499;
   reg _417500_417500 ; 
   reg __417500_417500;
   reg _417501_417501 ; 
   reg __417501_417501;
   reg _417502_417502 ; 
   reg __417502_417502;
   reg _417503_417503 ; 
   reg __417503_417503;
   reg _417504_417504 ; 
   reg __417504_417504;
   reg _417505_417505 ; 
   reg __417505_417505;
   reg _417506_417506 ; 
   reg __417506_417506;
   reg _417507_417507 ; 
   reg __417507_417507;
   reg _417508_417508 ; 
   reg __417508_417508;
   reg _417509_417509 ; 
   reg __417509_417509;
   reg _417510_417510 ; 
   reg __417510_417510;
   reg _417511_417511 ; 
   reg __417511_417511;
   reg _417512_417512 ; 
   reg __417512_417512;
   reg _417513_417513 ; 
   reg __417513_417513;
   reg _417514_417514 ; 
   reg __417514_417514;
   reg _417515_417515 ; 
   reg __417515_417515;
   reg _417516_417516 ; 
   reg __417516_417516;
   reg _417517_417517 ; 
   reg __417517_417517;
   reg _417518_417518 ; 
   reg __417518_417518;
   reg _417519_417519 ; 
   reg __417519_417519;
   reg _417520_417520 ; 
   reg __417520_417520;
   reg _417521_417521 ; 
   reg __417521_417521;
   reg _417522_417522 ; 
   reg __417522_417522;
   reg _417523_417523 ; 
   reg __417523_417523;
   reg _417524_417524 ; 
   reg __417524_417524;
   reg _417525_417525 ; 
   reg __417525_417525;
   reg _417526_417526 ; 
   reg __417526_417526;
   reg _417527_417527 ; 
   reg __417527_417527;
   reg _417528_417528 ; 
   reg __417528_417528;
   reg _417529_417529 ; 
   reg __417529_417529;
   reg _417530_417530 ; 
   reg __417530_417530;
   reg _417531_417531 ; 
   reg __417531_417531;
   reg _417532_417532 ; 
   reg __417532_417532;
   reg _417533_417533 ; 
   reg __417533_417533;
   reg _417534_417534 ; 
   reg __417534_417534;
   reg _417535_417535 ; 
   reg __417535_417535;
   reg _417536_417536 ; 
   reg __417536_417536;
   reg _417537_417537 ; 
   reg __417537_417537;
   reg _417538_417538 ; 
   reg __417538_417538;
   reg _417539_417539 ; 
   reg __417539_417539;
   reg _417540_417540 ; 
   reg __417540_417540;
   reg _417541_417541 ; 
   reg __417541_417541;
   reg _417542_417542 ; 
   reg __417542_417542;
   reg _417543_417543 ; 
   reg __417543_417543;
   reg _417544_417544 ; 
   reg __417544_417544;
   reg _417545_417545 ; 
   reg __417545_417545;
   reg _417546_417546 ; 
   reg __417546_417546;
   reg _417547_417547 ; 
   reg __417547_417547;
   reg _417548_417548 ; 
   reg __417548_417548;
   reg _417549_417549 ; 
   reg __417549_417549;
   reg _417550_417550 ; 
   reg __417550_417550;
   reg _417551_417551 ; 
   reg __417551_417551;
   reg _417552_417552 ; 
   reg __417552_417552;
   reg _417553_417553 ; 
   reg __417553_417553;
   reg _417554_417554 ; 
   reg __417554_417554;
   reg _417555_417555 ; 
   reg __417555_417555;
   reg _417556_417556 ; 
   reg __417556_417556;
   reg _417557_417557 ; 
   reg __417557_417557;
   reg _417558_417558 ; 
   reg __417558_417558;
   reg _417559_417559 ; 
   reg __417559_417559;
   reg _417560_417560 ; 
   reg __417560_417560;
   reg _417561_417561 ; 
   reg __417561_417561;
   reg _417562_417562 ; 
   reg __417562_417562;
   reg _417563_417563 ; 
   reg __417563_417563;
   reg _417564_417564 ; 
   reg __417564_417564;
   reg _417565_417565 ; 
   reg __417565_417565;
   reg _417566_417566 ; 
   reg __417566_417566;
   reg _417567_417567 ; 
   reg __417567_417567;
   reg _417568_417568 ; 
   reg __417568_417568;
   reg _417569_417569 ; 
   reg __417569_417569;
   reg _417570_417570 ; 
   reg __417570_417570;
   reg _417571_417571 ; 
   reg __417571_417571;
   reg _417572_417572 ; 
   reg __417572_417572;
   reg _417573_417573 ; 
   reg __417573_417573;
   reg _417574_417574 ; 
   reg __417574_417574;
   reg _417575_417575 ; 
   reg __417575_417575;
   reg _417576_417576 ; 
   reg __417576_417576;
   reg _417577_417577 ; 
   reg __417577_417577;
   reg _417578_417578 ; 
   reg __417578_417578;
   reg _417579_417579 ; 
   reg __417579_417579;
   reg _417580_417580 ; 
   reg __417580_417580;
   reg _417581_417581 ; 
   reg __417581_417581;
   reg _417582_417582 ; 
   reg __417582_417582;
   reg _417583_417583 ; 
   reg __417583_417583;
   reg _417584_417584 ; 
   reg __417584_417584;
   reg _417585_417585 ; 
   reg __417585_417585;
   reg _417586_417586 ; 
   reg __417586_417586;
   reg _417587_417587 ; 
   reg __417587_417587;
   reg _417588_417588 ; 
   reg __417588_417588;
   reg _417589_417589 ; 
   reg __417589_417589;
   reg _417590_417590 ; 
   reg __417590_417590;
   reg _417591_417591 ; 
   reg __417591_417591;
   reg _417592_417592 ; 
   reg __417592_417592;
   reg _417593_417593 ; 
   reg __417593_417593;
   reg _417594_417594 ; 
   reg __417594_417594;
   reg _417595_417595 ; 
   reg __417595_417595;
   reg _417596_417596 ; 
   reg __417596_417596;
   reg _417597_417597 ; 
   reg __417597_417597;
   reg _417598_417598 ; 
   reg __417598_417598;
   reg _417599_417599 ; 
   reg __417599_417599;
   reg _417600_417600 ; 
   reg __417600_417600;
   reg _417601_417601 ; 
   reg __417601_417601;
   reg _417602_417602 ; 
   reg __417602_417602;
   reg _417603_417603 ; 
   reg __417603_417603;
   reg _417604_417604 ; 
   reg __417604_417604;
   reg _417605_417605 ; 
   reg __417605_417605;
   reg _417606_417606 ; 
   reg __417606_417606;
   reg _417607_417607 ; 
   reg __417607_417607;
   reg _417608_417608 ; 
   reg __417608_417608;
   reg _417609_417609 ; 
   reg __417609_417609;
   reg _417610_417610 ; 
   reg __417610_417610;
   reg _417611_417611 ; 
   reg __417611_417611;
   reg _417612_417612 ; 
   reg __417612_417612;
   reg _417613_417613 ; 
   reg __417613_417613;
   reg _417614_417614 ; 
   reg __417614_417614;
   reg _417615_417615 ; 
   reg __417615_417615;
   reg _417616_417616 ; 
   reg __417616_417616;
   reg _417617_417617 ; 
   reg __417617_417617;
   reg _417618_417618 ; 
   reg __417618_417618;
   reg _417619_417619 ; 
   reg __417619_417619;
   reg _417620_417620 ; 
   reg __417620_417620;
   reg _417621_417621 ; 
   reg __417621_417621;
   reg _417622_417622 ; 
   reg __417622_417622;
   reg _417623_417623 ; 
   reg __417623_417623;
   reg _417624_417624 ; 
   reg __417624_417624;
   reg _417625_417625 ; 
   reg __417625_417625;
   reg _417626_417626 ; 
   reg __417626_417626;
   reg _417627_417627 ; 
   reg __417627_417627;
   reg _417628_417628 ; 
   reg __417628_417628;
   reg _417629_417629 ; 
   reg __417629_417629;
   reg _417630_417630 ; 
   reg __417630_417630;
   reg _417631_417631 ; 
   reg __417631_417631;
   reg _417632_417632 ; 
   reg __417632_417632;
   reg _417633_417633 ; 
   reg __417633_417633;
   reg _417634_417634 ; 
   reg __417634_417634;
   reg _417635_417635 ; 
   reg __417635_417635;
   reg _417636_417636 ; 
   reg __417636_417636;
   reg _417637_417637 ; 
   reg __417637_417637;
   reg _417638_417638 ; 
   reg __417638_417638;
   reg _417639_417639 ; 
   reg __417639_417639;
   reg _417640_417640 ; 
   reg __417640_417640;
   reg _417641_417641 ; 
   reg __417641_417641;
   reg _417642_417642 ; 
   reg __417642_417642;
   reg _417643_417643 ; 
   reg __417643_417643;
   reg _417644_417644 ; 
   reg __417644_417644;
   reg _417645_417645 ; 
   reg __417645_417645;
   reg _417646_417646 ; 
   reg __417646_417646;
   reg _417647_417647 ; 
   reg __417647_417647;
   reg _417648_417648 ; 
   reg __417648_417648;
   reg _417649_417649 ; 
   reg __417649_417649;
   reg _417650_417650 ; 
   reg __417650_417650;
   reg _417651_417651 ; 
   reg __417651_417651;
   reg _417652_417652 ; 
   reg __417652_417652;
   reg _417653_417653 ; 
   reg __417653_417653;
   reg _417654_417654 ; 
   reg __417654_417654;
   reg _417655_417655 ; 
   reg __417655_417655;
   reg _417656_417656 ; 
   reg __417656_417656;
   reg _417657_417657 ; 
   reg __417657_417657;
   reg _417658_417658 ; 
   reg __417658_417658;
   reg _417659_417659 ; 
   reg __417659_417659;
   reg _417660_417660 ; 
   reg __417660_417660;
   reg _417661_417661 ; 
   reg __417661_417661;
   reg _417662_417662 ; 
   reg __417662_417662;
   reg _417663_417663 ; 
   reg __417663_417663;
   reg _417664_417664 ; 
   reg __417664_417664;
   reg _417665_417665 ; 
   reg __417665_417665;
   reg _417666_417666 ; 
   reg __417666_417666;
   reg _417667_417667 ; 
   reg __417667_417667;
   reg _417668_417668 ; 
   reg __417668_417668;
   reg _417669_417669 ; 
   reg __417669_417669;
   reg _417670_417670 ; 
   reg __417670_417670;
   reg _417671_417671 ; 
   reg __417671_417671;
   reg _417672_417672 ; 
   reg __417672_417672;
   reg _417673_417673 ; 
   reg __417673_417673;
   reg _417674_417674 ; 
   reg __417674_417674;
   reg _417675_417675 ; 
   reg __417675_417675;
   reg _417676_417676 ; 
   reg __417676_417676;
   reg _417677_417677 ; 
   reg __417677_417677;
   reg _417678_417678 ; 
   reg __417678_417678;
   reg _417679_417679 ; 
   reg __417679_417679;
   reg _417680_417680 ; 
   reg __417680_417680;
   reg _417681_417681 ; 
   reg __417681_417681;
   reg _417682_417682 ; 
   reg __417682_417682;
   reg _417683_417683 ; 
   reg __417683_417683;
   reg _417684_417684 ; 
   reg __417684_417684;
   reg _417685_417685 ; 
   reg __417685_417685;
   reg _417686_417686 ; 
   reg __417686_417686;
   reg _417687_417687 ; 
   reg __417687_417687;
   reg _417688_417688 ; 
   reg __417688_417688;
   reg _417689_417689 ; 
   reg __417689_417689;
   reg _417690_417690 ; 
   reg __417690_417690;
   reg _417691_417691 ; 
   reg __417691_417691;
   reg _417692_417692 ; 
   reg __417692_417692;
   reg _417693_417693 ; 
   reg __417693_417693;
   reg _417694_417694 ; 
   reg __417694_417694;
   reg _417695_417695 ; 
   reg __417695_417695;
   reg _417696_417696 ; 
   reg __417696_417696;
   reg _417697_417697 ; 
   reg __417697_417697;
   reg _417698_417698 ; 
   reg __417698_417698;
   reg _417699_417699 ; 
   reg __417699_417699;
   reg _417700_417700 ; 
   reg __417700_417700;
   reg _417701_417701 ; 
   reg __417701_417701;
   reg _417702_417702 ; 
   reg __417702_417702;
   reg _417703_417703 ; 
   reg __417703_417703;
   reg _417704_417704 ; 
   reg __417704_417704;
   reg _417705_417705 ; 
   reg __417705_417705;
   reg _417706_417706 ; 
   reg __417706_417706;
   reg _417707_417707 ; 
   reg __417707_417707;
   reg _417708_417708 ; 
   reg __417708_417708;
   reg _417709_417709 ; 
   reg __417709_417709;
   reg _417710_417710 ; 
   reg __417710_417710;
   reg _417711_417711 ; 
   reg __417711_417711;
   reg _417712_417712 ; 
   reg __417712_417712;
   reg _417713_417713 ; 
   reg __417713_417713;
   reg _417714_417714 ; 
   reg __417714_417714;
   reg _417715_417715 ; 
   reg __417715_417715;
   reg _417716_417716 ; 
   reg __417716_417716;
   reg _417717_417717 ; 
   reg __417717_417717;
   reg _417718_417718 ; 
   reg __417718_417718;
   reg _417719_417719 ; 
   reg __417719_417719;
   reg _417720_417720 ; 
   reg __417720_417720;
   reg _417721_417721 ; 
   reg __417721_417721;
   reg _417722_417722 ; 
   reg __417722_417722;
   reg _417723_417723 ; 
   reg __417723_417723;
   reg _417724_417724 ; 
   reg __417724_417724;
   reg _417725_417725 ; 
   reg __417725_417725;
   reg _417726_417726 ; 
   reg __417726_417726;
   reg _417727_417727 ; 
   reg __417727_417727;
   reg _417728_417728 ; 
   reg __417728_417728;
   reg _417729_417729 ; 
   reg __417729_417729;
   reg _417730_417730 ; 
   reg __417730_417730;
   reg _417731_417731 ; 
   reg __417731_417731;
   reg _417732_417732 ; 
   reg __417732_417732;
   reg _417733_417733 ; 
   reg __417733_417733;
   reg _417734_417734 ; 
   reg __417734_417734;
   reg _417735_417735 ; 
   reg __417735_417735;
   reg _417736_417736 ; 
   reg __417736_417736;
   reg _417737_417737 ; 
   reg __417737_417737;
   reg _417738_417738 ; 
   reg __417738_417738;
   reg _417739_417739 ; 
   reg __417739_417739;
   reg _417740_417740 ; 
   reg __417740_417740;
   reg _417741_417741 ; 
   reg __417741_417741;
   reg _417742_417742 ; 
   reg __417742_417742;
   reg _417743_417743 ; 
   reg __417743_417743;
   reg _417744_417744 ; 
   reg __417744_417744;
   reg _417745_417745 ; 
   reg __417745_417745;
   reg _417746_417746 ; 
   reg __417746_417746;
   reg _417747_417747 ; 
   reg __417747_417747;
   reg _417748_417748 ; 
   reg __417748_417748;
   reg _417749_417749 ; 
   reg __417749_417749;
   reg _417750_417750 ; 
   reg __417750_417750;
   reg _417751_417751 ; 
   reg __417751_417751;
   reg _417752_417752 ; 
   reg __417752_417752;
   reg _417753_417753 ; 
   reg __417753_417753;
   reg _417754_417754 ; 
   reg __417754_417754;
   reg _417755_417755 ; 
   reg __417755_417755;
   reg _417756_417756 ; 
   reg __417756_417756;
   reg _417757_417757 ; 
   reg __417757_417757;
   reg _417758_417758 ; 
   reg __417758_417758;
   reg _417759_417759 ; 
   reg __417759_417759;
   reg _417760_417760 ; 
   reg __417760_417760;
   reg _417761_417761 ; 
   reg __417761_417761;
   reg _417762_417762 ; 
   reg __417762_417762;
   reg _417763_417763 ; 
   reg __417763_417763;
   reg _417764_417764 ; 
   reg __417764_417764;
   reg _417765_417765 ; 
   reg __417765_417765;
   reg _417766_417766 ; 
   reg __417766_417766;
   reg _417767_417767 ; 
   reg __417767_417767;
   reg _417768_417768 ; 
   reg __417768_417768;
   reg _417769_417769 ; 
   reg __417769_417769;
   reg _417770_417770 ; 
   reg __417770_417770;
   reg _417771_417771 ; 
   reg __417771_417771;
   reg _417772_417772 ; 
   reg __417772_417772;
   reg _417773_417773 ; 
   reg __417773_417773;
   reg _417774_417774 ; 
   reg __417774_417774;
   reg _417775_417775 ; 
   reg __417775_417775;
   reg _417776_417776 ; 
   reg __417776_417776;
   reg _417777_417777 ; 
   reg __417777_417777;
   reg _417778_417778 ; 
   reg __417778_417778;
   reg _417779_417779 ; 
   reg __417779_417779;
   reg _417780_417780 ; 
   reg __417780_417780;
   reg _417781_417781 ; 
   reg __417781_417781;
   reg _417782_417782 ; 
   reg __417782_417782;
   reg _417783_417783 ; 
   reg __417783_417783;
   reg _417784_417784 ; 
   reg __417784_417784;
   reg _417785_417785 ; 
   reg __417785_417785;
   reg _417786_417786 ; 
   reg __417786_417786;
   reg _417787_417787 ; 
   reg __417787_417787;
   reg _417788_417788 ; 
   reg __417788_417788;
   reg _417789_417789 ; 
   reg __417789_417789;
   reg _417790_417790 ; 
   reg __417790_417790;
   reg _417791_417791 ; 
   reg __417791_417791;
   reg _417792_417792 ; 
   reg __417792_417792;
   reg _417793_417793 ; 
   reg __417793_417793;
   reg _417794_417794 ; 
   reg __417794_417794;
   reg _417795_417795 ; 
   reg __417795_417795;
   reg _417796_417796 ; 
   reg __417796_417796;
   reg _417797_417797 ; 
   reg __417797_417797;
   reg _417798_417798 ; 
   reg __417798_417798;
   reg _417799_417799 ; 
   reg __417799_417799;
   reg _417800_417800 ; 
   reg __417800_417800;
   reg _417801_417801 ; 
   reg __417801_417801;
   reg _417802_417802 ; 
   reg __417802_417802;
   reg _417803_417803 ; 
   reg __417803_417803;
   reg _417804_417804 ; 
   reg __417804_417804;
   reg _417805_417805 ; 
   reg __417805_417805;
   reg _417806_417806 ; 
   reg __417806_417806;
   reg _417807_417807 ; 
   reg __417807_417807;
   reg _417808_417808 ; 
   reg __417808_417808;
   reg _417809_417809 ; 
   reg __417809_417809;
   reg _417810_417810 ; 
   reg __417810_417810;
   reg _417811_417811 ; 
   reg __417811_417811;
   reg _417812_417812 ; 
   reg __417812_417812;
   reg _417813_417813 ; 
   reg __417813_417813;
   reg _417814_417814 ; 
   reg __417814_417814;
   reg _417815_417815 ; 
   reg __417815_417815;
   reg _417816_417816 ; 
   reg __417816_417816;
   reg _417817_417817 ; 
   reg __417817_417817;
   reg _417818_417818 ; 
   reg __417818_417818;
   reg _417819_417819 ; 
   reg __417819_417819;
   reg _417820_417820 ; 
   reg __417820_417820;
   reg _417821_417821 ; 
   reg __417821_417821;
   reg _417822_417822 ; 
   reg __417822_417822;
   reg _417823_417823 ; 
   reg __417823_417823;
   reg _417824_417824 ; 
   reg __417824_417824;
   reg _417825_417825 ; 
   reg __417825_417825;
   reg _417826_417826 ; 
   reg __417826_417826;
   reg _417827_417827 ; 
   reg __417827_417827;
   reg _417828_417828 ; 
   reg __417828_417828;
   reg _417829_417829 ; 
   reg __417829_417829;
   reg _417830_417830 ; 
   reg __417830_417830;
   reg _417831_417831 ; 
   reg __417831_417831;
   reg _417832_417832 ; 
   reg __417832_417832;
   reg _417833_417833 ; 
   reg __417833_417833;
   reg _417834_417834 ; 
   reg __417834_417834;
   reg _417835_417835 ; 
   reg __417835_417835;
   reg _417836_417836 ; 
   reg __417836_417836;
   reg _417837_417837 ; 
   reg __417837_417837;
   reg _417838_417838 ; 
   reg __417838_417838;
   reg _417839_417839 ; 
   reg __417839_417839;
   reg _417840_417840 ; 
   reg __417840_417840;
   reg _417841_417841 ; 
   reg __417841_417841;
   reg _417842_417842 ; 
   reg __417842_417842;
   reg _417843_417843 ; 
   reg __417843_417843;
   reg _417844_417844 ; 
   reg __417844_417844;
   reg _417845_417845 ; 
   reg __417845_417845;
   reg _417846_417846 ; 
   reg __417846_417846;
   reg _417847_417847 ; 
   reg __417847_417847;
   reg _417848_417848 ; 
   reg __417848_417848;
   reg _417849_417849 ; 
   reg __417849_417849;
   reg _417850_417850 ; 
   reg __417850_417850;
   reg _417851_417851 ; 
   reg __417851_417851;
   reg _417852_417852 ; 
   reg __417852_417852;
   reg _417853_417853 ; 
   reg __417853_417853;
   reg _417854_417854 ; 
   reg __417854_417854;
   reg _417855_417855 ; 
   reg __417855_417855;
   reg _417856_417856 ; 
   reg __417856_417856;
   reg _417857_417857 ; 
   reg __417857_417857;
   reg _417858_417858 ; 
   reg __417858_417858;
   reg _417859_417859 ; 
   reg __417859_417859;
   reg _417860_417860 ; 
   reg __417860_417860;
   reg _417861_417861 ; 
   reg __417861_417861;
   reg _417862_417862 ; 
   reg __417862_417862;
   reg _417863_417863 ; 
   reg __417863_417863;
   reg _417864_417864 ; 
   reg __417864_417864;
   reg _417865_417865 ; 
   reg __417865_417865;
   reg _417866_417866 ; 
   reg __417866_417866;
   reg _417867_417867 ; 
   reg __417867_417867;
   reg _417868_417868 ; 
   reg __417868_417868;
   reg _417869_417869 ; 
   reg __417869_417869;
   reg _417870_417870 ; 
   reg __417870_417870;
   reg _417871_417871 ; 
   reg __417871_417871;
   reg _417872_417872 ; 
   reg __417872_417872;
   reg _417873_417873 ; 
   reg __417873_417873;
   reg _417874_417874 ; 
   reg __417874_417874;
   reg _417875_417875 ; 
   reg __417875_417875;
   reg _417876_417876 ; 
   reg __417876_417876;
   reg _417877_417877 ; 
   reg __417877_417877;
   reg _417878_417878 ; 
   reg __417878_417878;
   reg _417879_417879 ; 
   reg __417879_417879;
   reg _417880_417880 ; 
   reg __417880_417880;
   reg _417881_417881 ; 
   reg __417881_417881;
   reg _417882_417882 ; 
   reg __417882_417882;
   reg _417883_417883 ; 
   reg __417883_417883;
   reg _417884_417884 ; 
   reg __417884_417884;
   reg _417885_417885 ; 
   reg __417885_417885;
   reg _417886_417886 ; 
   reg __417886_417886;
   reg _417887_417887 ; 
   reg __417887_417887;
   reg _417888_417888 ; 
   reg __417888_417888;
   reg _417889_417889 ; 
   reg __417889_417889;
   reg _417890_417890 ; 
   reg __417890_417890;
   reg _417891_417891 ; 
   reg __417891_417891;
   reg _417892_417892 ; 
   reg __417892_417892;
   reg _417893_417893 ; 
   reg __417893_417893;
   reg _417894_417894 ; 
   reg __417894_417894;
   reg _417895_417895 ; 
   reg __417895_417895;
   reg _417896_417896 ; 
   reg __417896_417896;
   reg _417897_417897 ; 
   reg __417897_417897;
   reg _417898_417898 ; 
   reg __417898_417898;
   reg _417899_417899 ; 
   reg __417899_417899;
   reg _417900_417900 ; 
   reg __417900_417900;
   reg _417901_417901 ; 
   reg __417901_417901;
   reg _417902_417902 ; 
   reg __417902_417902;
   reg _417903_417903 ; 
   reg __417903_417903;
   reg _417904_417904 ; 
   reg __417904_417904;
   reg _417905_417905 ; 
   reg __417905_417905;
   reg _417906_417906 ; 
   reg __417906_417906;
   reg _417907_417907 ; 
   reg __417907_417907;
   reg _417908_417908 ; 
   reg __417908_417908;
   reg _417909_417909 ; 
   reg __417909_417909;
   reg _417910_417910 ; 
   reg __417910_417910;
   reg _417911_417911 ; 
   reg __417911_417911;
   reg _417912_417912 ; 
   reg __417912_417912;
   reg _417913_417913 ; 
   reg __417913_417913;
   reg _417914_417914 ; 
   reg __417914_417914;
   reg _417915_417915 ; 
   reg __417915_417915;
   reg _417916_417916 ; 
   reg __417916_417916;
   reg _417917_417917 ; 
   reg __417917_417917;
   reg _417918_417918 ; 
   reg __417918_417918;
   reg _417919_417919 ; 
   reg __417919_417919;
   reg _417920_417920 ; 
   reg __417920_417920;
   reg _417921_417921 ; 
   reg __417921_417921;
   reg _417922_417922 ; 
   reg __417922_417922;
   reg _417923_417923 ; 
   reg __417923_417923;
   reg _417924_417924 ; 
   reg __417924_417924;
   reg _417925_417925 ; 
   reg __417925_417925;
   reg _417926_417926 ; 
   reg __417926_417926;
   reg _417927_417927 ; 
   reg __417927_417927;
   reg _417928_417928 ; 
   reg __417928_417928;
   reg _417929_417929 ; 
   reg __417929_417929;
   reg _417930_417930 ; 
   reg __417930_417930;
   reg _417931_417931 ; 
   reg __417931_417931;
   reg _417932_417932 ; 
   reg __417932_417932;
   reg _417933_417933 ; 
   reg __417933_417933;
   reg _417934_417934 ; 
   reg __417934_417934;
   reg _417935_417935 ; 
   reg __417935_417935;
   reg _417936_417936 ; 
   reg __417936_417936;
   reg _417937_417937 ; 
   reg __417937_417937;
   reg _417938_417938 ; 
   reg __417938_417938;
   reg _417939_417939 ; 
   reg __417939_417939;
   reg _417940_417940 ; 
   reg __417940_417940;
   reg _417941_417941 ; 
   reg __417941_417941;
   reg _417942_417942 ; 
   reg __417942_417942;
   reg _417943_417943 ; 
   reg __417943_417943;
   reg _417944_417944 ; 
   reg __417944_417944;
   reg _417945_417945 ; 
   reg __417945_417945;
   reg _417946_417946 ; 
   reg __417946_417946;
   reg _417947_417947 ; 
   reg __417947_417947;
   reg _417948_417948 ; 
   reg __417948_417948;
   reg _417949_417949 ; 
   reg __417949_417949;
   reg _417950_417950 ; 
   reg __417950_417950;
   reg _417951_417951 ; 
   reg __417951_417951;
   reg _417952_417952 ; 
   reg __417952_417952;
   reg _417953_417953 ; 
   reg __417953_417953;
   reg _417954_417954 ; 
   reg __417954_417954;
   reg _417955_417955 ; 
   reg __417955_417955;
   reg _417956_417956 ; 
   reg __417956_417956;
   reg _417957_417957 ; 
   reg __417957_417957;
   reg _417958_417958 ; 
   reg __417958_417958;
   reg _417959_417959 ; 
   reg __417959_417959;
   reg _417960_417960 ; 
   reg __417960_417960;
   reg _417961_417961 ; 
   reg __417961_417961;
   reg _417962_417962 ; 
   reg __417962_417962;
   reg _417963_417963 ; 
   reg __417963_417963;
   reg _417964_417964 ; 
   reg __417964_417964;
   reg _417965_417965 ; 
   reg __417965_417965;
   reg _417966_417966 ; 
   reg __417966_417966;
   reg _417967_417967 ; 
   reg __417967_417967;
   reg _417968_417968 ; 
   reg __417968_417968;
   reg _417969_417969 ; 
   reg __417969_417969;
   reg _417970_417970 ; 
   reg __417970_417970;
   reg _417971_417971 ; 
   reg __417971_417971;
   reg _417972_417972 ; 
   reg __417972_417972;
   reg _417973_417973 ; 
   reg __417973_417973;
   reg _417974_417974 ; 
   reg __417974_417974;
   reg _417975_417975 ; 
   reg __417975_417975;
   reg _417976_417976 ; 
   reg __417976_417976;
   reg _417977_417977 ; 
   reg __417977_417977;
   reg _417978_417978 ; 
   reg __417978_417978;
   reg _417979_417979 ; 
   reg __417979_417979;
   reg _417980_417980 ; 
   reg __417980_417980;
   reg _417981_417981 ; 
   reg __417981_417981;
   reg _417982_417982 ; 
   reg __417982_417982;
   reg _417983_417983 ; 
   reg __417983_417983;
   reg _417984_417984 ; 
   reg __417984_417984;
   reg _417985_417985 ; 
   reg __417985_417985;
   reg _417986_417986 ; 
   reg __417986_417986;
   reg _417987_417987 ; 
   reg __417987_417987;
   reg _417988_417988 ; 
   reg __417988_417988;
   reg _417989_417989 ; 
   reg __417989_417989;
   reg _417990_417990 ; 
   reg __417990_417990;
   reg _417991_417991 ; 
   reg __417991_417991;
   reg _417992_417992 ; 
   reg __417992_417992;
   reg _417993_417993 ; 
   reg __417993_417993;
   reg _417994_417994 ; 
   reg __417994_417994;
   reg _417995_417995 ; 
   reg __417995_417995;
   reg _417996_417996 ; 
   reg __417996_417996;
   reg _417997_417997 ; 
   reg __417997_417997;
   reg _417998_417998 ; 
   reg __417998_417998;
   reg _417999_417999 ; 
   reg __417999_417999;
   reg _418000_418000 ; 
   reg __418000_418000;
   reg _418001_418001 ; 
   reg __418001_418001;
   reg _418002_418002 ; 
   reg __418002_418002;
   reg _418003_418003 ; 
   reg __418003_418003;
   reg _418004_418004 ; 
   reg __418004_418004;
   reg _418005_418005 ; 
   reg __418005_418005;
   reg _418006_418006 ; 
   reg __418006_418006;
   reg _418007_418007 ; 
   reg __418007_418007;
   reg _418008_418008 ; 
   reg __418008_418008;
   reg _418009_418009 ; 
   reg __418009_418009;
   reg _418010_418010 ; 
   reg __418010_418010;
   reg _418011_418011 ; 
   reg __418011_418011;
   reg _418012_418012 ; 
   reg __418012_418012;
   reg _418013_418013 ; 
   reg __418013_418013;
   reg _418014_418014 ; 
   reg __418014_418014;
   reg _418015_418015 ; 
   reg __418015_418015;
   reg _418016_418016 ; 
   reg __418016_418016;
   reg _418017_418017 ; 
   reg __418017_418017;
   reg _418018_418018 ; 
   reg __418018_418018;
   reg _418019_418019 ; 
   reg __418019_418019;
   reg _418020_418020 ; 
   reg __418020_418020;
   reg _418021_418021 ; 
   reg __418021_418021;
   reg _418022_418022 ; 
   reg __418022_418022;
   reg _418023_418023 ; 
   reg __418023_418023;
   reg _418024_418024 ; 
   reg __418024_418024;
   reg _418025_418025 ; 
   reg __418025_418025;
   reg _418026_418026 ; 
   reg __418026_418026;
   reg _418027_418027 ; 
   reg __418027_418027;
   reg _418028_418028 ; 
   reg __418028_418028;
   reg _418029_418029 ; 
   reg __418029_418029;
   reg _418030_418030 ; 
   reg __418030_418030;
   reg _418031_418031 ; 
   reg __418031_418031;
   reg _418032_418032 ; 
   reg __418032_418032;
   reg _418033_418033 ; 
   reg __418033_418033;
   reg _418034_418034 ; 
   reg __418034_418034;
   reg _418035_418035 ; 
   reg __418035_418035;
   reg _418036_418036 ; 
   reg __418036_418036;
   reg _418037_418037 ; 
   reg __418037_418037;
   reg _418038_418038 ; 
   reg __418038_418038;
   reg _418039_418039 ; 
   reg __418039_418039;
   reg _418040_418040 ; 
   reg __418040_418040;
   reg _418041_418041 ; 
   reg __418041_418041;
   reg _418042_418042 ; 
   reg __418042_418042;
   reg _418043_418043 ; 
   reg __418043_418043;
   reg _418044_418044 ; 
   reg __418044_418044;
   reg _418045_418045 ; 
   reg __418045_418045;
   reg _418046_418046 ; 
   reg __418046_418046;
   reg _418047_418047 ; 
   reg __418047_418047;
   reg _418048_418048 ; 
   reg __418048_418048;
   reg _418049_418049 ; 
   reg __418049_418049;
   reg _418050_418050 ; 
   reg __418050_418050;
   reg _418051_418051 ; 
   reg __418051_418051;
   reg _418052_418052 ; 
   reg __418052_418052;
   reg _418053_418053 ; 
   reg __418053_418053;
   reg _418054_418054 ; 
   reg __418054_418054;
   reg _418055_418055 ; 
   reg __418055_418055;
   reg _418056_418056 ; 
   reg __418056_418056;
   reg _418057_418057 ; 
   reg __418057_418057;
   reg _418058_418058 ; 
   reg __418058_418058;
   reg _418059_418059 ; 
   reg __418059_418059;
   reg _418060_418060 ; 
   reg __418060_418060;
   reg _418061_418061 ; 
   reg __418061_418061;
   reg _418062_418062 ; 
   reg __418062_418062;
   reg _418063_418063 ; 
   reg __418063_418063;
   reg _418064_418064 ; 
   reg __418064_418064;
   reg _418065_418065 ; 
   reg __418065_418065;
   reg _418066_418066 ; 
   reg __418066_418066;
   reg _418067_418067 ; 
   reg __418067_418067;
   reg _418068_418068 ; 
   reg __418068_418068;
   reg _418069_418069 ; 
   reg __418069_418069;
   reg _418070_418070 ; 
   reg __418070_418070;
   reg _418071_418071 ; 
   reg __418071_418071;
   reg _418072_418072 ; 
   reg __418072_418072;
   reg _418073_418073 ; 
   reg __418073_418073;
   reg _418074_418074 ; 
   reg __418074_418074;
   reg _418075_418075 ; 
   reg __418075_418075;
   reg _418076_418076 ; 
   reg __418076_418076;
   reg _418077_418077 ; 
   reg __418077_418077;
   reg _418078_418078 ; 
   reg __418078_418078;
   reg _418079_418079 ; 
   reg __418079_418079;
   reg _418080_418080 ; 
   reg __418080_418080;
   reg _418081_418081 ; 
   reg __418081_418081;
   reg _418082_418082 ; 
   reg __418082_418082;
   reg _418083_418083 ; 
   reg __418083_418083;
   reg _418084_418084 ; 
   reg __418084_418084;
   reg _418085_418085 ; 
   reg __418085_418085;
   reg _418086_418086 ; 
   reg __418086_418086;
   reg _418087_418087 ; 
   reg __418087_418087;
   reg _418088_418088 ; 
   reg __418088_418088;
   reg _418089_418089 ; 
   reg __418089_418089;
   reg _418090_418090 ; 
   reg __418090_418090;
   reg _418091_418091 ; 
   reg __418091_418091;
   reg _418092_418092 ; 
   reg __418092_418092;
   reg _418093_418093 ; 
   reg __418093_418093;
   reg _418094_418094 ; 
   reg __418094_418094;
   reg _418095_418095 ; 
   reg __418095_418095;
   reg _418096_418096 ; 
   reg __418096_418096;
   reg _418097_418097 ; 
   reg __418097_418097;
   reg _418098_418098 ; 
   reg __418098_418098;
   reg _418099_418099 ; 
   reg __418099_418099;
   reg _418100_418100 ; 
   reg __418100_418100;
   reg _418101_418101 ; 
   reg __418101_418101;
   reg _418102_418102 ; 
   reg __418102_418102;
   reg _418103_418103 ; 
   reg __418103_418103;
   reg _418104_418104 ; 
   reg __418104_418104;
   reg _418105_418105 ; 
   reg __418105_418105;
   reg _418106_418106 ; 
   reg __418106_418106;
   reg _418107_418107 ; 
   reg __418107_418107;
   reg _418108_418108 ; 
   reg __418108_418108;
   reg _418109_418109 ; 
   reg __418109_418109;
   reg _418110_418110 ; 
   reg __418110_418110;
   reg _418111_418111 ; 
   reg __418111_418111;
   reg _418112_418112 ; 
   reg __418112_418112;
   reg _418113_418113 ; 
   reg __418113_418113;
   reg _418114_418114 ; 
   reg __418114_418114;
   reg _418115_418115 ; 
   reg __418115_418115;
   reg _418116_418116 ; 
   reg __418116_418116;
   reg _418117_418117 ; 
   reg __418117_418117;
   reg _418118_418118 ; 
   reg __418118_418118;
   reg _418119_418119 ; 
   reg __418119_418119;
   reg _418120_418120 ; 
   reg __418120_418120;
   reg _418121_418121 ; 
   reg __418121_418121;
   reg _418122_418122 ; 
   reg __418122_418122;
   reg _418123_418123 ; 
   reg __418123_418123;
   reg _418124_418124 ; 
   reg __418124_418124;
   reg _418125_418125 ; 
   reg __418125_418125;
   reg _418126_418126 ; 
   reg __418126_418126;
   reg _418127_418127 ; 
   reg __418127_418127;
   reg _418128_418128 ; 
   reg __418128_418128;
   reg _418129_418129 ; 
   reg __418129_418129;
   reg _418130_418130 ; 
   reg __418130_418130;
   reg _418131_418131 ; 
   reg __418131_418131;
   reg _418132_418132 ; 
   reg __418132_418132;
   reg _418133_418133 ; 
   reg __418133_418133;
   reg _418134_418134 ; 
   reg __418134_418134;
   reg _418135_418135 ; 
   reg __418135_418135;
   reg _418136_418136 ; 
   reg __418136_418136;
   reg _418137_418137 ; 
   reg __418137_418137;
   reg _418138_418138 ; 
   reg __418138_418138;
   reg _418139_418139 ; 
   reg __418139_418139;
   reg _418140_418140 ; 
   reg __418140_418140;
   reg _418141_418141 ; 
   reg __418141_418141;
   reg _418142_418142 ; 
   reg __418142_418142;
   reg _418143_418143 ; 
   reg __418143_418143;
   reg _418144_418144 ; 
   reg __418144_418144;
   reg _418145_418145 ; 
   reg __418145_418145;
   reg _418146_418146 ; 
   reg __418146_418146;
   reg _418147_418147 ; 
   reg __418147_418147;
   reg _418148_418148 ; 
   reg __418148_418148;
   reg _418149_418149 ; 
   reg __418149_418149;
   reg _418150_418150 ; 
   reg __418150_418150;
   reg _418151_418151 ; 
   reg __418151_418151;
   reg _418152_418152 ; 
   reg __418152_418152;
   reg _418153_418153 ; 
   reg __418153_418153;
   reg _418154_418154 ; 
   reg __418154_418154;
   reg _418155_418155 ; 
   reg __418155_418155;
   reg _418156_418156 ; 
   reg __418156_418156;
   reg _418157_418157 ; 
   reg __418157_418157;
   reg _418158_418158 ; 
   reg __418158_418158;
   reg _418159_418159 ; 
   reg __418159_418159;
   reg _418160_418160 ; 
   reg __418160_418160;
   reg _418161_418161 ; 
   reg __418161_418161;
   reg _418162_418162 ; 
   reg __418162_418162;
   reg _418163_418163 ; 
   reg __418163_418163;
   reg _418164_418164 ; 
   reg __418164_418164;
   reg _418165_418165 ; 
   reg __418165_418165;
   reg _418166_418166 ; 
   reg __418166_418166;
   reg _418167_418167 ; 
   reg __418167_418167;
   reg _418168_418168 ; 
   reg __418168_418168;
   reg _418169_418169 ; 
   reg __418169_418169;
   reg _418170_418170 ; 
   reg __418170_418170;
   reg _418171_418171 ; 
   reg __418171_418171;
   reg _418172_418172 ; 
   reg __418172_418172;
   reg _418173_418173 ; 
   reg __418173_418173;
   reg _418174_418174 ; 
   reg __418174_418174;
   reg _418175_418175 ; 
   reg __418175_418175;
   reg _418176_418176 ; 
   reg __418176_418176;
   reg _418177_418177 ; 
   reg __418177_418177;
   reg _418178_418178 ; 
   reg __418178_418178;
   reg _418179_418179 ; 
   reg __418179_418179;
   reg _418180_418180 ; 
   reg __418180_418180;
   reg _418181_418181 ; 
   reg __418181_418181;
   reg _418182_418182 ; 
   reg __418182_418182;
   reg _418183_418183 ; 
   reg __418183_418183;
   reg _418184_418184 ; 
   reg __418184_418184;
   reg _418185_418185 ; 
   reg __418185_418185;
   reg _418186_418186 ; 
   reg __418186_418186;
   reg _418187_418187 ; 
   reg __418187_418187;
   reg _418188_418188 ; 
   reg __418188_418188;
   reg _418189_418189 ; 
   reg __418189_418189;
   reg _418190_418190 ; 
   reg __418190_418190;
   reg _418191_418191 ; 
   reg __418191_418191;
   reg _418192_418192 ; 
   reg __418192_418192;
   reg _418193_418193 ; 
   reg __418193_418193;
   reg _418194_418194 ; 
   reg __418194_418194;
   reg _418195_418195 ; 
   reg __418195_418195;
   reg _418196_418196 ; 
   reg __418196_418196;
   reg _418197_418197 ; 
   reg __418197_418197;
   reg _418198_418198 ; 
   reg __418198_418198;
   reg _418199_418199 ; 
   reg __418199_418199;
   reg _418200_418200 ; 
   reg __418200_418200;
   reg _418201_418201 ; 
   reg __418201_418201;
   reg _418202_418202 ; 
   reg __418202_418202;
   reg _418203_418203 ; 
   reg __418203_418203;
   reg _418204_418204 ; 
   reg __418204_418204;
   reg _418205_418205 ; 
   reg __418205_418205;
   reg _418206_418206 ; 
   reg __418206_418206;
   reg _418207_418207 ; 
   reg __418207_418207;
   reg _418208_418208 ; 
   reg __418208_418208;
   reg _418209_418209 ; 
   reg __418209_418209;
   reg _418210_418210 ; 
   reg __418210_418210;
   reg _418211_418211 ; 
   reg __418211_418211;
   reg _418212_418212 ; 
   reg __418212_418212;
   reg _418213_418213 ; 
   reg __418213_418213;
   reg _418214_418214 ; 
   reg __418214_418214;
   reg _418215_418215 ; 
   reg __418215_418215;
   reg _418216_418216 ; 
   reg __418216_418216;
   reg _418217_418217 ; 
   reg __418217_418217;
   reg _418218_418218 ; 
   reg __418218_418218;
   reg _418219_418219 ; 
   reg __418219_418219;
   reg _418220_418220 ; 
   reg __418220_418220;
   reg _418221_418221 ; 
   reg __418221_418221;
   reg _418222_418222 ; 
   reg __418222_418222;
   reg _418223_418223 ; 
   reg __418223_418223;
   reg _418224_418224 ; 
   reg __418224_418224;
   reg _418225_418225 ; 
   reg __418225_418225;
   reg _418226_418226 ; 
   reg __418226_418226;
   reg _418227_418227 ; 
   reg __418227_418227;
   reg _418228_418228 ; 
   reg __418228_418228;
   reg _418229_418229 ; 
   reg __418229_418229;
   reg _418230_418230 ; 
   reg __418230_418230;
   reg _418231_418231 ; 
   reg __418231_418231;
   reg _418232_418232 ; 
   reg __418232_418232;
   reg _418233_418233 ; 
   reg __418233_418233;
   reg _418234_418234 ; 
   reg __418234_418234;
   reg _418235_418235 ; 
   reg __418235_418235;
   reg _418236_418236 ; 
   reg __418236_418236;
   reg _418237_418237 ; 
   reg __418237_418237;
   reg _418238_418238 ; 
   reg __418238_418238;
   reg _418239_418239 ; 
   reg __418239_418239;
   reg _418240_418240 ; 
   reg __418240_418240;
   reg _418241_418241 ; 
   reg __418241_418241;
   reg _418242_418242 ; 
   reg __418242_418242;
   reg _418243_418243 ; 
   reg __418243_418243;
   reg _418244_418244 ; 
   reg __418244_418244;
   reg _418245_418245 ; 
   reg __418245_418245;
   reg _418246_418246 ; 
   reg __418246_418246;
   reg _418247_418247 ; 
   reg __418247_418247;
   reg _418248_418248 ; 
   reg __418248_418248;
   reg _418249_418249 ; 
   reg __418249_418249;
   reg _418250_418250 ; 
   reg __418250_418250;
   reg _418251_418251 ; 
   reg __418251_418251;
   reg _418252_418252 ; 
   reg __418252_418252;
   reg _418253_418253 ; 
   reg __418253_418253;
   reg _418254_418254 ; 
   reg __418254_418254;
   reg _418255_418255 ; 
   reg __418255_418255;
   reg _418256_418256 ; 
   reg __418256_418256;
   reg _418257_418257 ; 
   reg __418257_418257;
   reg _418258_418258 ; 
   reg __418258_418258;
   reg _418259_418259 ; 
   reg __418259_418259;
   reg _418260_418260 ; 
   reg __418260_418260;
   reg _418261_418261 ; 
   reg __418261_418261;
   reg _418262_418262 ; 
   reg __418262_418262;
   reg _418263_418263 ; 
   reg __418263_418263;
   reg _418264_418264 ; 
   reg __418264_418264;
   reg _418265_418265 ; 
   reg __418265_418265;
   reg _418266_418266 ; 
   reg __418266_418266;
   reg _418267_418267 ; 
   reg __418267_418267;
   reg _418268_418268 ; 
   reg __418268_418268;
   reg _418269_418269 ; 
   reg __418269_418269;
   reg _418270_418270 ; 
   reg __418270_418270;
   reg _418271_418271 ; 
   reg __418271_418271;
   reg _418272_418272 ; 
   reg __418272_418272;
   reg _418273_418273 ; 
   reg __418273_418273;
   reg _418274_418274 ; 
   reg __418274_418274;
   reg _418275_418275 ; 
   reg __418275_418275;
   reg _418276_418276 ; 
   reg __418276_418276;
   reg _418277_418277 ; 
   reg __418277_418277;
   reg _418278_418278 ; 
   reg __418278_418278;
   reg _418279_418279 ; 
   reg __418279_418279;
   reg _418280_418280 ; 
   reg __418280_418280;
   reg _418281_418281 ; 
   reg __418281_418281;
   reg _418282_418282 ; 
   reg __418282_418282;
   reg _418283_418283 ; 
   reg __418283_418283;
   reg _418284_418284 ; 
   reg __418284_418284;
   reg _418285_418285 ; 
   reg __418285_418285;
   reg _418286_418286 ; 
   reg __418286_418286;
   reg _418287_418287 ; 
   reg __418287_418287;
   reg _418288_418288 ; 
   reg __418288_418288;
   reg _418289_418289 ; 
   reg __418289_418289;
   reg _418290_418290 ; 
   reg __418290_418290;
   reg _418291_418291 ; 
   reg __418291_418291;
   reg _418292_418292 ; 
   reg __418292_418292;
   reg _418293_418293 ; 
   reg __418293_418293;
   reg _418294_418294 ; 
   reg __418294_418294;
   reg _418295_418295 ; 
   reg __418295_418295;
   reg _418296_418296 ; 
   reg __418296_418296;
   reg _418297_418297 ; 
   reg __418297_418297;
   reg _418298_418298 ; 
   reg __418298_418298;
   reg _418299_418299 ; 
   reg __418299_418299;
   reg _418300_418300 ; 
   reg __418300_418300;
   reg _418301_418301 ; 
   reg __418301_418301;
   reg _418302_418302 ; 
   reg __418302_418302;
   reg _418303_418303 ; 
   reg __418303_418303;
   reg _418304_418304 ; 
   reg __418304_418304;
   reg _418305_418305 ; 
   reg __418305_418305;
   reg _418306_418306 ; 
   reg __418306_418306;
   reg _418307_418307 ; 
   reg __418307_418307;
   reg _418308_418308 ; 
   reg __418308_418308;
   reg _418309_418309 ; 
   reg __418309_418309;
   reg _418310_418310 ; 
   reg __418310_418310;
   reg _418311_418311 ; 
   reg __418311_418311;
   reg _418312_418312 ; 
   reg __418312_418312;
   reg _418313_418313 ; 
   reg __418313_418313;
   reg _418314_418314 ; 
   reg __418314_418314;
   reg _418315_418315 ; 
   reg __418315_418315;
   reg _418316_418316 ; 
   reg __418316_418316;
   reg _418317_418317 ; 
   reg __418317_418317;
   reg _418318_418318 ; 
   reg __418318_418318;
   reg _418319_418319 ; 
   reg __418319_418319;
   reg _418320_418320 ; 
   reg __418320_418320;
   reg _418321_418321 ; 
   reg __418321_418321;
   reg _418322_418322 ; 
   reg __418322_418322;
   reg _418323_418323 ; 
   reg __418323_418323;
   reg _418324_418324 ; 
   reg __418324_418324;
   reg _418325_418325 ; 
   reg __418325_418325;
   reg _418326_418326 ; 
   reg __418326_418326;
   reg _418327_418327 ; 
   reg __418327_418327;
   reg _418328_418328 ; 
   reg __418328_418328;
   reg _418329_418329 ; 
   reg __418329_418329;
   reg _418330_418330 ; 
   reg __418330_418330;
   reg _418331_418331 ; 
   reg __418331_418331;
   reg _418332_418332 ; 
   reg __418332_418332;
   reg _418333_418333 ; 
   reg __418333_418333;
   reg _418334_418334 ; 
   reg __418334_418334;
   reg _418335_418335 ; 
   reg __418335_418335;
   reg _418336_418336 ; 
   reg __418336_418336;
   reg _418337_418337 ; 
   reg __418337_418337;
   reg _418338_418338 ; 
   reg __418338_418338;
   reg _418339_418339 ; 
   reg __418339_418339;
   reg _418340_418340 ; 
   reg __418340_418340;
   reg _418341_418341 ; 
   reg __418341_418341;
   reg _418342_418342 ; 
   reg __418342_418342;
   reg _418343_418343 ; 
   reg __418343_418343;
   reg _418344_418344 ; 
   reg __418344_418344;
   reg _418345_418345 ; 
   reg __418345_418345;
   reg _418346_418346 ; 
   reg __418346_418346;
   reg _418347_418347 ; 
   reg __418347_418347;
   reg _418348_418348 ; 
   reg __418348_418348;
   reg _418349_418349 ; 
   reg __418349_418349;
   reg _418350_418350 ; 
   reg __418350_418350;
   reg _418351_418351 ; 
   reg __418351_418351;
   reg _418352_418352 ; 
   reg __418352_418352;
   reg _418353_418353 ; 
   reg __418353_418353;
   reg _418354_418354 ; 
   reg __418354_418354;
   reg _418355_418355 ; 
   reg __418355_418355;
   reg _418356_418356 ; 
   reg __418356_418356;
   reg _418357_418357 ; 
   reg __418357_418357;
   reg _418358_418358 ; 
   reg __418358_418358;
   reg _418359_418359 ; 
   reg __418359_418359;
   reg _418360_418360 ; 
   reg __418360_418360;
   reg _418361_418361 ; 
   reg __418361_418361;
   reg _418362_418362 ; 
   reg __418362_418362;
   reg _418363_418363 ; 
   reg __418363_418363;
   reg _418364_418364 ; 
   reg __418364_418364;
   reg _418365_418365 ; 
   reg __418365_418365;
   reg _418366_418366 ; 
   reg __418366_418366;
   reg _418367_418367 ; 
   reg __418367_418367;
   reg _418368_418368 ; 
   reg __418368_418368;
   reg _418369_418369 ; 
   reg __418369_418369;
   reg _418370_418370 ; 
   reg __418370_418370;
   reg _418371_418371 ; 
   reg __418371_418371;
   reg _418372_418372 ; 
   reg __418372_418372;
   reg _418373_418373 ; 
   reg __418373_418373;
   reg _418374_418374 ; 
   reg __418374_418374;
   reg _418375_418375 ; 
   reg __418375_418375;
   reg _418376_418376 ; 
   reg __418376_418376;
   reg _418377_418377 ; 
   reg __418377_418377;
   reg _418378_418378 ; 
   reg __418378_418378;
   reg _418379_418379 ; 
   reg __418379_418379;
   reg _418380_418380 ; 
   reg __418380_418380;
   reg _418381_418381 ; 
   reg __418381_418381;
   reg _418382_418382 ; 
   reg __418382_418382;
   reg _418383_418383 ; 
   reg __418383_418383;
   reg _418384_418384 ; 
   reg __418384_418384;
   reg _418385_418385 ; 
   reg __418385_418385;
   reg _418386_418386 ; 
   reg __418386_418386;
   reg _418387_418387 ; 
   reg __418387_418387;
   reg _418388_418388 ; 
   reg __418388_418388;
   reg _418389_418389 ; 
   reg __418389_418389;
   reg _418390_418390 ; 
   reg __418390_418390;
   reg _418391_418391 ; 
   reg __418391_418391;
   reg _418392_418392 ; 
   reg __418392_418392;
   reg _418393_418393 ; 
   reg __418393_418393;
   reg _418394_418394 ; 
   reg __418394_418394;
   reg _418395_418395 ; 
   reg __418395_418395;
   reg _418396_418396 ; 
   reg __418396_418396;
   reg _418397_418397 ; 
   reg __418397_418397;
   reg _418398_418398 ; 
   reg __418398_418398;
   reg _418399_418399 ; 
   reg __418399_418399;
   reg _418400_418400 ; 
   reg __418400_418400;
   reg _418401_418401 ; 
   reg __418401_418401;
   reg _418402_418402 ; 
   reg __418402_418402;
   reg _418403_418403 ; 
   reg __418403_418403;
   reg _418404_418404 ; 
   reg __418404_418404;
   reg _418405_418405 ; 
   reg __418405_418405;
   reg _418406_418406 ; 
   reg __418406_418406;
   reg _418407_418407 ; 
   reg __418407_418407;
   reg _418408_418408 ; 
   reg __418408_418408;
   reg _418409_418409 ; 
   reg __418409_418409;
   reg _418410_418410 ; 
   reg __418410_418410;
   reg _418411_418411 ; 
   reg __418411_418411;
   reg _418412_418412 ; 
   reg __418412_418412;
   reg _418413_418413 ; 
   reg __418413_418413;
   reg _418414_418414 ; 
   reg __418414_418414;
   reg _418415_418415 ; 
   reg __418415_418415;
   reg _418416_418416 ; 
   reg __418416_418416;
   reg _418417_418417 ; 
   reg __418417_418417;
   reg _418418_418418 ; 
   reg __418418_418418;
   reg _418419_418419 ; 
   reg __418419_418419;
   reg _418420_418420 ; 
   reg __418420_418420;
   reg _418421_418421 ; 
   reg __418421_418421;
   reg _418422_418422 ; 
   reg __418422_418422;
   reg _418423_418423 ; 
   reg __418423_418423;
   reg _418424_418424 ; 
   reg __418424_418424;
   reg _418425_418425 ; 
   reg __418425_418425;
   reg _418426_418426 ; 
   reg __418426_418426;
   reg _418427_418427 ; 
   reg __418427_418427;
   reg _418428_418428 ; 
   reg __418428_418428;
   reg _418429_418429 ; 
   reg __418429_418429;
   reg _418430_418430 ; 
   reg __418430_418430;
   reg _418431_418431 ; 
   reg __418431_418431;
   reg _418432_418432 ; 
   reg __418432_418432;
   reg _418433_418433 ; 
   reg __418433_418433;
   reg _418434_418434 ; 
   reg __418434_418434;
   reg _418435_418435 ; 
   reg __418435_418435;
   reg _418436_418436 ; 
   reg __418436_418436;
   reg _418437_418437 ; 
   reg __418437_418437;
   reg _418438_418438 ; 
   reg __418438_418438;
   reg _418439_418439 ; 
   reg __418439_418439;
   reg _418440_418440 ; 
   reg __418440_418440;
   reg _418441_418441 ; 
   reg __418441_418441;
   reg _418442_418442 ; 
   reg __418442_418442;
   reg _418443_418443 ; 
   reg __418443_418443;
   reg _418444_418444 ; 
   reg __418444_418444;
   reg _418445_418445 ; 
   reg __418445_418445;
   reg _418446_418446 ; 
   reg __418446_418446;
   reg _418447_418447 ; 
   reg __418447_418447;
   reg _418448_418448 ; 
   reg __418448_418448;
   reg _418449_418449 ; 
   reg __418449_418449;
   reg _418450_418450 ; 
   reg __418450_418450;
   reg _418451_418451 ; 
   reg __418451_418451;
   reg _418452_418452 ; 
   reg __418452_418452;
   reg _418453_418453 ; 
   reg __418453_418453;
   reg _418454_418454 ; 
   reg __418454_418454;
   reg _418455_418455 ; 
   reg __418455_418455;
   reg _418456_418456 ; 
   reg __418456_418456;
   reg _418457_418457 ; 
   reg __418457_418457;
   reg _418458_418458 ; 
   reg __418458_418458;
   reg _418459_418459 ; 
   reg __418459_418459;
   reg _418460_418460 ; 
   reg __418460_418460;
   reg _418461_418461 ; 
   reg __418461_418461;
   reg _418462_418462 ; 
   reg __418462_418462;
   reg _418463_418463 ; 
   reg __418463_418463;
   reg _418464_418464 ; 
   reg __418464_418464;
   reg _418465_418465 ; 
   reg __418465_418465;
   reg _418466_418466 ; 
   reg __418466_418466;
   reg _418467_418467 ; 
   reg __418467_418467;
   reg _418468_418468 ; 
   reg __418468_418468;
   reg _418469_418469 ; 
   reg __418469_418469;
   reg _418470_418470 ; 
   reg __418470_418470;
   reg _418471_418471 ; 
   reg __418471_418471;
   reg _418472_418472 ; 
   reg __418472_418472;
   reg _418473_418473 ; 
   reg __418473_418473;
   reg _418474_418474 ; 
   reg __418474_418474;
   reg _418475_418475 ; 
   reg __418475_418475;
   reg _418476_418476 ; 
   reg __418476_418476;
   reg _418477_418477 ; 
   reg __418477_418477;
   reg _418478_418478 ; 
   reg __418478_418478;
   reg _418479_418479 ; 
   reg __418479_418479;
   reg _418480_418480 ; 
   reg __418480_418480;
   reg _418481_418481 ; 
   reg __418481_418481;
   reg _418482_418482 ; 
   reg __418482_418482;
   reg _418483_418483 ; 
   reg __418483_418483;
   reg _418484_418484 ; 
   reg __418484_418484;
   reg _418485_418485 ; 
   reg __418485_418485;
   reg _418486_418486 ; 
   reg __418486_418486;
   reg _418487_418487 ; 
   reg __418487_418487;
   reg _418488_418488 ; 
   reg __418488_418488;
   reg _418489_418489 ; 
   reg __418489_418489;
   reg _418490_418490 ; 
   reg __418490_418490;
   reg _418491_418491 ; 
   reg __418491_418491;
   reg _418492_418492 ; 
   reg __418492_418492;
   reg _418493_418493 ; 
   reg __418493_418493;
   reg _418494_418494 ; 
   reg __418494_418494;
   reg _418495_418495 ; 
   reg __418495_418495;
   reg _418496_418496 ; 
   reg __418496_418496;
   reg _418497_418497 ; 
   reg __418497_418497;
   reg _418498_418498 ; 
   reg __418498_418498;
   reg _418499_418499 ; 
   reg __418499_418499;
   reg _418500_418500 ; 
   reg __418500_418500;
   reg _418501_418501 ; 
   reg __418501_418501;
   reg _418502_418502 ; 
   reg __418502_418502;
   reg _418503_418503 ; 
   reg __418503_418503;
   reg _418504_418504 ; 
   reg __418504_418504;
   reg _418505_418505 ; 
   reg __418505_418505;
   reg _418506_418506 ; 
   reg __418506_418506;
   reg _418507_418507 ; 
   reg __418507_418507;
   reg _418508_418508 ; 
   reg __418508_418508;
   reg _418509_418509 ; 
   reg __418509_418509;
   reg _418510_418510 ; 
   reg __418510_418510;
   reg _418511_418511 ; 
   reg __418511_418511;
   reg _418512_418512 ; 
   reg __418512_418512;
   reg _418513_418513 ; 
   reg __418513_418513;
   reg _418514_418514 ; 
   reg __418514_418514;
   reg _418515_418515 ; 
   reg __418515_418515;
   reg _418516_418516 ; 
   reg __418516_418516;
   reg _418517_418517 ; 
   reg __418517_418517;
   reg _418518_418518 ; 
   reg __418518_418518;
   reg _418519_418519 ; 
   reg __418519_418519;
   reg _418520_418520 ; 
   reg __418520_418520;
   reg _418521_418521 ; 
   reg __418521_418521;
   reg _418522_418522 ; 
   reg __418522_418522;
   reg _418523_418523 ; 
   reg __418523_418523;
   reg _418524_418524 ; 
   reg __418524_418524;
   reg _418525_418525 ; 
   reg __418525_418525;
   reg _418526_418526 ; 
   reg __418526_418526;
   reg _418527_418527 ; 
   reg __418527_418527;
   reg _418528_418528 ; 
   reg __418528_418528;
   reg _418529_418529 ; 
   reg __418529_418529;
   reg _418530_418530 ; 
   reg __418530_418530;
   reg _418531_418531 ; 
   reg __418531_418531;
   reg _418532_418532 ; 
   reg __418532_418532;
   reg _418533_418533 ; 
   reg __418533_418533;
   reg _418534_418534 ; 
   reg __418534_418534;
   reg _418535_418535 ; 
   reg __418535_418535;
   reg _418536_418536 ; 
   reg __418536_418536;
   reg _418537_418537 ; 
   reg __418537_418537;
   reg _418538_418538 ; 
   reg __418538_418538;
   reg _418539_418539 ; 
   reg __418539_418539;
   reg _418540_418540 ; 
   reg __418540_418540;
   reg _418541_418541 ; 
   reg __418541_418541;
   reg _418542_418542 ; 
   reg __418542_418542;
   reg _418543_418543 ; 
   reg __418543_418543;
   reg _418544_418544 ; 
   reg __418544_418544;
   reg _418545_418545 ; 
   reg __418545_418545;
   reg _418546_418546 ; 
   reg __418546_418546;
   reg _418547_418547 ; 
   reg __418547_418547;
   reg _418548_418548 ; 
   reg __418548_418548;
   reg _418549_418549 ; 
   reg __418549_418549;
   reg _418550_418550 ; 
   reg __418550_418550;
   reg _418551_418551 ; 
   reg __418551_418551;
   reg _418552_418552 ; 
   reg __418552_418552;
   reg _418553_418553 ; 
   reg __418553_418553;
   reg _418554_418554 ; 
   reg __418554_418554;
   reg _418555_418555 ; 
   reg __418555_418555;
   reg _418556_418556 ; 
   reg __418556_418556;
   reg _418557_418557 ; 
   reg __418557_418557;
   reg _418558_418558 ; 
   reg __418558_418558;
   reg _418559_418559 ; 
   reg __418559_418559;
   reg _418560_418560 ; 
   reg __418560_418560;
   reg _418561_418561 ; 
   reg __418561_418561;
   reg _418562_418562 ; 
   reg __418562_418562;
   reg _418563_418563 ; 
   reg __418563_418563;
   reg _418564_418564 ; 
   reg __418564_418564;
   reg _418565_418565 ; 
   reg __418565_418565;
   reg _418566_418566 ; 
   reg __418566_418566;
   reg _418567_418567 ; 
   reg __418567_418567;
   reg _418568_418568 ; 
   reg __418568_418568;
   reg _418569_418569 ; 
   reg __418569_418569;
   reg _418570_418570 ; 
   reg __418570_418570;
   reg _418571_418571 ; 
   reg __418571_418571;
   reg _418572_418572 ; 
   reg __418572_418572;
   reg _418573_418573 ; 
   reg __418573_418573;
   reg _418574_418574 ; 
   reg __418574_418574;
   reg _418575_418575 ; 
   reg __418575_418575;
   reg _418576_418576 ; 
   reg __418576_418576;
   reg _418577_418577 ; 
   reg __418577_418577;
   reg _418578_418578 ; 
   reg __418578_418578;
   reg _418579_418579 ; 
   reg __418579_418579;
   reg _418580_418580 ; 
   reg __418580_418580;
   reg _418581_418581 ; 
   reg __418581_418581;
   reg _418582_418582 ; 
   reg __418582_418582;
   reg _418583_418583 ; 
   reg __418583_418583;
   reg _418584_418584 ; 
   reg __418584_418584;
   reg _418585_418585 ; 
   reg __418585_418585;
   reg _418586_418586 ; 
   reg __418586_418586;
   reg _418587_418587 ; 
   reg __418587_418587;
   reg _418588_418588 ; 
   reg __418588_418588;
   reg _418589_418589 ; 
   reg __418589_418589;
   reg _418590_418590 ; 
   reg __418590_418590;
   reg _418591_418591 ; 
   reg __418591_418591;
   reg _418592_418592 ; 
   reg __418592_418592;
   reg _418593_418593 ; 
   reg __418593_418593;
   reg _418594_418594 ; 
   reg __418594_418594;
   reg _418595_418595 ; 
   reg __418595_418595;
   reg _418596_418596 ; 
   reg __418596_418596;
   reg _418597_418597 ; 
   reg __418597_418597;
   reg _418598_418598 ; 
   reg __418598_418598;
   reg _418599_418599 ; 
   reg __418599_418599;
   reg _418600_418600 ; 
   reg __418600_418600;
   reg _418601_418601 ; 
   reg __418601_418601;
   reg _418602_418602 ; 
   reg __418602_418602;
   reg _418603_418603 ; 
   reg __418603_418603;
   reg _418604_418604 ; 
   reg __418604_418604;
   reg _418605_418605 ; 
   reg __418605_418605;
   reg _418606_418606 ; 
   reg __418606_418606;
   reg _418607_418607 ; 
   reg __418607_418607;
   reg _418608_418608 ; 
   reg __418608_418608;
   reg _418609_418609 ; 
   reg __418609_418609;
   reg _418610_418610 ; 
   reg __418610_418610;
   reg _418611_418611 ; 
   reg __418611_418611;
   reg _418612_418612 ; 
   reg __418612_418612;
   reg _418613_418613 ; 
   reg __418613_418613;
   reg _418614_418614 ; 
   reg __418614_418614;
   reg _418615_418615 ; 
   reg __418615_418615;
   reg _418616_418616 ; 
   reg __418616_418616;
   reg _418617_418617 ; 
   reg __418617_418617;
   reg _418618_418618 ; 
   reg __418618_418618;
   reg _418619_418619 ; 
   reg __418619_418619;
   reg _418620_418620 ; 
   reg __418620_418620;
   reg _418621_418621 ; 
   reg __418621_418621;
   reg _418622_418622 ; 
   reg __418622_418622;
   reg _418623_418623 ; 
   reg __418623_418623;
   reg _418624_418624 ; 
   reg __418624_418624;
   reg _418625_418625 ; 
   reg __418625_418625;
   reg _418626_418626 ; 
   reg __418626_418626;
   reg _418627_418627 ; 
   reg __418627_418627;
   reg _418628_418628 ; 
   reg __418628_418628;
   reg _418629_418629 ; 
   reg __418629_418629;
   reg _418630_418630 ; 
   reg __418630_418630;
   reg _418631_418631 ; 
   reg __418631_418631;
   reg _418632_418632 ; 
   reg __418632_418632;
   reg _418633_418633 ; 
   reg __418633_418633;
   reg _418634_418634 ; 
   reg __418634_418634;
   reg _418635_418635 ; 
   reg __418635_418635;
   reg _418636_418636 ; 
   reg __418636_418636;
   reg _418637_418637 ; 
   reg __418637_418637;
   reg _418638_418638 ; 
   reg __418638_418638;
   reg _418639_418639 ; 
   reg __418639_418639;
   reg _418640_418640 ; 
   reg __418640_418640;
   reg _418641_418641 ; 
   reg __418641_418641;
   reg _418642_418642 ; 
   reg __418642_418642;
   reg _418643_418643 ; 
   reg __418643_418643;
   reg _418644_418644 ; 
   reg __418644_418644;
   reg _418645_418645 ; 
   reg __418645_418645;
   reg _418646_418646 ; 
   reg __418646_418646;
   reg _418647_418647 ; 
   reg __418647_418647;
   reg _418648_418648 ; 
   reg __418648_418648;
   reg _418649_418649 ; 
   reg __418649_418649;
   reg _418650_418650 ; 
   reg __418650_418650;
   reg _418651_418651 ; 
   reg __418651_418651;
   reg _418652_418652 ; 
   reg __418652_418652;
   reg _418653_418653 ; 
   reg __418653_418653;
   reg _418654_418654 ; 
   reg __418654_418654;
   reg _418655_418655 ; 
   reg __418655_418655;
   reg _418656_418656 ; 
   reg __418656_418656;
   reg _418657_418657 ; 
   reg __418657_418657;
   reg _418658_418658 ; 
   reg __418658_418658;
   reg _418659_418659 ; 
   reg __418659_418659;
   reg _418660_418660 ; 
   reg __418660_418660;
   reg _418661_418661 ; 
   reg __418661_418661;
   reg _418662_418662 ; 
   reg __418662_418662;
   reg _418663_418663 ; 
   reg __418663_418663;
   reg _418664_418664 ; 
   reg __418664_418664;
   reg _418665_418665 ; 
   reg __418665_418665;
   reg _418666_418666 ; 
   reg __418666_418666;
   reg _418667_418667 ; 
   reg __418667_418667;
   reg _418668_418668 ; 
   reg __418668_418668;
   reg _418669_418669 ; 
   reg __418669_418669;
   reg _418670_418670 ; 
   reg __418670_418670;
   reg _418671_418671 ; 
   reg __418671_418671;
   reg _418672_418672 ; 
   reg __418672_418672;
   reg _418673_418673 ; 
   reg __418673_418673;
   reg _418674_418674 ; 
   reg __418674_418674;
   reg _418675_418675 ; 
   reg __418675_418675;
   reg _418676_418676 ; 
   reg __418676_418676;
   reg _418677_418677 ; 
   reg __418677_418677;
   reg _418678_418678 ; 
   reg __418678_418678;
   reg _418679_418679 ; 
   reg __418679_418679;
   reg _418680_418680 ; 
   reg __418680_418680;
   reg _418681_418681 ; 
   reg __418681_418681;
   reg _418682_418682 ; 
   reg __418682_418682;
   reg _418683_418683 ; 
   reg __418683_418683;
   reg _418684_418684 ; 
   reg __418684_418684;
   reg _418685_418685 ; 
   reg __418685_418685;
   reg _418686_418686 ; 
   reg __418686_418686;
   reg _418687_418687 ; 
   reg __418687_418687;
   reg _418688_418688 ; 
   reg __418688_418688;
   reg _418689_418689 ; 
   reg __418689_418689;
   reg _418690_418690 ; 
   reg __418690_418690;
   reg _418691_418691 ; 
   reg __418691_418691;
   reg _418692_418692 ; 
   reg __418692_418692;
   reg _418693_418693 ; 
   reg __418693_418693;
   reg _418694_418694 ; 
   reg __418694_418694;
   reg _418695_418695 ; 
   reg __418695_418695;
   reg _418696_418696 ; 
   reg __418696_418696;
   reg _418697_418697 ; 
   reg __418697_418697;
   reg _418698_418698 ; 
   reg __418698_418698;
   reg _418699_418699 ; 
   reg __418699_418699;
   reg _418700_418700 ; 
   reg __418700_418700;
   reg _418701_418701 ; 
   reg __418701_418701;
   reg _418702_418702 ; 
   reg __418702_418702;
   reg _418703_418703 ; 
   reg __418703_418703;
   reg _418704_418704 ; 
   reg __418704_418704;
   reg _418705_418705 ; 
   reg __418705_418705;
   reg _418706_418706 ; 
   reg __418706_418706;
   reg _418707_418707 ; 
   reg __418707_418707;
   reg _418708_418708 ; 
   reg __418708_418708;
   reg _418709_418709 ; 
   reg __418709_418709;
   reg _418710_418710 ; 
   reg __418710_418710;
   reg _418711_418711 ; 
   reg __418711_418711;
   reg _418712_418712 ; 
   reg __418712_418712;
   reg _418713_418713 ; 
   reg __418713_418713;
   reg _418714_418714 ; 
   reg __418714_418714;
   reg _418715_418715 ; 
   reg __418715_418715;
   reg _418716_418716 ; 
   reg __418716_418716;
   reg _418717_418717 ; 
   reg __418717_418717;
   reg _418718_418718 ; 
   reg __418718_418718;
   reg _418719_418719 ; 
   reg __418719_418719;
   reg _418720_418720 ; 
   reg __418720_418720;
   reg _418721_418721 ; 
   reg __418721_418721;
   reg _418722_418722 ; 
   reg __418722_418722;
   reg _418723_418723 ; 
   reg __418723_418723;
   reg _418724_418724 ; 
   reg __418724_418724;
   reg _418725_418725 ; 
   reg __418725_418725;
   reg _418726_418726 ; 
   reg __418726_418726;
   reg _418727_418727 ; 
   reg __418727_418727;
   reg _418728_418728 ; 
   reg __418728_418728;
   reg _418729_418729 ; 
   reg __418729_418729;
   reg _418730_418730 ; 
   reg __418730_418730;
   reg _418731_418731 ; 
   reg __418731_418731;
   reg _418732_418732 ; 
   reg __418732_418732;
   reg _418733_418733 ; 
   reg __418733_418733;
   reg _418734_418734 ; 
   reg __418734_418734;
   reg _418735_418735 ; 
   reg __418735_418735;
   reg _418736_418736 ; 
   reg __418736_418736;
   reg _418737_418737 ; 
   reg __418737_418737;
   reg _418738_418738 ; 
   reg __418738_418738;
   reg _418739_418739 ; 
   reg __418739_418739;
   reg _418740_418740 ; 
   reg __418740_418740;
   reg _418741_418741 ; 
   reg __418741_418741;
   reg _418742_418742 ; 
   reg __418742_418742;
   reg _418743_418743 ; 
   reg __418743_418743;
   reg _418744_418744 ; 
   reg __418744_418744;
   reg _418745_418745 ; 
   reg __418745_418745;
   reg _418746_418746 ; 
   reg __418746_418746;
   reg _418747_418747 ; 
   reg __418747_418747;
   reg _418748_418748 ; 
   reg __418748_418748;
   reg _418749_418749 ; 
   reg __418749_418749;
   reg _418750_418750 ; 
   reg __418750_418750;
   reg _418751_418751 ; 
   reg __418751_418751;
   reg _418752_418752 ; 
   reg __418752_418752;
   reg _418753_418753 ; 
   reg __418753_418753;
   reg _418754_418754 ; 
   reg __418754_418754;
   reg _418755_418755 ; 
   reg __418755_418755;
   reg _418756_418756 ; 
   reg __418756_418756;
   reg _418757_418757 ; 
   reg __418757_418757;
   reg _418758_418758 ; 
   reg __418758_418758;
   reg _418759_418759 ; 
   reg __418759_418759;
   reg _418760_418760 ; 
   reg __418760_418760;
   reg _418761_418761 ; 
   reg __418761_418761;
   reg _418762_418762 ; 
   reg __418762_418762;
   reg _418763_418763 ; 
   reg __418763_418763;
   reg _418764_418764 ; 
   reg __418764_418764;
   reg _418765_418765 ; 
   reg __418765_418765;
   reg _418766_418766 ; 
   reg __418766_418766;
   reg _418767_418767 ; 
   reg __418767_418767;
   reg _418768_418768 ; 
   reg __418768_418768;
   reg _418769_418769 ; 
   reg __418769_418769;
   reg _418770_418770 ; 
   reg __418770_418770;
   reg _418771_418771 ; 
   reg __418771_418771;
   reg _418772_418772 ; 
   reg __418772_418772;
   reg _418773_418773 ; 
   reg __418773_418773;
   reg _418774_418774 ; 
   reg __418774_418774;
   reg _418775_418775 ; 
   reg __418775_418775;
   reg _418776_418776 ; 
   reg __418776_418776;
   reg _418777_418777 ; 
   reg __418777_418777;
   reg _418778_418778 ; 
   reg __418778_418778;
   reg _418779_418779 ; 
   reg __418779_418779;
   reg _418780_418780 ; 
   reg __418780_418780;
   reg _418781_418781 ; 
   reg __418781_418781;
   reg _418782_418782 ; 
   reg __418782_418782;
   reg _418783_418783 ; 
   reg __418783_418783;
   reg _418784_418784 ; 
   reg __418784_418784;
   reg _418785_418785 ; 
   reg __418785_418785;
   reg _418786_418786 ; 
   reg __418786_418786;
   reg _418787_418787 ; 
   reg __418787_418787;
   reg _418788_418788 ; 
   reg __418788_418788;
   reg _418789_418789 ; 
   reg __418789_418789;
   reg _418790_418790 ; 
   reg __418790_418790;
   reg _418791_418791 ; 
   reg __418791_418791;
   reg _418792_418792 ; 
   reg __418792_418792;
   reg _418793_418793 ; 
   reg __418793_418793;
   reg _418794_418794 ; 
   reg __418794_418794;
   reg _418795_418795 ; 
   reg __418795_418795;
   reg _418796_418796 ; 
   reg __418796_418796;
   reg _418797_418797 ; 
   reg __418797_418797;
   reg _418798_418798 ; 
   reg __418798_418798;
   reg _418799_418799 ; 
   reg __418799_418799;
   reg _418800_418800 ; 
   reg __418800_418800;
   reg _418801_418801 ; 
   reg __418801_418801;
   reg _418802_418802 ; 
   reg __418802_418802;
   reg _418803_418803 ; 
   reg __418803_418803;
   reg _418804_418804 ; 
   reg __418804_418804;
   reg _418805_418805 ; 
   reg __418805_418805;
   reg _418806_418806 ; 
   reg __418806_418806;
   reg _418807_418807 ; 
   reg __418807_418807;
   reg _418808_418808 ; 
   reg __418808_418808;
   reg _418809_418809 ; 
   reg __418809_418809;
   reg _418810_418810 ; 
   reg __418810_418810;
   reg _418811_418811 ; 
   reg __418811_418811;
   reg _418812_418812 ; 
   reg __418812_418812;
   reg _418813_418813 ; 
   reg __418813_418813;
   reg _418814_418814 ; 
   reg __418814_418814;
   reg _418815_418815 ; 
   reg __418815_418815;
   reg _418816_418816 ; 
   reg __418816_418816;
   reg _418817_418817 ; 
   reg __418817_418817;
   reg _418818_418818 ; 
   reg __418818_418818;
   reg _418819_418819 ; 
   reg __418819_418819;
   reg _418820_418820 ; 
   reg __418820_418820;
   reg _418821_418821 ; 
   reg __418821_418821;
   reg _418822_418822 ; 
   reg __418822_418822;
   reg _418823_418823 ; 
   reg __418823_418823;
   reg _418824_418824 ; 
   reg __418824_418824;
   reg _418825_418825 ; 
   reg __418825_418825;
   reg _418826_418826 ; 
   reg __418826_418826;
   reg _418827_418827 ; 
   reg __418827_418827;
   reg _418828_418828 ; 
   reg __418828_418828;
   reg _418829_418829 ; 
   reg __418829_418829;
   reg _418830_418830 ; 
   reg __418830_418830;
   reg _418831_418831 ; 
   reg __418831_418831;
   reg _418832_418832 ; 
   reg __418832_418832;
   reg _418833_418833 ; 
   reg __418833_418833;
   reg _418834_418834 ; 
   reg __418834_418834;
   reg _418835_418835 ; 
   reg __418835_418835;
   reg _418836_418836 ; 
   reg __418836_418836;
   reg _418837_418837 ; 
   reg __418837_418837;
   reg _418838_418838 ; 
   reg __418838_418838;
   reg _418839_418839 ; 
   reg __418839_418839;
   reg _418840_418840 ; 
   reg __418840_418840;
   reg _418841_418841 ; 
   reg __418841_418841;
   reg _418842_418842 ; 
   reg __418842_418842;
   reg _418843_418843 ; 
   reg __418843_418843;
   reg _418844_418844 ; 
   reg __418844_418844;
   reg _418845_418845 ; 
   reg __418845_418845;
   reg _418846_418846 ; 
   reg __418846_418846;
   reg _418847_418847 ; 
   reg __418847_418847;
   reg _418848_418848 ; 
   reg __418848_418848;
   reg _418849_418849 ; 
   reg __418849_418849;
   reg _418850_418850 ; 
   reg __418850_418850;
   reg _418851_418851 ; 
   reg __418851_418851;
   reg _418852_418852 ; 
   reg __418852_418852;
   reg _418853_418853 ; 
   reg __418853_418853;
   reg _418854_418854 ; 
   reg __418854_418854;
   reg _418855_418855 ; 
   reg __418855_418855;
   reg _418856_418856 ; 
   reg __418856_418856;
   reg _418857_418857 ; 
   reg __418857_418857;
   reg _418858_418858 ; 
   reg __418858_418858;
   reg _418859_418859 ; 
   reg __418859_418859;
   reg _418860_418860 ; 
   reg __418860_418860;
   reg _418861_418861 ; 
   reg __418861_418861;
   reg _418862_418862 ; 
   reg __418862_418862;
   reg _418863_418863 ; 
   reg __418863_418863;
   reg _418864_418864 ; 
   reg __418864_418864;
   reg _418865_418865 ; 
   reg __418865_418865;
   reg _418866_418866 ; 
   reg __418866_418866;
   reg _418867_418867 ; 
   reg __418867_418867;
   reg _418868_418868 ; 
   reg __418868_418868;
   reg _418869_418869 ; 
   reg __418869_418869;
   reg _418870_418870 ; 
   reg __418870_418870;
   reg _418871_418871 ; 
   reg __418871_418871;
   reg _418872_418872 ; 
   reg __418872_418872;
   reg _418873_418873 ; 
   reg __418873_418873;
   reg _418874_418874 ; 
   reg __418874_418874;
   reg _418875_418875 ; 
   reg __418875_418875;
   reg _418876_418876 ; 
   reg __418876_418876;
   reg _418877_418877 ; 
   reg __418877_418877;
   reg _418878_418878 ; 
   reg __418878_418878;
   reg _418879_418879 ; 
   reg __418879_418879;
   reg _418880_418880 ; 
   reg __418880_418880;
   reg _418881_418881 ; 
   reg __418881_418881;
   reg _418882_418882 ; 
   reg __418882_418882;
   reg _418883_418883 ; 
   reg __418883_418883;
   reg _418884_418884 ; 
   reg __418884_418884;
   reg _418885_418885 ; 
   reg __418885_418885;
   reg _418886_418886 ; 
   reg __418886_418886;
   reg _418887_418887 ; 
   reg __418887_418887;
   reg _418888_418888 ; 
   reg __418888_418888;
   reg _418889_418889 ; 
   reg __418889_418889;
   reg _418890_418890 ; 
   reg __418890_418890;
   reg _418891_418891 ; 
   reg __418891_418891;
   reg _418892_418892 ; 
   reg __418892_418892;
   reg _418893_418893 ; 
   reg __418893_418893;
   reg _418894_418894 ; 
   reg __418894_418894;
   reg _418895_418895 ; 
   reg __418895_418895;
   reg _418896_418896 ; 
   reg __418896_418896;
   reg _418897_418897 ; 
   reg __418897_418897;
   reg _418898_418898 ; 
   reg __418898_418898;
   reg _418899_418899 ; 
   reg __418899_418899;
   reg _418900_418900 ; 
   reg __418900_418900;
   reg _418901_418901 ; 
   reg __418901_418901;
   reg _418902_418902 ; 
   reg __418902_418902;
   reg _418903_418903 ; 
   reg __418903_418903;
   reg _418904_418904 ; 
   reg __418904_418904;
   reg _418905_418905 ; 
   reg __418905_418905;
   reg _418906_418906 ; 
   reg __418906_418906;
   reg _418907_418907 ; 
   reg __418907_418907;
   reg _418908_418908 ; 
   reg __418908_418908;
   reg _418909_418909 ; 
   reg __418909_418909;
   reg _418910_418910 ; 
   reg __418910_418910;
   reg _418911_418911 ; 
   reg __418911_418911;
   reg _418912_418912 ; 
   reg __418912_418912;
   reg _418913_418913 ; 
   reg __418913_418913;
   reg _418914_418914 ; 
   reg __418914_418914;
   reg _418915_418915 ; 
   reg __418915_418915;
   reg _418916_418916 ; 
   reg __418916_418916;
   reg _418917_418917 ; 
   reg __418917_418917;
   reg _418918_418918 ; 
   reg __418918_418918;
   reg _418919_418919 ; 
   reg __418919_418919;
   reg _418920_418920 ; 
   reg __418920_418920;
   reg _418921_418921 ; 
   reg __418921_418921;
   reg _418922_418922 ; 
   reg __418922_418922;
   reg _418923_418923 ; 
   reg __418923_418923;
   reg _418924_418924 ; 
   reg __418924_418924;
   reg _418925_418925 ; 
   reg __418925_418925;
   reg _418926_418926 ; 
   reg __418926_418926;
   reg _418927_418927 ; 
   reg __418927_418927;
   reg _418928_418928 ; 
   reg __418928_418928;
   reg _418929_418929 ; 
   reg __418929_418929;
   reg _418930_418930 ; 
   reg __418930_418930;
   reg _418931_418931 ; 
   reg __418931_418931;
   reg _418932_418932 ; 
   reg __418932_418932;
   reg _418933_418933 ; 
   reg __418933_418933;
   reg _418934_418934 ; 
   reg __418934_418934;
   reg _418935_418935 ; 
   reg __418935_418935;
   reg _418936_418936 ; 
   reg __418936_418936;
   reg _418937_418937 ; 
   reg __418937_418937;
   reg _418938_418938 ; 
   reg __418938_418938;
   reg _418939_418939 ; 
   reg __418939_418939;
   reg _418940_418940 ; 
   reg __418940_418940;
   reg _418941_418941 ; 
   reg __418941_418941;
   reg _418942_418942 ; 
   reg __418942_418942;
   reg _418943_418943 ; 
   reg __418943_418943;
   reg _418944_418944 ; 
   reg __418944_418944;
   reg _418945_418945 ; 
   reg __418945_418945;
   reg _418946_418946 ; 
   reg __418946_418946;
   reg _418947_418947 ; 
   reg __418947_418947;
   reg _418948_418948 ; 
   reg __418948_418948;
   reg _418949_418949 ; 
   reg __418949_418949;
   reg _418950_418950 ; 
   reg __418950_418950;
   reg _418951_418951 ; 
   reg __418951_418951;
   reg _418952_418952 ; 
   reg __418952_418952;
   reg _418953_418953 ; 
   reg __418953_418953;
   reg _418954_418954 ; 
   reg __418954_418954;
   reg _418955_418955 ; 
   reg __418955_418955;
   reg _418956_418956 ; 
   reg __418956_418956;
   reg _418957_418957 ; 
   reg __418957_418957;
   reg _418958_418958 ; 
   reg __418958_418958;
   reg _418959_418959 ; 
   reg __418959_418959;
   reg _418960_418960 ; 
   reg __418960_418960;
   reg _418961_418961 ; 
   reg __418961_418961;
   reg _418962_418962 ; 
   reg __418962_418962;
   reg _418963_418963 ; 
   reg __418963_418963;
   reg _418964_418964 ; 
   reg __418964_418964;
   reg _418965_418965 ; 
   reg __418965_418965;
   reg _418966_418966 ; 
   reg __418966_418966;
   reg _418967_418967 ; 
   reg __418967_418967;
   reg _418968_418968 ; 
   reg __418968_418968;
   reg _418969_418969 ; 
   reg __418969_418969;
   reg _418970_418970 ; 
   reg __418970_418970;
   reg _418971_418971 ; 
   reg __418971_418971;
   reg _418972_418972 ; 
   reg __418972_418972;
   reg _418973_418973 ; 
   reg __418973_418973;
   reg _418974_418974 ; 
   reg __418974_418974;
   reg _418975_418975 ; 
   reg __418975_418975;
   reg _418976_418976 ; 
   reg __418976_418976;
   reg _418977_418977 ; 
   reg __418977_418977;
   reg _418978_418978 ; 
   reg __418978_418978;
   reg _418979_418979 ; 
   reg __418979_418979;
   reg _418980_418980 ; 
   reg __418980_418980;
   reg _418981_418981 ; 
   reg __418981_418981;
   reg _418982_418982 ; 
   reg __418982_418982;
   reg _418983_418983 ; 
   reg __418983_418983;
   reg _418984_418984 ; 
   reg __418984_418984;
   reg _418985_418985 ; 
   reg __418985_418985;
   reg _418986_418986 ; 
   reg __418986_418986;
   reg _418987_418987 ; 
   reg __418987_418987;
   reg _418988_418988 ; 
   reg __418988_418988;
   reg _418989_418989 ; 
   reg __418989_418989;
   reg _418990_418990 ; 
   reg __418990_418990;
   reg _418991_418991 ; 
   reg __418991_418991;
   reg _418992_418992 ; 
   reg __418992_418992;
   reg _418993_418993 ; 
   reg __418993_418993;
   reg _418994_418994 ; 
   reg __418994_418994;
   reg _418995_418995 ; 
   reg __418995_418995;
   reg _418996_418996 ; 
   reg __418996_418996;
   reg _418997_418997 ; 
   reg __418997_418997;
   reg _418998_418998 ; 
   reg __418998_418998;
   reg _418999_418999 ; 
   reg __418999_418999;
   reg _419000_419000 ; 
   reg __419000_419000;
   reg _419001_419001 ; 
   reg __419001_419001;
   reg _419002_419002 ; 
   reg __419002_419002;
   reg _419003_419003 ; 
   reg __419003_419003;
   reg _419004_419004 ; 
   reg __419004_419004;
   reg _419005_419005 ; 
   reg __419005_419005;
   reg _419006_419006 ; 
   reg __419006_419006;
   reg _419007_419007 ; 
   reg __419007_419007;
   reg _419008_419008 ; 
   reg __419008_419008;
   reg _419009_419009 ; 
   reg __419009_419009;
   reg _419010_419010 ; 
   reg __419010_419010;
   reg _419011_419011 ; 
   reg __419011_419011;
   reg _419012_419012 ; 
   reg __419012_419012;
   reg _419013_419013 ; 
   reg __419013_419013;
   reg _419014_419014 ; 
   reg __419014_419014;
   reg _419015_419015 ; 
   reg __419015_419015;
   reg _419016_419016 ; 
   reg __419016_419016;
   reg _419017_419017 ; 
   reg __419017_419017;
   reg _419018_419018 ; 
   reg __419018_419018;
   reg _419019_419019 ; 
   reg __419019_419019;
   reg _419020_419020 ; 
   reg __419020_419020;
   reg _419021_419021 ; 
   reg __419021_419021;
   reg _419022_419022 ; 
   reg __419022_419022;
   reg _419023_419023 ; 
   reg __419023_419023;
   reg _419024_419024 ; 
   reg __419024_419024;
   reg _419025_419025 ; 
   reg __419025_419025;
   reg _419026_419026 ; 
   reg __419026_419026;
   reg _419027_419027 ; 
   reg __419027_419027;
   reg _419028_419028 ; 
   reg __419028_419028;
   reg _419029_419029 ; 
   reg __419029_419029;
   reg _419030_419030 ; 
   reg __419030_419030;
   reg _419031_419031 ; 
   reg __419031_419031;
   reg _419032_419032 ; 
   reg __419032_419032;
   reg _419033_419033 ; 
   reg __419033_419033;
   reg _419034_419034 ; 
   reg __419034_419034;
   reg _419035_419035 ; 
   reg __419035_419035;
   reg _419036_419036 ; 
   reg __419036_419036;
   reg _419037_419037 ; 
   reg __419037_419037;
   reg _419038_419038 ; 
   reg __419038_419038;
   reg _419039_419039 ; 
   reg __419039_419039;
   reg _419040_419040 ; 
   reg __419040_419040;
   reg _419041_419041 ; 
   reg __419041_419041;
   reg _419042_419042 ; 
   reg __419042_419042;
   reg _419043_419043 ; 
   reg __419043_419043;
   reg _419044_419044 ; 
   reg __419044_419044;
   reg _419045_419045 ; 
   reg __419045_419045;
   reg _419046_419046 ; 
   reg __419046_419046;
   reg _419047_419047 ; 
   reg __419047_419047;
   reg _419048_419048 ; 
   reg __419048_419048;
   reg _419049_419049 ; 
   reg __419049_419049;
   reg _419050_419050 ; 
   reg __419050_419050;
   reg _419051_419051 ; 
   reg __419051_419051;
   reg _419052_419052 ; 
   reg __419052_419052;
   reg _419053_419053 ; 
   reg __419053_419053;
   reg _419054_419054 ; 
   reg __419054_419054;
   reg _419055_419055 ; 
   reg __419055_419055;
   reg _419056_419056 ; 
   reg __419056_419056;
   reg _419057_419057 ; 
   reg __419057_419057;
   reg _419058_419058 ; 
   reg __419058_419058;
   reg _419059_419059 ; 
   reg __419059_419059;
   reg _419060_419060 ; 
   reg __419060_419060;
   reg _419061_419061 ; 
   reg __419061_419061;
   reg _419062_419062 ; 
   reg __419062_419062;
   reg _419063_419063 ; 
   reg __419063_419063;
   reg _419064_419064 ; 
   reg __419064_419064;
   reg _419065_419065 ; 
   reg __419065_419065;
   reg _419066_419066 ; 
   reg __419066_419066;
   reg _419067_419067 ; 
   reg __419067_419067;
   reg _419068_419068 ; 
   reg __419068_419068;
   reg _419069_419069 ; 
   reg __419069_419069;
   reg _419070_419070 ; 
   reg __419070_419070;
   reg _419071_419071 ; 
   reg __419071_419071;
   reg _419072_419072 ; 
   reg __419072_419072;
   reg _419073_419073 ; 
   reg __419073_419073;
   reg _419074_419074 ; 
   reg __419074_419074;
   reg _419075_419075 ; 
   reg __419075_419075;
   reg _419076_419076 ; 
   reg __419076_419076;
   reg _419077_419077 ; 
   reg __419077_419077;
   reg _419078_419078 ; 
   reg __419078_419078;
   reg _419079_419079 ; 
   reg __419079_419079;
   reg _419080_419080 ; 
   reg __419080_419080;
   reg _419081_419081 ; 
   reg __419081_419081;
   reg _419082_419082 ; 
   reg __419082_419082;
   reg _419083_419083 ; 
   reg __419083_419083;
   reg _419084_419084 ; 
   reg __419084_419084;
   reg _419085_419085 ; 
   reg __419085_419085;
   reg _419086_419086 ; 
   reg __419086_419086;
   reg _419087_419087 ; 
   reg __419087_419087;
   reg _419088_419088 ; 
   reg __419088_419088;
   reg _419089_419089 ; 
   reg __419089_419089;
   reg _419090_419090 ; 
   reg __419090_419090;
   reg _419091_419091 ; 
   reg __419091_419091;
   reg _419092_419092 ; 
   reg __419092_419092;
   reg _419093_419093 ; 
   reg __419093_419093;
   reg _419094_419094 ; 
   reg __419094_419094;
   reg _419095_419095 ; 
   reg __419095_419095;
   reg _419096_419096 ; 
   reg __419096_419096;
   reg _419097_419097 ; 
   reg __419097_419097;
   reg _419098_419098 ; 
   reg __419098_419098;
   reg _419099_419099 ; 
   reg __419099_419099;
   reg _419100_419100 ; 
   reg __419100_419100;
   reg _419101_419101 ; 
   reg __419101_419101;
   reg _419102_419102 ; 
   reg __419102_419102;
   reg _419103_419103 ; 
   reg __419103_419103;
   reg _419104_419104 ; 
   reg __419104_419104;
   reg _419105_419105 ; 
   reg __419105_419105;
   reg _419106_419106 ; 
   reg __419106_419106;
   reg _419107_419107 ; 
   reg __419107_419107;
   reg _419108_419108 ; 
   reg __419108_419108;
   reg _419109_419109 ; 
   reg __419109_419109;
   reg _419110_419110 ; 
   reg __419110_419110;
   reg _419111_419111 ; 
   reg __419111_419111;
   reg _419112_419112 ; 
   reg __419112_419112;
   reg _419113_419113 ; 
   reg __419113_419113;
   reg _419114_419114 ; 
   reg __419114_419114;
   reg _419115_419115 ; 
   reg __419115_419115;
   reg _419116_419116 ; 
   reg __419116_419116;
   reg _419117_419117 ; 
   reg __419117_419117;
   reg _419118_419118 ; 
   reg __419118_419118;
   reg _419119_419119 ; 
   reg __419119_419119;
   reg _419120_419120 ; 
   reg __419120_419120;
   reg _419121_419121 ; 
   reg __419121_419121;
   reg _419122_419122 ; 
   reg __419122_419122;
   reg _419123_419123 ; 
   reg __419123_419123;
   reg _419124_419124 ; 
   reg __419124_419124;
   reg _419125_419125 ; 
   reg __419125_419125;
   reg _419126_419126 ; 
   reg __419126_419126;
   reg _419127_419127 ; 
   reg __419127_419127;
   reg _419128_419128 ; 
   reg __419128_419128;
   reg _419129_419129 ; 
   reg __419129_419129;
   reg _419130_419130 ; 
   reg __419130_419130;
   reg _419131_419131 ; 
   reg __419131_419131;
   reg _419132_419132 ; 
   reg __419132_419132;
   reg _419133_419133 ; 
   reg __419133_419133;
   reg _419134_419134 ; 
   reg __419134_419134;
   reg _419135_419135 ; 
   reg __419135_419135;
   reg _419136_419136 ; 
   reg __419136_419136;
   reg _419137_419137 ; 
   reg __419137_419137;
   reg _419138_419138 ; 
   reg __419138_419138;
   reg _419139_419139 ; 
   reg __419139_419139;
   reg _419140_419140 ; 
   reg __419140_419140;
   reg _419141_419141 ; 
   reg __419141_419141;
   reg _419142_419142 ; 
   reg __419142_419142;
   reg _419143_419143 ; 
   reg __419143_419143;
   reg _419144_419144 ; 
   reg __419144_419144;
   reg _419145_419145 ; 
   reg __419145_419145;
   reg _419146_419146 ; 
   reg __419146_419146;
   reg _419147_419147 ; 
   reg __419147_419147;
   reg _419148_419148 ; 
   reg __419148_419148;
   reg _419149_419149 ; 
   reg __419149_419149;
   reg _419150_419150 ; 
   reg __419150_419150;
   reg _419151_419151 ; 
   reg __419151_419151;
   reg _419152_419152 ; 
   reg __419152_419152;
   reg _419153_419153 ; 
   reg __419153_419153;
   reg _419154_419154 ; 
   reg __419154_419154;
   reg _419155_419155 ; 
   reg __419155_419155;
   reg _419156_419156 ; 
   reg __419156_419156;
   reg _419157_419157 ; 
   reg __419157_419157;
   reg _419158_419158 ; 
   reg __419158_419158;
   reg _419159_419159 ; 
   reg __419159_419159;
   reg _419160_419160 ; 
   reg __419160_419160;
   reg _419161_419161 ; 
   reg __419161_419161;
   reg _419162_419162 ; 
   reg __419162_419162;
   reg _419163_419163 ; 
   reg __419163_419163;
   reg _419164_419164 ; 
   reg __419164_419164;
   reg _419165_419165 ; 
   reg __419165_419165;
   reg _419166_419166 ; 
   reg __419166_419166;
   reg _419167_419167 ; 
   reg __419167_419167;
   reg _419168_419168 ; 
   reg __419168_419168;
   reg _419169_419169 ; 
   reg __419169_419169;
   reg _419170_419170 ; 
   reg __419170_419170;
   reg _419171_419171 ; 
   reg __419171_419171;
   reg _419172_419172 ; 
   reg __419172_419172;
   reg _419173_419173 ; 
   reg __419173_419173;
   reg _419174_419174 ; 
   reg __419174_419174;
   reg _419175_419175 ; 
   reg __419175_419175;
   reg _419176_419176 ; 
   reg __419176_419176;
   reg _419177_419177 ; 
   reg __419177_419177;
   reg _419178_419178 ; 
   reg __419178_419178;
   reg _419179_419179 ; 
   reg __419179_419179;
   reg _419180_419180 ; 
   reg __419180_419180;
   reg _419181_419181 ; 
   reg __419181_419181;
   reg _419182_419182 ; 
   reg __419182_419182;
   reg _419183_419183 ; 
   reg __419183_419183;
   reg _419184_419184 ; 
   reg __419184_419184;
   reg _419185_419185 ; 
   reg __419185_419185;
   reg _419186_419186 ; 
   reg __419186_419186;
   reg _419187_419187 ; 
   reg __419187_419187;
   reg _419188_419188 ; 
   reg __419188_419188;
   reg _419189_419189 ; 
   reg __419189_419189;
   reg _419190_419190 ; 
   reg __419190_419190;
   reg _419191_419191 ; 
   reg __419191_419191;
   reg _419192_419192 ; 
   reg __419192_419192;
   reg _419193_419193 ; 
   reg __419193_419193;
   reg _419194_419194 ; 
   reg __419194_419194;
   reg _419195_419195 ; 
   reg __419195_419195;
   reg _419196_419196 ; 
   reg __419196_419196;
   reg _419197_419197 ; 
   reg __419197_419197;
   reg _419198_419198 ; 
   reg __419198_419198;
   reg _419199_419199 ; 
   reg __419199_419199;
   reg _419200_419200 ; 
   reg __419200_419200;
   reg _419201_419201 ; 
   reg __419201_419201;
   reg _419202_419202 ; 
   reg __419202_419202;
   reg _419203_419203 ; 
   reg __419203_419203;
   reg _419204_419204 ; 
   reg __419204_419204;
   reg _419205_419205 ; 
   reg __419205_419205;
   reg _419206_419206 ; 
   reg __419206_419206;
   reg _419207_419207 ; 
   reg __419207_419207;
   reg _419208_419208 ; 
   reg __419208_419208;
   reg _419209_419209 ; 
   reg __419209_419209;
   reg _419210_419210 ; 
   reg __419210_419210;
   reg _419211_419211 ; 
   reg __419211_419211;
   reg _419212_419212 ; 
   reg __419212_419212;
   reg _419213_419213 ; 
   reg __419213_419213;
   reg _419214_419214 ; 
   reg __419214_419214;
   reg _419215_419215 ; 
   reg __419215_419215;
   reg _419216_419216 ; 
   reg __419216_419216;
   reg _419217_419217 ; 
   reg __419217_419217;
   reg _419218_419218 ; 
   reg __419218_419218;
   reg _419219_419219 ; 
   reg __419219_419219;
   reg _419220_419220 ; 
   reg __419220_419220;
   reg _419221_419221 ; 
   reg __419221_419221;
   reg _419222_419222 ; 
   reg __419222_419222;
   reg _419223_419223 ; 
   reg __419223_419223;
   reg _419224_419224 ; 
   reg __419224_419224;
   reg _419225_419225 ; 
   reg __419225_419225;
   reg _419226_419226 ; 
   reg __419226_419226;
   reg _419227_419227 ; 
   reg __419227_419227;
   reg _419228_419228 ; 
   reg __419228_419228;
   reg _419229_419229 ; 
   reg __419229_419229;
   reg _419230_419230 ; 
   reg __419230_419230;
   reg _419231_419231 ; 
   reg __419231_419231;
   reg _419232_419232 ; 
   reg __419232_419232;
   reg _419233_419233 ; 
   reg __419233_419233;
   reg _419234_419234 ; 
   reg __419234_419234;
   reg _419235_419235 ; 
   reg __419235_419235;
   reg _419236_419236 ; 
   reg __419236_419236;
   reg _419237_419237 ; 
   reg __419237_419237;
   reg _419238_419238 ; 
   reg __419238_419238;
   reg _419239_419239 ; 
   reg __419239_419239;
   reg _419240_419240 ; 
   reg __419240_419240;
   reg _419241_419241 ; 
   reg __419241_419241;
   reg _419242_419242 ; 
   reg __419242_419242;
   reg _419243_419243 ; 
   reg __419243_419243;
   reg _419244_419244 ; 
   reg __419244_419244;
   reg _419245_419245 ; 
   reg __419245_419245;
   reg _419246_419246 ; 
   reg __419246_419246;
   reg _419247_419247 ; 
   reg __419247_419247;
   reg _419248_419248 ; 
   reg __419248_419248;
   reg _419249_419249 ; 
   reg __419249_419249;
   reg _419250_419250 ; 
   reg __419250_419250;
   reg _419251_419251 ; 
   reg __419251_419251;
   reg _419252_419252 ; 
   reg __419252_419252;
   reg _419253_419253 ; 
   reg __419253_419253;
   reg _419254_419254 ; 
   reg __419254_419254;
   reg _419255_419255 ; 
   reg __419255_419255;
   reg _419256_419256 ; 
   reg __419256_419256;
   reg _419257_419257 ; 
   reg __419257_419257;
   reg _419258_419258 ; 
   reg __419258_419258;
   reg _419259_419259 ; 
   reg __419259_419259;
   reg _419260_419260 ; 
   reg __419260_419260;
   reg _419261_419261 ; 
   reg __419261_419261;
   reg _419262_419262 ; 
   reg __419262_419262;
   reg _419263_419263 ; 
   reg __419263_419263;
   reg _419264_419264 ; 
   reg __419264_419264;
   reg _419265_419265 ; 
   reg __419265_419265;
   reg _419266_419266 ; 
   reg __419266_419266;
   reg _419267_419267 ; 
   reg __419267_419267;
   reg _419268_419268 ; 
   reg __419268_419268;
   reg _419269_419269 ; 
   reg __419269_419269;
   reg _419270_419270 ; 
   reg __419270_419270;
   reg _419271_419271 ; 
   reg __419271_419271;
   reg _419272_419272 ; 
   reg __419272_419272;
   reg _419273_419273 ; 
   reg __419273_419273;
   reg _419274_419274 ; 
   reg __419274_419274;
   reg _419275_419275 ; 
   reg __419275_419275;
   reg _419276_419276 ; 
   reg __419276_419276;
   reg _419277_419277 ; 
   reg __419277_419277;
   reg _419278_419278 ; 
   reg __419278_419278;
   reg _419279_419279 ; 
   reg __419279_419279;
   reg _419280_419280 ; 
   reg __419280_419280;
   reg _419281_419281 ; 
   reg __419281_419281;
   reg _419282_419282 ; 
   reg __419282_419282;
   reg _419283_419283 ; 
   reg __419283_419283;
   reg _419284_419284 ; 
   reg __419284_419284;
   reg _419285_419285 ; 
   reg __419285_419285;
   reg _419286_419286 ; 
   reg __419286_419286;
   reg _419287_419287 ; 
   reg __419287_419287;
   reg _419288_419288 ; 
   reg __419288_419288;
   reg _419289_419289 ; 
   reg __419289_419289;
   reg _419290_419290 ; 
   reg __419290_419290;
   reg _419291_419291 ; 
   reg __419291_419291;
   reg _419292_419292 ; 
   reg __419292_419292;
   reg _419293_419293 ; 
   reg __419293_419293;
   reg _419294_419294 ; 
   reg __419294_419294;
   reg _419295_419295 ; 
   reg __419295_419295;
   reg _419296_419296 ; 
   reg __419296_419296;
   reg _419297_419297 ; 
   reg __419297_419297;
   reg _419298_419298 ; 
   reg __419298_419298;
   reg _419299_419299 ; 
   reg __419299_419299;
   reg _419300_419300 ; 
   reg __419300_419300;
   reg _419301_419301 ; 
   reg __419301_419301;
   reg _419302_419302 ; 
   reg __419302_419302;
   reg _419303_419303 ; 
   reg __419303_419303;
   reg _419304_419304 ; 
   reg __419304_419304;
   reg _419305_419305 ; 
   reg __419305_419305;
   reg _419306_419306 ; 
   reg __419306_419306;
   reg _419307_419307 ; 
   reg __419307_419307;
   reg _419308_419308 ; 
   reg __419308_419308;
   reg _419309_419309 ; 
   reg __419309_419309;
   reg _419310_419310 ; 
   reg __419310_419310;
   reg _419311_419311 ; 
   reg __419311_419311;
   reg _419312_419312 ; 
   reg __419312_419312;
   reg _419313_419313 ; 
   reg __419313_419313;
   reg _419314_419314 ; 
   reg __419314_419314;
   reg _419315_419315 ; 
   reg __419315_419315;
   reg _419316_419316 ; 
   reg __419316_419316;
   reg _419317_419317 ; 
   reg __419317_419317;
   reg _419318_419318 ; 
   reg __419318_419318;
   reg _419319_419319 ; 
   reg __419319_419319;
   reg _419320_419320 ; 
   reg __419320_419320;
   reg _419321_419321 ; 
   reg __419321_419321;
   reg _419322_419322 ; 
   reg __419322_419322;
   reg _419323_419323 ; 
   reg __419323_419323;
   reg _419324_419324 ; 
   reg __419324_419324;
   reg _419325_419325 ; 
   reg __419325_419325;
   reg _419326_419326 ; 
   reg __419326_419326;
   reg _419327_419327 ; 
   reg __419327_419327;
   reg _419328_419328 ; 
   reg __419328_419328;
   reg _419329_419329 ; 
   reg __419329_419329;
   reg _419330_419330 ; 
   reg __419330_419330;
   reg _419331_419331 ; 
   reg __419331_419331;
   reg _419332_419332 ; 
   reg __419332_419332;
   reg _419333_419333 ; 
   reg __419333_419333;
   reg _419334_419334 ; 
   reg __419334_419334;
   reg _419335_419335 ; 
   reg __419335_419335;
   reg _419336_419336 ; 
   reg __419336_419336;
   reg _419337_419337 ; 
   reg __419337_419337;
   reg _419338_419338 ; 
   reg __419338_419338;
   reg _419339_419339 ; 
   reg __419339_419339;
   reg _419340_419340 ; 
   reg __419340_419340;
   reg _419341_419341 ; 
   reg __419341_419341;
   reg _419342_419342 ; 
   reg __419342_419342;
   reg _419343_419343 ; 
   reg __419343_419343;
   reg _419344_419344 ; 
   reg __419344_419344;
   reg _419345_419345 ; 
   reg __419345_419345;
   reg _419346_419346 ; 
   reg __419346_419346;
   reg _419347_419347 ; 
   reg __419347_419347;
   reg _419348_419348 ; 
   reg __419348_419348;
   reg _419349_419349 ; 
   reg __419349_419349;
   reg _419350_419350 ; 
   reg __419350_419350;
   reg _419351_419351 ; 
   reg __419351_419351;
   reg _419352_419352 ; 
   reg __419352_419352;
   reg _419353_419353 ; 
   reg __419353_419353;
   reg _419354_419354 ; 
   reg __419354_419354;
   reg _419355_419355 ; 
   reg __419355_419355;
   reg _419356_419356 ; 
   reg __419356_419356;
   reg _419357_419357 ; 
   reg __419357_419357;
   reg _419358_419358 ; 
   reg __419358_419358;
   reg _419359_419359 ; 
   reg __419359_419359;
   reg _419360_419360 ; 
   reg __419360_419360;
   reg _419361_419361 ; 
   reg __419361_419361;
   reg _419362_419362 ; 
   reg __419362_419362;
   reg _419363_419363 ; 
   reg __419363_419363;
   reg _419364_419364 ; 
   reg __419364_419364;
   reg _419365_419365 ; 
   reg __419365_419365;
   reg _419366_419366 ; 
   reg __419366_419366;
   reg _419367_419367 ; 
   reg __419367_419367;
   reg _419368_419368 ; 
   reg __419368_419368;
   reg _419369_419369 ; 
   reg __419369_419369;
   reg _419370_419370 ; 
   reg __419370_419370;
   reg _419371_419371 ; 
   reg __419371_419371;
   reg _419372_419372 ; 
   reg __419372_419372;
   reg _419373_419373 ; 
   reg __419373_419373;
   reg _419374_419374 ; 
   reg __419374_419374;
   reg _419375_419375 ; 
   reg __419375_419375;
   reg _419376_419376 ; 
   reg __419376_419376;
   reg _419377_419377 ; 
   reg __419377_419377;
   reg _419378_419378 ; 
   reg __419378_419378;
   reg _419379_419379 ; 
   reg __419379_419379;
   reg _419380_419380 ; 
   reg __419380_419380;
   reg _419381_419381 ; 
   reg __419381_419381;
   reg _419382_419382 ; 
   reg __419382_419382;
   reg _419383_419383 ; 
   reg __419383_419383;
   reg _419384_419384 ; 
   reg __419384_419384;
   reg _419385_419385 ; 
   reg __419385_419385;
   reg _419386_419386 ; 
   reg __419386_419386;
   reg _419387_419387 ; 
   reg __419387_419387;
   reg _419388_419388 ; 
   reg __419388_419388;
   reg _419389_419389 ; 
   reg __419389_419389;
   reg _419390_419390 ; 
   reg __419390_419390;
   reg _419391_419391 ; 
   reg __419391_419391;
   reg _419392_419392 ; 
   reg __419392_419392;
   reg _419393_419393 ; 
   reg __419393_419393;
   reg _419394_419394 ; 
   reg __419394_419394;
   reg _419395_419395 ; 
   reg __419395_419395;
   reg _419396_419396 ; 
   reg __419396_419396;
   reg _419397_419397 ; 
   reg __419397_419397;
   reg _419398_419398 ; 
   reg __419398_419398;
   reg _419399_419399 ; 
   reg __419399_419399;
   reg _419400_419400 ; 
   reg __419400_419400;
   reg _419401_419401 ; 
   reg __419401_419401;
   reg _419402_419402 ; 
   reg __419402_419402;
   reg _419403_419403 ; 
   reg __419403_419403;
   reg _419404_419404 ; 
   reg __419404_419404;
   reg _419405_419405 ; 
   reg __419405_419405;
   reg _419406_419406 ; 
   reg __419406_419406;
   reg _419407_419407 ; 
   reg __419407_419407;
   reg _419408_419408 ; 
   reg __419408_419408;
   reg _419409_419409 ; 
   reg __419409_419409;
   reg _419410_419410 ; 
   reg __419410_419410;
   reg _419411_419411 ; 
   reg __419411_419411;
   reg _419412_419412 ; 
   reg __419412_419412;
   reg _419413_419413 ; 
   reg __419413_419413;
   reg _419414_419414 ; 
   reg __419414_419414;
   reg _419415_419415 ; 
   reg __419415_419415;
   reg _419416_419416 ; 
   reg __419416_419416;
   reg _419417_419417 ; 
   reg __419417_419417;
   reg _419418_419418 ; 
   reg __419418_419418;
   reg _419419_419419 ; 
   reg __419419_419419;
   reg _419420_419420 ; 
   reg __419420_419420;
   reg _419421_419421 ; 
   reg __419421_419421;
   reg _419422_419422 ; 
   reg __419422_419422;
   reg _419423_419423 ; 
   reg __419423_419423;
   reg _419424_419424 ; 
   reg __419424_419424;
   reg _419425_419425 ; 
   reg __419425_419425;
   reg _419426_419426 ; 
   reg __419426_419426;
   reg _419427_419427 ; 
   reg __419427_419427;
   reg _419428_419428 ; 
   reg __419428_419428;
   reg _419429_419429 ; 
   reg __419429_419429;
   reg _419430_419430 ; 
   reg __419430_419430;
   reg _419431_419431 ; 
   reg __419431_419431;
   reg _419432_419432 ; 
   reg __419432_419432;
   reg _419433_419433 ; 
   reg __419433_419433;
   reg _419434_419434 ; 
   reg __419434_419434;
   reg _419435_419435 ; 
   reg __419435_419435;
   reg _419436_419436 ; 
   reg __419436_419436;
   reg _419437_419437 ; 
   reg __419437_419437;
   reg _419438_419438 ; 
   reg __419438_419438;
   reg _419439_419439 ; 
   reg __419439_419439;
   reg _419440_419440 ; 
   reg __419440_419440;
   reg _419441_419441 ; 
   reg __419441_419441;
   reg _419442_419442 ; 
   reg __419442_419442;
   reg _419443_419443 ; 
   reg __419443_419443;
   reg _419444_419444 ; 
   reg __419444_419444;
   reg _419445_419445 ; 
   reg __419445_419445;
   reg _419446_419446 ; 
   reg __419446_419446;
   reg _419447_419447 ; 
   reg __419447_419447;
   reg _419448_419448 ; 
   reg __419448_419448;
   reg _419449_419449 ; 
   reg __419449_419449;
   reg _419450_419450 ; 
   reg __419450_419450;
   reg _419451_419451 ; 
   reg __419451_419451;
   reg _419452_419452 ; 
   reg __419452_419452;
   reg _419453_419453 ; 
   reg __419453_419453;
   reg _419454_419454 ; 
   reg __419454_419454;
   reg _419455_419455 ; 
   reg __419455_419455;
   reg _419456_419456 ; 
   reg __419456_419456;
   reg _419457_419457 ; 
   reg __419457_419457;
   reg _419458_419458 ; 
   reg __419458_419458;
   reg _419459_419459 ; 
   reg __419459_419459;
   reg _419460_419460 ; 
   reg __419460_419460;
   reg _419461_419461 ; 
   reg __419461_419461;
   reg _419462_419462 ; 
   reg __419462_419462;
   reg _419463_419463 ; 
   reg __419463_419463;
   reg _419464_419464 ; 
   reg __419464_419464;
   reg _419465_419465 ; 
   reg __419465_419465;
   reg _419466_419466 ; 
   reg __419466_419466;
   reg _419467_419467 ; 
   reg __419467_419467;
   reg _419468_419468 ; 
   reg __419468_419468;
   reg _419469_419469 ; 
   reg __419469_419469;
   reg _419470_419470 ; 
   reg __419470_419470;
   reg _419471_419471 ; 
   reg __419471_419471;
   reg _419472_419472 ; 
   reg __419472_419472;
   reg _419473_419473 ; 
   reg __419473_419473;
   reg _419474_419474 ; 
   reg __419474_419474;
   reg _419475_419475 ; 
   reg __419475_419475;
   reg _419476_419476 ; 
   reg __419476_419476;
   reg _419477_419477 ; 
   reg __419477_419477;
   reg _419478_419478 ; 
   reg __419478_419478;
   reg _419479_419479 ; 
   reg __419479_419479;
   reg _419480_419480 ; 
   reg __419480_419480;
   reg _419481_419481 ; 
   reg __419481_419481;
   reg _419482_419482 ; 
   reg __419482_419482;
   reg _419483_419483 ; 
   reg __419483_419483;
   reg _419484_419484 ; 
   reg __419484_419484;
   reg _419485_419485 ; 
   reg __419485_419485;
   reg _419486_419486 ; 
   reg __419486_419486;
   reg _419487_419487 ; 
   reg __419487_419487;
   reg _419488_419488 ; 
   reg __419488_419488;
   reg _419489_419489 ; 
   reg __419489_419489;
   reg _419490_419490 ; 
   reg __419490_419490;
   reg _419491_419491 ; 
   reg __419491_419491;
   reg _419492_419492 ; 
   reg __419492_419492;
   reg _419493_419493 ; 
   reg __419493_419493;
   reg _419494_419494 ; 
   reg __419494_419494;
   reg _419495_419495 ; 
   reg __419495_419495;
   reg _419496_419496 ; 
   reg __419496_419496;
   reg _419497_419497 ; 
   reg __419497_419497;
   reg _419498_419498 ; 
   reg __419498_419498;
   reg _419499_419499 ; 
   reg __419499_419499;
   reg _419500_419500 ; 
   reg __419500_419500;
   reg _419501_419501 ; 
   reg __419501_419501;
   reg _419502_419502 ; 
   reg __419502_419502;
   reg _419503_419503 ; 
   reg __419503_419503;
   reg _419504_419504 ; 
   reg __419504_419504;
   reg _419505_419505 ; 
   reg __419505_419505;
   reg _419506_419506 ; 
   reg __419506_419506;
   reg _419507_419507 ; 
   reg __419507_419507;
   reg _419508_419508 ; 
   reg __419508_419508;
   reg _419509_419509 ; 
   reg __419509_419509;
   reg _419510_419510 ; 
   reg __419510_419510;
   reg _419511_419511 ; 
   reg __419511_419511;
   reg _419512_419512 ; 
   reg __419512_419512;
   reg _419513_419513 ; 
   reg __419513_419513;
   reg _419514_419514 ; 
   reg __419514_419514;
   reg _419515_419515 ; 
   reg __419515_419515;
   reg _419516_419516 ; 
   reg __419516_419516;
   reg _419517_419517 ; 
   reg __419517_419517;
   reg _419518_419518 ; 
   reg __419518_419518;
   reg _419519_419519 ; 
   reg __419519_419519;
   reg _419520_419520 ; 
   reg __419520_419520;
   reg _419521_419521 ; 
   reg __419521_419521;
   reg _419522_419522 ; 
   reg __419522_419522;
   reg _419523_419523 ; 
   reg __419523_419523;
   reg _419524_419524 ; 
   reg __419524_419524;
   reg _419525_419525 ; 
   reg __419525_419525;
   reg _419526_419526 ; 
   reg __419526_419526;
   reg _419527_419527 ; 
   reg __419527_419527;
   reg _419528_419528 ; 
   reg __419528_419528;
   reg _419529_419529 ; 
   reg __419529_419529;
   reg _419530_419530 ; 
   reg __419530_419530;
   reg _419531_419531 ; 
   reg __419531_419531;
   reg _419532_419532 ; 
   reg __419532_419532;
   reg _419533_419533 ; 
   reg __419533_419533;
   reg _419534_419534 ; 
   reg __419534_419534;
   reg _419535_419535 ; 
   reg __419535_419535;
   reg _419536_419536 ; 
   reg __419536_419536;
   reg _419537_419537 ; 
   reg __419537_419537;
   reg _419538_419538 ; 
   reg __419538_419538;
   reg _419539_419539 ; 
   reg __419539_419539;
   reg _419540_419540 ; 
   reg __419540_419540;
   reg _419541_419541 ; 
   reg __419541_419541;
   reg _419542_419542 ; 
   reg __419542_419542;
   reg _419543_419543 ; 
   reg __419543_419543;
   reg _419544_419544 ; 
   reg __419544_419544;
   reg _419545_419545 ; 
   reg __419545_419545;
   reg _419546_419546 ; 
   reg __419546_419546;
   reg _419547_419547 ; 
   reg __419547_419547;
   reg _419548_419548 ; 
   reg __419548_419548;
   reg _419549_419549 ; 
   reg __419549_419549;
   reg _419550_419550 ; 
   reg __419550_419550;
   reg _419551_419551 ; 
   reg __419551_419551;
   reg _419552_419552 ; 
   reg __419552_419552;
   reg _419553_419553 ; 
   reg __419553_419553;
   reg _419554_419554 ; 
   reg __419554_419554;
   reg _419555_419555 ; 
   reg __419555_419555;
   reg _419556_419556 ; 
   reg __419556_419556;
   reg _419557_419557 ; 
   reg __419557_419557;
   reg _419558_419558 ; 
   reg __419558_419558;
   reg _419559_419559 ; 
   reg __419559_419559;
   reg _419560_419560 ; 
   reg __419560_419560;
   reg _419561_419561 ; 
   reg __419561_419561;
   reg _419562_419562 ; 
   reg __419562_419562;
   reg _419563_419563 ; 
   reg __419563_419563;
   reg _419564_419564 ; 
   reg __419564_419564;
   reg _419565_419565 ; 
   reg __419565_419565;
   reg _419566_419566 ; 
   reg __419566_419566;
   reg _419567_419567 ; 
   reg __419567_419567;
   reg _419568_419568 ; 
   reg __419568_419568;
   reg _419569_419569 ; 
   reg __419569_419569;
   reg _419570_419570 ; 
   reg __419570_419570;
   reg _419571_419571 ; 
   reg __419571_419571;
   reg _419572_419572 ; 
   reg __419572_419572;
   reg _419573_419573 ; 
   reg __419573_419573;
   reg _419574_419574 ; 
   reg __419574_419574;
   reg _419575_419575 ; 
   reg __419575_419575;
   reg _419576_419576 ; 
   reg __419576_419576;
   reg _419577_419577 ; 
   reg __419577_419577;
   reg _419578_419578 ; 
   reg __419578_419578;
   reg _419579_419579 ; 
   reg __419579_419579;
   reg _419580_419580 ; 
   reg __419580_419580;
   reg _419581_419581 ; 
   reg __419581_419581;
   reg _419582_419582 ; 
   reg __419582_419582;
   reg _419583_419583 ; 
   reg __419583_419583;
   reg _419584_419584 ; 
   reg __419584_419584;
   reg _419585_419585 ; 
   reg __419585_419585;
   reg _419586_419586 ; 
   reg __419586_419586;
   reg _419587_419587 ; 
   reg __419587_419587;
   reg _419588_419588 ; 
   reg __419588_419588;
   reg _419589_419589 ; 
   reg __419589_419589;
   reg _419590_419590 ; 
   reg __419590_419590;
   reg _419591_419591 ; 
   reg __419591_419591;
   reg _419592_419592 ; 
   reg __419592_419592;
   reg _419593_419593 ; 
   reg __419593_419593;
   reg _419594_419594 ; 
   reg __419594_419594;
   reg _419595_419595 ; 
   reg __419595_419595;
   reg _419596_419596 ; 
   reg __419596_419596;
   reg _419597_419597 ; 
   reg __419597_419597;
   reg _419598_419598 ; 
   reg __419598_419598;
   reg _419599_419599 ; 
   reg __419599_419599;
   reg _419600_419600 ; 
   reg __419600_419600;
   reg _419601_419601 ; 
   reg __419601_419601;
   reg _419602_419602 ; 
   reg __419602_419602;
   reg _419603_419603 ; 
   reg __419603_419603;
   reg _419604_419604 ; 
   reg __419604_419604;
   reg _419605_419605 ; 
   reg __419605_419605;
   reg _419606_419606 ; 
   reg __419606_419606;
   reg _419607_419607 ; 
   reg __419607_419607;
   reg _419608_419608 ; 
   reg __419608_419608;
   reg _419609_419609 ; 
   reg __419609_419609;
   reg _419610_419610 ; 
   reg __419610_419610;
   reg _419611_419611 ; 
   reg __419611_419611;
   reg _419612_419612 ; 
   reg __419612_419612;
   reg _419613_419613 ; 
   reg __419613_419613;
   reg _419614_419614 ; 
   reg __419614_419614;
   reg _419615_419615 ; 
   reg __419615_419615;
   reg _419616_419616 ; 
   reg __419616_419616;
   reg _419617_419617 ; 
   reg __419617_419617;
   reg _419618_419618 ; 
   reg __419618_419618;
   reg _419619_419619 ; 
   reg __419619_419619;
   reg _419620_419620 ; 
   reg __419620_419620;
   reg _419621_419621 ; 
   reg __419621_419621;
   reg _419622_419622 ; 
   reg __419622_419622;
   reg _419623_419623 ; 
   reg __419623_419623;
   reg _419624_419624 ; 
   reg __419624_419624;
   reg _419625_419625 ; 
   reg __419625_419625;
   reg _419626_419626 ; 
   reg __419626_419626;
   reg _419627_419627 ; 
   reg __419627_419627;
   reg _419628_419628 ; 
   reg __419628_419628;
   reg _419629_419629 ; 
   reg __419629_419629;
   reg _419630_419630 ; 
   reg __419630_419630;
   reg _419631_419631 ; 
   reg __419631_419631;
   reg _419632_419632 ; 
   reg __419632_419632;
   reg _419633_419633 ; 
   reg __419633_419633;
   reg _419634_419634 ; 
   reg __419634_419634;
   reg _419635_419635 ; 
   reg __419635_419635;
   reg _419636_419636 ; 
   reg __419636_419636;
   reg _419637_419637 ; 
   reg __419637_419637;
   reg _419638_419638 ; 
   reg __419638_419638;
   reg _419639_419639 ; 
   reg __419639_419639;
   reg _419640_419640 ; 
   reg __419640_419640;
   reg _419641_419641 ; 
   reg __419641_419641;
   reg _419642_419642 ; 
   reg __419642_419642;
   reg _419643_419643 ; 
   reg __419643_419643;
   reg _419644_419644 ; 
   reg __419644_419644;
   reg _419645_419645 ; 
   reg __419645_419645;
   reg _419646_419646 ; 
   reg __419646_419646;
   reg _419647_419647 ; 
   reg __419647_419647;
   reg _419648_419648 ; 
   reg __419648_419648;
   reg _419649_419649 ; 
   reg __419649_419649;
   reg _419650_419650 ; 
   reg __419650_419650;
   reg _419651_419651 ; 
   reg __419651_419651;
   reg _419652_419652 ; 
   reg __419652_419652;
   reg _419653_419653 ; 
   reg __419653_419653;
   reg _419654_419654 ; 
   reg __419654_419654;
   reg _419655_419655 ; 
   reg __419655_419655;
   reg _419656_419656 ; 
   reg __419656_419656;
   reg _419657_419657 ; 
   reg __419657_419657;
   reg _419658_419658 ; 
   reg __419658_419658;
   reg _419659_419659 ; 
   reg __419659_419659;
   reg _419660_419660 ; 
   reg __419660_419660;
   reg _419661_419661 ; 
   reg __419661_419661;
   reg _419662_419662 ; 
   reg __419662_419662;
   reg _419663_419663 ; 
   reg __419663_419663;
   reg _419664_419664 ; 
   reg __419664_419664;
   reg _419665_419665 ; 
   reg __419665_419665;
   reg _419666_419666 ; 
   reg __419666_419666;
   reg _419667_419667 ; 
   reg __419667_419667;
   reg _419668_419668 ; 
   reg __419668_419668;
   reg _419669_419669 ; 
   reg __419669_419669;
   reg _419670_419670 ; 
   reg __419670_419670;
   reg _419671_419671 ; 
   reg __419671_419671;
   reg _419672_419672 ; 
   reg __419672_419672;
   reg _419673_419673 ; 
   reg __419673_419673;
   reg _419674_419674 ; 
   reg __419674_419674;
   reg _419675_419675 ; 
   reg __419675_419675;
   reg _419676_419676 ; 
   reg __419676_419676;
   reg _419677_419677 ; 
   reg __419677_419677;
   reg _419678_419678 ; 
   reg __419678_419678;
   reg _419679_419679 ; 
   reg __419679_419679;
   reg _419680_419680 ; 
   reg __419680_419680;
   reg _419681_419681 ; 
   reg __419681_419681;
   reg _419682_419682 ; 
   reg __419682_419682;
   reg _419683_419683 ; 
   reg __419683_419683;
   reg _419684_419684 ; 
   reg __419684_419684;
   reg _419685_419685 ; 
   reg __419685_419685;
   reg _419686_419686 ; 
   reg __419686_419686;
   reg _419687_419687 ; 
   reg __419687_419687;
   reg _419688_419688 ; 
   reg __419688_419688;
   reg _419689_419689 ; 
   reg __419689_419689;
   reg _419690_419690 ; 
   reg __419690_419690;
   reg _419691_419691 ; 
   reg __419691_419691;
   reg _419692_419692 ; 
   reg __419692_419692;
   reg _419693_419693 ; 
   reg __419693_419693;
   reg _419694_419694 ; 
   reg __419694_419694;
   reg _419695_419695 ; 
   reg __419695_419695;
   reg _419696_419696 ; 
   reg __419696_419696;
   reg _419697_419697 ; 
   reg __419697_419697;
   reg _419698_419698 ; 
   reg __419698_419698;
   reg _419699_419699 ; 
   reg __419699_419699;
   reg _419700_419700 ; 
   reg __419700_419700;
   reg _419701_419701 ; 
   reg __419701_419701;
   reg _419702_419702 ; 
   reg __419702_419702;
   reg _419703_419703 ; 
   reg __419703_419703;
   reg _419704_419704 ; 
   reg __419704_419704;
   reg _419705_419705 ; 
   reg __419705_419705;
   reg _419706_419706 ; 
   reg __419706_419706;
   reg _419707_419707 ; 
   reg __419707_419707;
   reg _419708_419708 ; 
   reg __419708_419708;
   reg _419709_419709 ; 
   reg __419709_419709;
   reg _419710_419710 ; 
   reg __419710_419710;
   reg _419711_419711 ; 
   reg __419711_419711;
   reg _419712_419712 ; 
   reg __419712_419712;
   reg _419713_419713 ; 
   reg __419713_419713;
   reg _419714_419714 ; 
   reg __419714_419714;
   reg _419715_419715 ; 
   reg __419715_419715;
   reg _419716_419716 ; 
   reg __419716_419716;
   reg _419717_419717 ; 
   reg __419717_419717;
   reg _419718_419718 ; 
   reg __419718_419718;
   reg _419719_419719 ; 
   reg __419719_419719;
   reg _419720_419720 ; 
   reg __419720_419720;
   reg _419721_419721 ; 
   reg __419721_419721;
   reg _419722_419722 ; 
   reg __419722_419722;
   reg _419723_419723 ; 
   reg __419723_419723;
   reg _419724_419724 ; 
   reg __419724_419724;
   reg _419725_419725 ; 
   reg __419725_419725;
   reg _419726_419726 ; 
   reg __419726_419726;
   reg _419727_419727 ; 
   reg __419727_419727;
   reg _419728_419728 ; 
   reg __419728_419728;
   reg _419729_419729 ; 
   reg __419729_419729;
   reg _419730_419730 ; 
   reg __419730_419730;
   reg _419731_419731 ; 
   reg __419731_419731;
   reg _419732_419732 ; 
   reg __419732_419732;
   reg _419733_419733 ; 
   reg __419733_419733;
   reg _419734_419734 ; 
   reg __419734_419734;
   reg _419735_419735 ; 
   reg __419735_419735;
   reg _419736_419736 ; 
   reg __419736_419736;
   reg _419737_419737 ; 
   reg __419737_419737;
   reg _419738_419738 ; 
   reg __419738_419738;
   reg _419739_419739 ; 
   reg __419739_419739;
   reg _419740_419740 ; 
   reg __419740_419740;
   reg _419741_419741 ; 
   reg __419741_419741;
   reg _419742_419742 ; 
   reg __419742_419742;
   reg _419743_419743 ; 
   reg __419743_419743;
   reg _419744_419744 ; 
   reg __419744_419744;
   reg _419745_419745 ; 
   reg __419745_419745;
   reg _419746_419746 ; 
   reg __419746_419746;
   reg _419747_419747 ; 
   reg __419747_419747;
   reg _419748_419748 ; 
   reg __419748_419748;
   reg _419749_419749 ; 
   reg __419749_419749;
   reg _419750_419750 ; 
   reg __419750_419750;
   reg _419751_419751 ; 
   reg __419751_419751;
   reg _419752_419752 ; 
   reg __419752_419752;
   reg _419753_419753 ; 
   reg __419753_419753;
   reg _419754_419754 ; 
   reg __419754_419754;
   reg _419755_419755 ; 
   reg __419755_419755;
   reg _419756_419756 ; 
   reg __419756_419756;
   reg _419757_419757 ; 
   reg __419757_419757;
   reg _419758_419758 ; 
   reg __419758_419758;
   reg _419759_419759 ; 
   reg __419759_419759;
   reg _419760_419760 ; 
   reg __419760_419760;
   reg _419761_419761 ; 
   reg __419761_419761;
   reg _419762_419762 ; 
   reg __419762_419762;
   reg _419763_419763 ; 
   reg __419763_419763;
   reg _419764_419764 ; 
   reg __419764_419764;
   reg _419765_419765 ; 
   reg __419765_419765;
   reg _419766_419766 ; 
   reg __419766_419766;
   reg _419767_419767 ; 
   reg __419767_419767;
   reg _419768_419768 ; 
   reg __419768_419768;
   reg _419769_419769 ; 
   reg __419769_419769;
   reg _419770_419770 ; 
   reg __419770_419770;
   reg _419771_419771 ; 
   reg __419771_419771;
   reg _419772_419772 ; 
   reg __419772_419772;
   reg _419773_419773 ; 
   reg __419773_419773;
   reg _419774_419774 ; 
   reg __419774_419774;
   reg _419775_419775 ; 
   reg __419775_419775;
   reg _419776_419776 ; 
   reg __419776_419776;
   reg _419777_419777 ; 
   reg __419777_419777;
   reg _419778_419778 ; 
   reg __419778_419778;
   reg _419779_419779 ; 
   reg __419779_419779;
   reg _419780_419780 ; 
   reg __419780_419780;
   reg _419781_419781 ; 
   reg __419781_419781;
   reg _419782_419782 ; 
   reg __419782_419782;
   reg _419783_419783 ; 
   reg __419783_419783;
   reg _419784_419784 ; 
   reg __419784_419784;
   reg _419785_419785 ; 
   reg __419785_419785;
   reg _419786_419786 ; 
   reg __419786_419786;
   reg _419787_419787 ; 
   reg __419787_419787;
   reg _419788_419788 ; 
   reg __419788_419788;
   reg _419789_419789 ; 
   reg __419789_419789;
   reg _419790_419790 ; 
   reg __419790_419790;
   reg _419791_419791 ; 
   reg __419791_419791;
   reg _419792_419792 ; 
   reg __419792_419792;
   reg _419793_419793 ; 
   reg __419793_419793;
   reg _419794_419794 ; 
   reg __419794_419794;
   reg _419795_419795 ; 
   reg __419795_419795;
   reg _419796_419796 ; 
   reg __419796_419796;
   reg _419797_419797 ; 
   reg __419797_419797;
   reg _419798_419798 ; 
   reg __419798_419798;
   reg _419799_419799 ; 
   reg __419799_419799;
   reg _419800_419800 ; 
   reg __419800_419800;
   reg _419801_419801 ; 
   reg __419801_419801;
   reg _419802_419802 ; 
   reg __419802_419802;
   reg _419803_419803 ; 
   reg __419803_419803;
   reg _419804_419804 ; 
   reg __419804_419804;
   reg _419805_419805 ; 
   reg __419805_419805;
   reg _419806_419806 ; 
   reg __419806_419806;
   reg _419807_419807 ; 
   reg __419807_419807;
   reg _419808_419808 ; 
   reg __419808_419808;
   reg _419809_419809 ; 
   reg __419809_419809;
   reg _419810_419810 ; 
   reg __419810_419810;
   reg _419811_419811 ; 
   reg __419811_419811;
   reg _419812_419812 ; 
   reg __419812_419812;
   reg _419813_419813 ; 
   reg __419813_419813;
   reg _419814_419814 ; 
   reg __419814_419814;
   reg _419815_419815 ; 
   reg __419815_419815;
   reg _419816_419816 ; 
   reg __419816_419816;
   reg _419817_419817 ; 
   reg __419817_419817;
   reg _419818_419818 ; 
   reg __419818_419818;
   reg _419819_419819 ; 
   reg __419819_419819;
   reg _419820_419820 ; 
   reg __419820_419820;
   reg _419821_419821 ; 
   reg __419821_419821;
   reg _419822_419822 ; 
   reg __419822_419822;
   reg _419823_419823 ; 
   reg __419823_419823;
   reg _419824_419824 ; 
   reg __419824_419824;
   reg _419825_419825 ; 
   reg __419825_419825;
   reg _419826_419826 ; 
   reg __419826_419826;
   reg _419827_419827 ; 
   reg __419827_419827;
   reg _419828_419828 ; 
   reg __419828_419828;
   reg _419829_419829 ; 
   reg __419829_419829;
   reg _419830_419830 ; 
   reg __419830_419830;
   reg _419831_419831 ; 
   reg __419831_419831;
   reg _419832_419832 ; 
   reg __419832_419832;
   reg _419833_419833 ; 
   reg __419833_419833;
   reg _419834_419834 ; 
   reg __419834_419834;
   reg _419835_419835 ; 
   reg __419835_419835;
   reg _419836_419836 ; 
   reg __419836_419836;
   reg _419837_419837 ; 
   reg __419837_419837;
   reg _419838_419838 ; 
   reg __419838_419838;
   reg _419839_419839 ; 
   reg __419839_419839;
   reg _419840_419840 ; 
   reg __419840_419840;
   reg _419841_419841 ; 
   reg __419841_419841;
   reg _419842_419842 ; 
   reg __419842_419842;
   reg _419843_419843 ; 
   reg __419843_419843;
   reg _419844_419844 ; 
   reg __419844_419844;
   reg _419845_419845 ; 
   reg __419845_419845;
   reg _419846_419846 ; 
   reg __419846_419846;
   reg _419847_419847 ; 
   reg __419847_419847;
   reg _419848_419848 ; 
   reg __419848_419848;
   reg _419849_419849 ; 
   reg __419849_419849;
   reg _419850_419850 ; 
   reg __419850_419850;
   reg _419851_419851 ; 
   reg __419851_419851;
   reg _419852_419852 ; 
   reg __419852_419852;
   reg _419853_419853 ; 
   reg __419853_419853;
   reg _419854_419854 ; 
   reg __419854_419854;
   reg _419855_419855 ; 
   reg __419855_419855;
   reg _419856_419856 ; 
   reg __419856_419856;
   reg _419857_419857 ; 
   reg __419857_419857;
   reg _419858_419858 ; 
   reg __419858_419858;
   reg _419859_419859 ; 
   reg __419859_419859;
   reg _419860_419860 ; 
   reg __419860_419860;
   reg _419861_419861 ; 
   reg __419861_419861;
   reg _419862_419862 ; 
   reg __419862_419862;
   reg _419863_419863 ; 
   reg __419863_419863;
   reg _419864_419864 ; 
   reg __419864_419864;
   reg _419865_419865 ; 
   reg __419865_419865;
   reg _419866_419866 ; 
   reg __419866_419866;
   reg _419867_419867 ; 
   reg __419867_419867;
   reg _419868_419868 ; 
   reg __419868_419868;
   reg _419869_419869 ; 
   reg __419869_419869;
   reg _419870_419870 ; 
   reg __419870_419870;
   reg _419871_419871 ; 
   reg __419871_419871;
   reg _419872_419872 ; 
   reg __419872_419872;
   reg _419873_419873 ; 
   reg __419873_419873;
   reg _419874_419874 ; 
   reg __419874_419874;
   reg _419875_419875 ; 
   reg __419875_419875;
   reg _419876_419876 ; 
   reg __419876_419876;
   reg _419877_419877 ; 
   reg __419877_419877;
   reg _419878_419878 ; 
   reg __419878_419878;
   reg _419879_419879 ; 
   reg __419879_419879;
   reg _419880_419880 ; 
   reg __419880_419880;
   reg _419881_419881 ; 
   reg __419881_419881;
   reg _419882_419882 ; 
   reg __419882_419882;
   reg _419883_419883 ; 
   reg __419883_419883;
   reg _419884_419884 ; 
   reg __419884_419884;
   reg _419885_419885 ; 
   reg __419885_419885;
   reg _419886_419886 ; 
   reg __419886_419886;
   reg _419887_419887 ; 
   reg __419887_419887;
   reg _419888_419888 ; 
   reg __419888_419888;
   reg _419889_419889 ; 
   reg __419889_419889;
   reg _419890_419890 ; 
   reg __419890_419890;
   reg _419891_419891 ; 
   reg __419891_419891;
   reg _419892_419892 ; 
   reg __419892_419892;
   reg _419893_419893 ; 
   reg __419893_419893;
   reg _419894_419894 ; 
   reg __419894_419894;
   reg _419895_419895 ; 
   reg __419895_419895;
   reg _419896_419896 ; 
   reg __419896_419896;
   reg _419897_419897 ; 
   reg __419897_419897;
   reg _419898_419898 ; 
   reg __419898_419898;
   reg _419899_419899 ; 
   reg __419899_419899;
   reg _419900_419900 ; 
   reg __419900_419900;
   reg _419901_419901 ; 
   reg __419901_419901;
   reg _419902_419902 ; 
   reg __419902_419902;
   reg _419903_419903 ; 
   reg __419903_419903;
   reg _419904_419904 ; 
   reg __419904_419904;
   reg _419905_419905 ; 
   reg __419905_419905;
   reg _419906_419906 ; 
   reg __419906_419906;
   reg _419907_419907 ; 
   reg __419907_419907;
   reg _419908_419908 ; 
   reg __419908_419908;
   reg _419909_419909 ; 
   reg __419909_419909;
   reg _419910_419910 ; 
   reg __419910_419910;
   reg _419911_419911 ; 
   reg __419911_419911;
   reg _419912_419912 ; 
   reg __419912_419912;
   reg _419913_419913 ; 
   reg __419913_419913;
   reg _419914_419914 ; 
   reg __419914_419914;
   reg _419915_419915 ; 
   reg __419915_419915;
   reg _419916_419916 ; 
   reg __419916_419916;
   reg _419917_419917 ; 
   reg __419917_419917;
   reg _419918_419918 ; 
   reg __419918_419918;
   reg _419919_419919 ; 
   reg __419919_419919;
   reg _419920_419920 ; 
   reg __419920_419920;
   reg _419921_419921 ; 
   reg __419921_419921;
   reg _419922_419922 ; 
   reg __419922_419922;
   reg _419923_419923 ; 
   reg __419923_419923;
   reg _419924_419924 ; 
   reg __419924_419924;
   reg _419925_419925 ; 
   reg __419925_419925;
   reg _419926_419926 ; 
   reg __419926_419926;
   reg _419927_419927 ; 
   reg __419927_419927;
   reg _419928_419928 ; 
   reg __419928_419928;
   reg _419929_419929 ; 
   reg __419929_419929;
   reg _419930_419930 ; 
   reg __419930_419930;
   reg _419931_419931 ; 
   reg __419931_419931;
   reg _419932_419932 ; 
   reg __419932_419932;
   reg _419933_419933 ; 
   reg __419933_419933;
   reg _419934_419934 ; 
   reg __419934_419934;
   reg _419935_419935 ; 
   reg __419935_419935;
   reg _419936_419936 ; 
   reg __419936_419936;
   reg _419937_419937 ; 
   reg __419937_419937;
   reg _419938_419938 ; 
   reg __419938_419938;
   reg _419939_419939 ; 
   reg __419939_419939;
   reg _419940_419940 ; 
   reg __419940_419940;
   reg _419941_419941 ; 
   reg __419941_419941;
   reg _419942_419942 ; 
   reg __419942_419942;
   reg _419943_419943 ; 
   reg __419943_419943;
   reg _419944_419944 ; 
   reg __419944_419944;
   reg _419945_419945 ; 
   reg __419945_419945;
   reg _419946_419946 ; 
   reg __419946_419946;
   reg _419947_419947 ; 
   reg __419947_419947;
   reg _419948_419948 ; 
   reg __419948_419948;
   reg _419949_419949 ; 
   reg __419949_419949;
   reg _419950_419950 ; 
   reg __419950_419950;
   reg _419951_419951 ; 
   reg __419951_419951;
   reg _419952_419952 ; 
   reg __419952_419952;
   reg _419953_419953 ; 
   reg __419953_419953;
   reg _419954_419954 ; 
   reg __419954_419954;
   reg _419955_419955 ; 
   reg __419955_419955;
   reg _419956_419956 ; 
   reg __419956_419956;
   reg _419957_419957 ; 
   reg __419957_419957;
   reg _419958_419958 ; 
   reg __419958_419958;
   reg _419959_419959 ; 
   reg __419959_419959;
   reg _419960_419960 ; 
   reg __419960_419960;
   reg _419961_419961 ; 
   reg __419961_419961;
   reg _419962_419962 ; 
   reg __419962_419962;
   reg _419963_419963 ; 
   reg __419963_419963;
   reg _419964_419964 ; 
   reg __419964_419964;
   reg _419965_419965 ; 
   reg __419965_419965;
   reg _419966_419966 ; 
   reg __419966_419966;
   reg _419967_419967 ; 
   reg __419967_419967;
   reg _419968_419968 ; 
   reg __419968_419968;
   reg _419969_419969 ; 
   reg __419969_419969;
   reg _419970_419970 ; 
   reg __419970_419970;
   reg _419971_419971 ; 
   reg __419971_419971;
   reg _419972_419972 ; 
   reg __419972_419972;
   reg _419973_419973 ; 
   reg __419973_419973;
   reg _419974_419974 ; 
   reg __419974_419974;
   reg _419975_419975 ; 
   reg __419975_419975;
   reg _419976_419976 ; 
   reg __419976_419976;
   reg _419977_419977 ; 
   reg __419977_419977;
   reg _419978_419978 ; 
   reg __419978_419978;
   reg _419979_419979 ; 
   reg __419979_419979;
   reg _419980_419980 ; 
   reg __419980_419980;
   reg _419981_419981 ; 
   reg __419981_419981;
   reg _419982_419982 ; 
   reg __419982_419982;
   reg _419983_419983 ; 
   reg __419983_419983;
   reg _419984_419984 ; 
   reg __419984_419984;
   reg _419985_419985 ; 
   reg __419985_419985;
   reg _419986_419986 ; 
   reg __419986_419986;
   reg _419987_419987 ; 
   reg __419987_419987;
   reg _419988_419988 ; 
   reg __419988_419988;
   reg _419989_419989 ; 
   reg __419989_419989;
   reg _419990_419990 ; 
   reg __419990_419990;
   reg _419991_419991 ; 
   reg __419991_419991;
   reg _419992_419992 ; 
   reg __419992_419992;
   reg _419993_419993 ; 
   reg __419993_419993;
   reg _419994_419994 ; 
   reg __419994_419994;
   reg _419995_419995 ; 
   reg __419995_419995;
   reg _419996_419996 ; 
   reg __419996_419996;
   reg _419997_419997 ; 
   reg __419997_419997;
   reg _419998_419998 ; 
   reg __419998_419998;
   reg _419999_419999 ; 
   reg __419999_419999;
   reg _420000_420000 ; 
   reg __420000_420000;
   reg _420001_420001 ; 
   reg __420001_420001;
   reg _420002_420002 ; 
   reg __420002_420002;
   reg _420003_420003 ; 
   reg __420003_420003;
   reg _420004_420004 ; 
   reg __420004_420004;
   reg _420005_420005 ; 
   reg __420005_420005;
   reg _420006_420006 ; 
   reg __420006_420006;
   reg _420007_420007 ; 
   reg __420007_420007;
   reg _420008_420008 ; 
   reg __420008_420008;
   reg _420009_420009 ; 
   reg __420009_420009;
   reg _420010_420010 ; 
   reg __420010_420010;
   reg _420011_420011 ; 
   reg __420011_420011;
   reg _420012_420012 ; 
   reg __420012_420012;
   reg _420013_420013 ; 
   reg __420013_420013;
   reg _420014_420014 ; 
   reg __420014_420014;
   reg _420015_420015 ; 
   reg __420015_420015;
   reg _420016_420016 ; 
   reg __420016_420016;
   reg _420017_420017 ; 
   reg __420017_420017;
   reg _420018_420018 ; 
   reg __420018_420018;
   reg _420019_420019 ; 
   reg __420019_420019;
   reg _420020_420020 ; 
   reg __420020_420020;
   reg _420021_420021 ; 
   reg __420021_420021;
   reg _420022_420022 ; 
   reg __420022_420022;
   reg _420023_420023 ; 
   reg __420023_420023;
   reg _420024_420024 ; 
   reg __420024_420024;
   reg _420025_420025 ; 
   reg __420025_420025;
   reg _420026_420026 ; 
   reg __420026_420026;
   reg _420027_420027 ; 
   reg __420027_420027;
   reg _420028_420028 ; 
   reg __420028_420028;
   reg _420029_420029 ; 
   reg __420029_420029;
   reg _420030_420030 ; 
   reg __420030_420030;
   reg _420031_420031 ; 
   reg __420031_420031;
   reg _420032_420032 ; 
   reg __420032_420032;
   reg _420033_420033 ; 
   reg __420033_420033;
   reg _420034_420034 ; 
   reg __420034_420034;
   reg _420035_420035 ; 
   reg __420035_420035;
   reg _420036_420036 ; 
   reg __420036_420036;
   reg _420037_420037 ; 
   reg __420037_420037;
   reg _420038_420038 ; 
   reg __420038_420038;
   reg _420039_420039 ; 
   reg __420039_420039;
   reg _420040_420040 ; 
   reg __420040_420040;
   reg _420041_420041 ; 
   reg __420041_420041;
   reg _420042_420042 ; 
   reg __420042_420042;
   reg _420043_420043 ; 
   reg __420043_420043;
   reg _420044_420044 ; 
   reg __420044_420044;
   reg _420045_420045 ; 
   reg __420045_420045;
   reg _420046_420046 ; 
   reg __420046_420046;
   reg _420047_420047 ; 
   reg __420047_420047;
   reg _420048_420048 ; 
   reg __420048_420048;
   reg _420049_420049 ; 
   reg __420049_420049;
   reg _420050_420050 ; 
   reg __420050_420050;
   reg _420051_420051 ; 
   reg __420051_420051;
   reg _420052_420052 ; 
   reg __420052_420052;
   reg _420053_420053 ; 
   reg __420053_420053;
   reg _420054_420054 ; 
   reg __420054_420054;
   reg _420055_420055 ; 
   reg __420055_420055;
   reg _420056_420056 ; 
   reg __420056_420056;
   reg _420057_420057 ; 
   reg __420057_420057;
   reg _420058_420058 ; 
   reg __420058_420058;
   reg _420059_420059 ; 
   reg __420059_420059;
   reg _420060_420060 ; 
   reg __420060_420060;
   reg _420061_420061 ; 
   reg __420061_420061;
   reg _420062_420062 ; 
   reg __420062_420062;
   reg _420063_420063 ; 
   reg __420063_420063;
   reg _420064_420064 ; 
   reg __420064_420064;
   reg _420065_420065 ; 
   reg __420065_420065;
   reg _420066_420066 ; 
   reg __420066_420066;
   reg _420067_420067 ; 
   reg __420067_420067;
   reg _420068_420068 ; 
   reg __420068_420068;
   reg _420069_420069 ; 
   reg __420069_420069;
   reg _420070_420070 ; 
   reg __420070_420070;
   reg _420071_420071 ; 
   reg __420071_420071;
   reg _420072_420072 ; 
   reg __420072_420072;
   reg _420073_420073 ; 
   reg __420073_420073;
   reg _420074_420074 ; 
   reg __420074_420074;
   reg _420075_420075 ; 
   reg __420075_420075;
   reg _420076_420076 ; 
   reg __420076_420076;
   reg _420077_420077 ; 
   reg __420077_420077;
   reg _420078_420078 ; 
   reg __420078_420078;
   reg _420079_420079 ; 
   reg __420079_420079;
   reg _420080_420080 ; 
   reg __420080_420080;
   reg _420081_420081 ; 
   reg __420081_420081;
   reg _420082_420082 ; 
   reg __420082_420082;
   reg _420083_420083 ; 
   reg __420083_420083;
   reg _420084_420084 ; 
   reg __420084_420084;
   reg _420085_420085 ; 
   reg __420085_420085;
   reg _420086_420086 ; 
   reg __420086_420086;
   reg _420087_420087 ; 
   reg __420087_420087;
   reg _420088_420088 ; 
   reg __420088_420088;
   reg _420089_420089 ; 
   reg __420089_420089;
   reg _420090_420090 ; 
   reg __420090_420090;
   reg _420091_420091 ; 
   reg __420091_420091;
   reg _420092_420092 ; 
   reg __420092_420092;
   reg _420093_420093 ; 
   reg __420093_420093;
   reg _420094_420094 ; 
   reg __420094_420094;
   reg _420095_420095 ; 
   reg __420095_420095;
   reg _420096_420096 ; 
   reg __420096_420096;
   reg _420097_420097 ; 
   reg __420097_420097;
   reg _420098_420098 ; 
   reg __420098_420098;
   reg _420099_420099 ; 
   reg __420099_420099;
   reg _420100_420100 ; 
   reg __420100_420100;
   reg _420101_420101 ; 
   reg __420101_420101;
   reg _420102_420102 ; 
   reg __420102_420102;
   reg _420103_420103 ; 
   reg __420103_420103;
   reg _420104_420104 ; 
   reg __420104_420104;
   reg _420105_420105 ; 
   reg __420105_420105;
   reg _420106_420106 ; 
   reg __420106_420106;
   reg _420107_420107 ; 
   reg __420107_420107;
   reg _420108_420108 ; 
   reg __420108_420108;
   reg _420109_420109 ; 
   reg __420109_420109;
   reg _420110_420110 ; 
   reg __420110_420110;
   reg _420111_420111 ; 
   reg __420111_420111;
   reg _420112_420112 ; 
   reg __420112_420112;
   reg _420113_420113 ; 
   reg __420113_420113;
   reg _420114_420114 ; 
   reg __420114_420114;
   reg _420115_420115 ; 
   reg __420115_420115;
   reg _420116_420116 ; 
   reg __420116_420116;
   reg _420117_420117 ; 
   reg __420117_420117;
   reg _420118_420118 ; 
   reg __420118_420118;
   reg _420119_420119 ; 
   reg __420119_420119;
   reg _420120_420120 ; 
   reg __420120_420120;
   reg _420121_420121 ; 
   reg __420121_420121;
   reg _420122_420122 ; 
   reg __420122_420122;
   reg _420123_420123 ; 
   reg __420123_420123;
   reg _420124_420124 ; 
   reg __420124_420124;
   reg _420125_420125 ; 
   reg __420125_420125;
   reg _420126_420126 ; 
   reg __420126_420126;
   reg _420127_420127 ; 
   reg __420127_420127;
   reg _420128_420128 ; 
   reg __420128_420128;
   reg _420129_420129 ; 
   reg __420129_420129;
   reg _420130_420130 ; 
   reg __420130_420130;
   reg _420131_420131 ; 
   reg __420131_420131;
   reg _420132_420132 ; 
   reg __420132_420132;
   reg _420133_420133 ; 
   reg __420133_420133;
   reg _420134_420134 ; 
   reg __420134_420134;
   reg _420135_420135 ; 
   reg __420135_420135;
   reg _420136_420136 ; 
   reg __420136_420136;
   reg _420137_420137 ; 
   reg __420137_420137;
   reg _420138_420138 ; 
   reg __420138_420138;
   reg _420139_420139 ; 
   reg __420139_420139;
   reg _420140_420140 ; 
   reg __420140_420140;
   reg _420141_420141 ; 
   reg __420141_420141;
   reg _420142_420142 ; 
   reg __420142_420142;
   reg _420143_420143 ; 
   reg __420143_420143;
   reg _420144_420144 ; 
   reg __420144_420144;
   reg _420145_420145 ; 
   reg __420145_420145;
   reg _420146_420146 ; 
   reg __420146_420146;
   reg _420147_420147 ; 
   reg __420147_420147;
   reg _420148_420148 ; 
   reg __420148_420148;
   reg _420149_420149 ; 
   reg __420149_420149;
   reg _420150_420150 ; 
   reg __420150_420150;
   reg _420151_420151 ; 
   reg __420151_420151;
   reg _420152_420152 ; 
   reg __420152_420152;
   reg _420153_420153 ; 
   reg __420153_420153;
   reg _420154_420154 ; 
   reg __420154_420154;
   reg _420155_420155 ; 
   reg __420155_420155;
   reg _420156_420156 ; 
   reg __420156_420156;
   reg _420157_420157 ; 
   reg __420157_420157;
   reg _420158_420158 ; 
   reg __420158_420158;
   reg _420159_420159 ; 
   reg __420159_420159;
   reg _420160_420160 ; 
   reg __420160_420160;
   reg _420161_420161 ; 
   reg __420161_420161;
   reg _420162_420162 ; 
   reg __420162_420162;
   reg _420163_420163 ; 
   reg __420163_420163;
   reg _420164_420164 ; 
   reg __420164_420164;
   reg _420165_420165 ; 
   reg __420165_420165;
   reg _420166_420166 ; 
   reg __420166_420166;
   reg _420167_420167 ; 
   reg __420167_420167;
   reg _420168_420168 ; 
   reg __420168_420168;
   reg _420169_420169 ; 
   reg __420169_420169;
   reg _420170_420170 ; 
   reg __420170_420170;
   reg _420171_420171 ; 
   reg __420171_420171;
   reg _420172_420172 ; 
   reg __420172_420172;
   reg _420173_420173 ; 
   reg __420173_420173;
   reg _420174_420174 ; 
   reg __420174_420174;
   reg _420175_420175 ; 
   reg __420175_420175;
   reg _420176_420176 ; 
   reg __420176_420176;
   reg _420177_420177 ; 
   reg __420177_420177;
   reg _420178_420178 ; 
   reg __420178_420178;
   reg _420179_420179 ; 
   reg __420179_420179;
   reg _420180_420180 ; 
   reg __420180_420180;
   reg _420181_420181 ; 
   reg __420181_420181;
   reg _420182_420182 ; 
   reg __420182_420182;
   reg _420183_420183 ; 
   reg __420183_420183;
   reg _420184_420184 ; 
   reg __420184_420184;
   reg _420185_420185 ; 
   reg __420185_420185;
   reg _420186_420186 ; 
   reg __420186_420186;
   reg _420187_420187 ; 
   reg __420187_420187;
   reg _420188_420188 ; 
   reg __420188_420188;
   reg _420189_420189 ; 
   reg __420189_420189;
   reg _420190_420190 ; 
   reg __420190_420190;
   reg _420191_420191 ; 
   reg __420191_420191;
   reg _420192_420192 ; 
   reg __420192_420192;
   reg _420193_420193 ; 
   reg __420193_420193;
   reg _420194_420194 ; 
   reg __420194_420194;
   reg _420195_420195 ; 
   reg __420195_420195;
   reg _420196_420196 ; 
   reg __420196_420196;
   reg _420197_420197 ; 
   reg __420197_420197;
   reg _420198_420198 ; 
   reg __420198_420198;
   reg _420199_420199 ; 
   reg __420199_420199;
   reg _420200_420200 ; 
   reg __420200_420200;
   reg _420201_420201 ; 
   reg __420201_420201;
   reg _420202_420202 ; 
   reg __420202_420202;
   reg _420203_420203 ; 
   reg __420203_420203;
   reg _420204_420204 ; 
   reg __420204_420204;
   reg _420205_420205 ; 
   reg __420205_420205;
   reg _420206_420206 ; 
   reg __420206_420206;
   reg _420207_420207 ; 
   reg __420207_420207;
   reg _420208_420208 ; 
   reg __420208_420208;
   reg _420209_420209 ; 
   reg __420209_420209;
   reg _420210_420210 ; 
   reg __420210_420210;
   reg _420211_420211 ; 
   reg __420211_420211;
   reg _420212_420212 ; 
   reg __420212_420212;
   reg _420213_420213 ; 
   reg __420213_420213;
   reg _420214_420214 ; 
   reg __420214_420214;
   reg _420215_420215 ; 
   reg __420215_420215;
   reg _420216_420216 ; 
   reg __420216_420216;
   reg _420217_420217 ; 
   reg __420217_420217;
   reg _420218_420218 ; 
   reg __420218_420218;
   reg _420219_420219 ; 
   reg __420219_420219;
   reg _420220_420220 ; 
   reg __420220_420220;
   reg _420221_420221 ; 
   reg __420221_420221;
   reg _420222_420222 ; 
   reg __420222_420222;
   reg _420223_420223 ; 
   reg __420223_420223;
   reg _420224_420224 ; 
   reg __420224_420224;
   reg _420225_420225 ; 
   reg __420225_420225;
   reg _420226_420226 ; 
   reg __420226_420226;
   reg _420227_420227 ; 
   reg __420227_420227;
   reg _420228_420228 ; 
   reg __420228_420228;
   reg _420229_420229 ; 
   reg __420229_420229;
   reg _420230_420230 ; 
   reg __420230_420230;
   reg _420231_420231 ; 
   reg __420231_420231;
   reg _420232_420232 ; 
   reg __420232_420232;
   reg _420233_420233 ; 
   reg __420233_420233;
   reg _420234_420234 ; 
   reg __420234_420234;
   reg _420235_420235 ; 
   reg __420235_420235;
   reg _420236_420236 ; 
   reg __420236_420236;
   reg _420237_420237 ; 
   reg __420237_420237;
   reg _420238_420238 ; 
   reg __420238_420238;
   reg _420239_420239 ; 
   reg __420239_420239;
   reg _420240_420240 ; 
   reg __420240_420240;
   reg _420241_420241 ; 
   reg __420241_420241;
   reg _420242_420242 ; 
   reg __420242_420242;
   reg _420243_420243 ; 
   reg __420243_420243;
   reg _420244_420244 ; 
   reg __420244_420244;
   reg _420245_420245 ; 
   reg __420245_420245;
   reg _420246_420246 ; 
   reg __420246_420246;
   reg _420247_420247 ; 
   reg __420247_420247;
   reg _420248_420248 ; 
   reg __420248_420248;
   reg _420249_420249 ; 
   reg __420249_420249;
   reg _420250_420250 ; 
   reg __420250_420250;
   reg _420251_420251 ; 
   reg __420251_420251;
   reg _420252_420252 ; 
   reg __420252_420252;
   reg _420253_420253 ; 
   reg __420253_420253;
   reg _420254_420254 ; 
   reg __420254_420254;
   reg _420255_420255 ; 
   reg __420255_420255;
   reg _420256_420256 ; 
   reg __420256_420256;
   reg _420257_420257 ; 
   reg __420257_420257;
   reg _420258_420258 ; 
   reg __420258_420258;
   reg _420259_420259 ; 
   reg __420259_420259;
   reg _420260_420260 ; 
   reg __420260_420260;
   reg _420261_420261 ; 
   reg __420261_420261;
   reg _420262_420262 ; 
   reg __420262_420262;
   reg _420263_420263 ; 
   reg __420263_420263;
   reg _420264_420264 ; 
   reg __420264_420264;
   reg _420265_420265 ; 
   reg __420265_420265;
   reg _420266_420266 ; 
   reg __420266_420266;
   reg _420267_420267 ; 
   reg __420267_420267;
   reg _420268_420268 ; 
   reg __420268_420268;
   reg _420269_420269 ; 
   reg __420269_420269;
   reg _420270_420270 ; 
   reg __420270_420270;
   reg _420271_420271 ; 
   reg __420271_420271;
   reg _420272_420272 ; 
   reg __420272_420272;
   reg _420273_420273 ; 
   reg __420273_420273;
   reg _420274_420274 ; 
   reg __420274_420274;
   reg _420275_420275 ; 
   reg __420275_420275;
   reg _420276_420276 ; 
   reg __420276_420276;
   reg _420277_420277 ; 
   reg __420277_420277;
   reg _420278_420278 ; 
   reg __420278_420278;
   reg _420279_420279 ; 
   reg __420279_420279;
   reg _420280_420280 ; 
   reg __420280_420280;
   reg _420281_420281 ; 
   reg __420281_420281;
   reg _420282_420282 ; 
   reg __420282_420282;
   reg _420283_420283 ; 
   reg __420283_420283;
   reg _420284_420284 ; 
   reg __420284_420284;
   reg _420285_420285 ; 
   reg __420285_420285;
   reg _420286_420286 ; 
   reg __420286_420286;
   reg _420287_420287 ; 
   reg __420287_420287;
   reg _420288_420288 ; 
   reg __420288_420288;
   reg _420289_420289 ; 
   reg __420289_420289;
   reg _420290_420290 ; 
   reg __420290_420290;
   reg _420291_420291 ; 
   reg __420291_420291;
   reg _420292_420292 ; 
   reg __420292_420292;
   reg _420293_420293 ; 
   reg __420293_420293;
   reg _420294_420294 ; 
   reg __420294_420294;
   reg _420295_420295 ; 
   reg __420295_420295;
   reg _420296_420296 ; 
   reg __420296_420296;
   reg _420297_420297 ; 
   reg __420297_420297;
   reg _420298_420298 ; 
   reg __420298_420298;
   reg _420299_420299 ; 
   reg __420299_420299;
   reg _420300_420300 ; 
   reg __420300_420300;
   reg _420301_420301 ; 
   reg __420301_420301;
   reg _420302_420302 ; 
   reg __420302_420302;
   reg _420303_420303 ; 
   reg __420303_420303;
   reg _420304_420304 ; 
   reg __420304_420304;
   reg _420305_420305 ; 
   reg __420305_420305;
   reg _420306_420306 ; 
   reg __420306_420306;
   reg _420307_420307 ; 
   reg __420307_420307;
   reg _420308_420308 ; 
   reg __420308_420308;
   reg _420309_420309 ; 
   reg __420309_420309;
   reg _420310_420310 ; 
   reg __420310_420310;
   reg _420311_420311 ; 
   reg __420311_420311;
   reg _420312_420312 ; 
   reg __420312_420312;
   reg _420313_420313 ; 
   reg __420313_420313;
   reg _420314_420314 ; 
   reg __420314_420314;
   reg _420315_420315 ; 
   reg __420315_420315;
   reg _420316_420316 ; 
   reg __420316_420316;
   reg _420317_420317 ; 
   reg __420317_420317;
   reg _420318_420318 ; 
   reg __420318_420318;
   reg _420319_420319 ; 
   reg __420319_420319;
   reg _420320_420320 ; 
   reg __420320_420320;
   reg _420321_420321 ; 
   reg __420321_420321;
   reg _420322_420322 ; 
   reg __420322_420322;
   reg _420323_420323 ; 
   reg __420323_420323;
   reg _420324_420324 ; 
   reg __420324_420324;
   reg _420325_420325 ; 
   reg __420325_420325;
   reg _420326_420326 ; 
   reg __420326_420326;
   reg _420327_420327 ; 
   reg __420327_420327;
   reg _420328_420328 ; 
   reg __420328_420328;
   reg _420329_420329 ; 
   reg __420329_420329;
   reg _420330_420330 ; 
   reg __420330_420330;
   reg _420331_420331 ; 
   reg __420331_420331;
   reg _420332_420332 ; 
   reg __420332_420332;
   reg _420333_420333 ; 
   reg __420333_420333;
   reg _420334_420334 ; 
   reg __420334_420334;
   reg _420335_420335 ; 
   reg __420335_420335;
   reg _420336_420336 ; 
   reg __420336_420336;
   reg _420337_420337 ; 
   reg __420337_420337;
   reg _420338_420338 ; 
   reg __420338_420338;
   reg _420339_420339 ; 
   reg __420339_420339;
   reg _420340_420340 ; 
   reg __420340_420340;
   reg _420341_420341 ; 
   reg __420341_420341;
   reg _420342_420342 ; 
   reg __420342_420342;
   reg _420343_420343 ; 
   reg __420343_420343;
   reg _420344_420344 ; 
   reg __420344_420344;
   reg _420345_420345 ; 
   reg __420345_420345;
   reg _420346_420346 ; 
   reg __420346_420346;
   reg _420347_420347 ; 
   reg __420347_420347;
   reg _420348_420348 ; 
   reg __420348_420348;
   reg _420349_420349 ; 
   reg __420349_420349;
   reg _420350_420350 ; 
   reg __420350_420350;
   reg _420351_420351 ; 
   reg __420351_420351;
   reg _420352_420352 ; 
   reg __420352_420352;
   reg _420353_420353 ; 
   reg __420353_420353;
   reg _420354_420354 ; 
   reg __420354_420354;
   reg _420355_420355 ; 
   reg __420355_420355;
   reg _420356_420356 ; 
   reg __420356_420356;
   reg _420357_420357 ; 
   reg __420357_420357;
   reg _420358_420358 ; 
   reg __420358_420358;
   reg _420359_420359 ; 
   reg __420359_420359;
   reg _420360_420360 ; 
   reg __420360_420360;
   reg _420361_420361 ; 
   reg __420361_420361;
   reg _420362_420362 ; 
   reg __420362_420362;
   reg _420363_420363 ; 
   reg __420363_420363;
   reg _420364_420364 ; 
   reg __420364_420364;
   reg _420365_420365 ; 
   reg __420365_420365;
   reg _420366_420366 ; 
   reg __420366_420366;
   reg _420367_420367 ; 
   reg __420367_420367;
   reg _420368_420368 ; 
   reg __420368_420368;
   reg _420369_420369 ; 
   reg __420369_420369;
   reg _420370_420370 ; 
   reg __420370_420370;
   reg _420371_420371 ; 
   reg __420371_420371;
   reg _420372_420372 ; 
   reg __420372_420372;
   reg _420373_420373 ; 
   reg __420373_420373;
   reg _420374_420374 ; 
   reg __420374_420374;
   reg _420375_420375 ; 
   reg __420375_420375;
   reg _420376_420376 ; 
   reg __420376_420376;
   reg _420377_420377 ; 
   reg __420377_420377;
   reg _420378_420378 ; 
   reg __420378_420378;
   reg _420379_420379 ; 
   reg __420379_420379;
   reg _420380_420380 ; 
   reg __420380_420380;
   reg _420381_420381 ; 
   reg __420381_420381;
   reg _420382_420382 ; 
   reg __420382_420382;
   reg _420383_420383 ; 
   reg __420383_420383;
   reg _420384_420384 ; 
   reg __420384_420384;
   reg _420385_420385 ; 
   reg __420385_420385;
   reg _420386_420386 ; 
   reg __420386_420386;
   reg _420387_420387 ; 
   reg __420387_420387;
   reg _420388_420388 ; 
   reg __420388_420388;
   reg _420389_420389 ; 
   reg __420389_420389;
   reg _420390_420390 ; 
   reg __420390_420390;
   reg _420391_420391 ; 
   reg __420391_420391;
   reg _420392_420392 ; 
   reg __420392_420392;
   reg _420393_420393 ; 
   reg __420393_420393;
   reg _420394_420394 ; 
   reg __420394_420394;
   reg _420395_420395 ; 
   reg __420395_420395;
   reg _420396_420396 ; 
   reg __420396_420396;
   reg _420397_420397 ; 
   reg __420397_420397;
   reg _420398_420398 ; 
   reg __420398_420398;
   reg _420399_420399 ; 
   reg __420399_420399;
   reg _420400_420400 ; 
   reg __420400_420400;
   reg _420401_420401 ; 
   reg __420401_420401;
   reg _420402_420402 ; 
   reg __420402_420402;
   reg _420403_420403 ; 
   reg __420403_420403;
   reg _420404_420404 ; 
   reg __420404_420404;
   reg _420405_420405 ; 
   reg __420405_420405;
   reg _420406_420406 ; 
   reg __420406_420406;
   reg _420407_420407 ; 
   reg __420407_420407;
   reg _420408_420408 ; 
   reg __420408_420408;
   reg _420409_420409 ; 
   reg __420409_420409;
   reg _420410_420410 ; 
   reg __420410_420410;
   reg _420411_420411 ; 
   reg __420411_420411;
   reg _420412_420412 ; 
   reg __420412_420412;
   reg _420413_420413 ; 
   reg __420413_420413;
   reg _420414_420414 ; 
   reg __420414_420414;
   reg _420415_420415 ; 
   reg __420415_420415;
   reg _420416_420416 ; 
   reg __420416_420416;
   reg _420417_420417 ; 
   reg __420417_420417;
   reg _420418_420418 ; 
   reg __420418_420418;
   reg _420419_420419 ; 
   reg __420419_420419;
   reg _420420_420420 ; 
   reg __420420_420420;
   reg _420421_420421 ; 
   reg __420421_420421;
   reg _420422_420422 ; 
   reg __420422_420422;
   reg _420423_420423 ; 
   reg __420423_420423;
   reg _420424_420424 ; 
   reg __420424_420424;
   reg _420425_420425 ; 
   reg __420425_420425;
   reg _420426_420426 ; 
   reg __420426_420426;
   reg _420427_420427 ; 
   reg __420427_420427;
   reg _420428_420428 ; 
   reg __420428_420428;
   reg _420429_420429 ; 
   reg __420429_420429;
   reg _420430_420430 ; 
   reg __420430_420430;
   reg _420431_420431 ; 
   reg __420431_420431;
   reg _420432_420432 ; 
   reg __420432_420432;
   reg _420433_420433 ; 
   reg __420433_420433;
   reg _420434_420434 ; 
   reg __420434_420434;
   reg _420435_420435 ; 
   reg __420435_420435;
   reg _420436_420436 ; 
   reg __420436_420436;
   reg _420437_420437 ; 
   reg __420437_420437;
   reg _420438_420438 ; 
   reg __420438_420438;
   reg _420439_420439 ; 
   reg __420439_420439;
   reg _420440_420440 ; 
   reg __420440_420440;
   reg _420441_420441 ; 
   reg __420441_420441;
   reg _420442_420442 ; 
   reg __420442_420442;
   reg _420443_420443 ; 
   reg __420443_420443;
   reg _420444_420444 ; 
   reg __420444_420444;
   reg _420445_420445 ; 
   reg __420445_420445;
   reg _420446_420446 ; 
   reg __420446_420446;
   reg _420447_420447 ; 
   reg __420447_420447;
   reg _420448_420448 ; 
   reg __420448_420448;
   reg _420449_420449 ; 
   reg __420449_420449;
   reg _420450_420450 ; 
   reg __420450_420450;
   reg _420451_420451 ; 
   reg __420451_420451;
   reg _420452_420452 ; 
   reg __420452_420452;
   reg _420453_420453 ; 
   reg __420453_420453;
   reg _420454_420454 ; 
   reg __420454_420454;
   reg _420455_420455 ; 
   reg __420455_420455;
   reg _420456_420456 ; 
   reg __420456_420456;
   reg _420457_420457 ; 
   reg __420457_420457;
   reg _420458_420458 ; 
   reg __420458_420458;
   reg _420459_420459 ; 
   reg __420459_420459;
   reg _420460_420460 ; 
   reg __420460_420460;
   reg _420461_420461 ; 
   reg __420461_420461;
   reg _420462_420462 ; 
   reg __420462_420462;
   reg _420463_420463 ; 
   reg __420463_420463;
   reg _420464_420464 ; 
   reg __420464_420464;
   reg _420465_420465 ; 
   reg __420465_420465;
   reg _420466_420466 ; 
   reg __420466_420466;
   reg _420467_420467 ; 
   reg __420467_420467;
   reg _420468_420468 ; 
   reg __420468_420468;
   reg _420469_420469 ; 
   reg __420469_420469;
   reg _420470_420470 ; 
   reg __420470_420470;
   reg _420471_420471 ; 
   reg __420471_420471;
   reg _420472_420472 ; 
   reg __420472_420472;
   reg _420473_420473 ; 
   reg __420473_420473;
   reg _420474_420474 ; 
   reg __420474_420474;
   reg _420475_420475 ; 
   reg __420475_420475;
   reg _420476_420476 ; 
   reg __420476_420476;
   reg _420477_420477 ; 
   reg __420477_420477;
   reg _420478_420478 ; 
   reg __420478_420478;
   reg _420479_420479 ; 
   reg __420479_420479;
   reg _420480_420480 ; 
   reg __420480_420480;
   reg _420481_420481 ; 
   reg __420481_420481;
   reg _420482_420482 ; 
   reg __420482_420482;
   reg _420483_420483 ; 
   reg __420483_420483;
   reg _420484_420484 ; 
   reg __420484_420484;
   reg _420485_420485 ; 
   reg __420485_420485;
   reg _420486_420486 ; 
   reg __420486_420486;
   reg _420487_420487 ; 
   reg __420487_420487;
   reg _420488_420488 ; 
   reg __420488_420488;
   reg _420489_420489 ; 
   reg __420489_420489;
   reg _420490_420490 ; 
   reg __420490_420490;
   reg _420491_420491 ; 
   reg __420491_420491;
   reg _420492_420492 ; 
   reg __420492_420492;
   reg _420493_420493 ; 
   reg __420493_420493;
   reg _420494_420494 ; 
   reg __420494_420494;
   reg _420495_420495 ; 
   reg __420495_420495;
   reg _420496_420496 ; 
   reg __420496_420496;
   reg _420497_420497 ; 
   reg __420497_420497;
   reg _420498_420498 ; 
   reg __420498_420498;
   reg _420499_420499 ; 
   reg __420499_420499;
   reg _420500_420500 ; 
   reg __420500_420500;
   reg _420501_420501 ; 
   reg __420501_420501;
   reg _420502_420502 ; 
   reg __420502_420502;
   reg _420503_420503 ; 
   reg __420503_420503;
   reg _420504_420504 ; 
   reg __420504_420504;
   reg _420505_420505 ; 
   reg __420505_420505;
   reg _420506_420506 ; 
   reg __420506_420506;
   reg _420507_420507 ; 
   reg __420507_420507;
   reg _420508_420508 ; 
   reg __420508_420508;
   reg _420509_420509 ; 
   reg __420509_420509;
   reg _420510_420510 ; 
   reg __420510_420510;
   reg _420511_420511 ; 
   reg __420511_420511;
   reg _420512_420512 ; 
   reg __420512_420512;
   reg _420513_420513 ; 
   reg __420513_420513;
   reg _420514_420514 ; 
   reg __420514_420514;
   reg _420515_420515 ; 
   reg __420515_420515;
   reg _420516_420516 ; 
   reg __420516_420516;
   reg _420517_420517 ; 
   reg __420517_420517;
   reg _420518_420518 ; 
   reg __420518_420518;
   reg _420519_420519 ; 
   reg __420519_420519;
   reg _420520_420520 ; 
   reg __420520_420520;
   reg _420521_420521 ; 
   reg __420521_420521;
   reg _420522_420522 ; 
   reg __420522_420522;
   reg _420523_420523 ; 
   reg __420523_420523;
   reg _420524_420524 ; 
   reg __420524_420524;
   reg _420525_420525 ; 
   reg __420525_420525;
   reg _420526_420526 ; 
   reg __420526_420526;
   reg _420527_420527 ; 
   reg __420527_420527;
   reg _420528_420528 ; 
   reg __420528_420528;
   reg _420529_420529 ; 
   reg __420529_420529;
   reg _420530_420530 ; 
   reg __420530_420530;
   reg _420531_420531 ; 
   reg __420531_420531;
   reg _420532_420532 ; 
   reg __420532_420532;
   reg _420533_420533 ; 
   reg __420533_420533;
   reg _420534_420534 ; 
   reg __420534_420534;
   reg _420535_420535 ; 
   reg __420535_420535;
   reg _420536_420536 ; 
   reg __420536_420536;
   reg _420537_420537 ; 
   reg __420537_420537;
   reg _420538_420538 ; 
   reg __420538_420538;
   reg _420539_420539 ; 
   reg __420539_420539;
   reg _420540_420540 ; 
   reg __420540_420540;
   reg _420541_420541 ; 
   reg __420541_420541;
   reg _420542_420542 ; 
   reg __420542_420542;
   reg _420543_420543 ; 
   reg __420543_420543;
   reg _420544_420544 ; 
   reg __420544_420544;
   reg _420545_420545 ; 
   reg __420545_420545;
   reg _420546_420546 ; 
   reg __420546_420546;
   reg _420547_420547 ; 
   reg __420547_420547;
   reg _420548_420548 ; 
   reg __420548_420548;
   reg _420549_420549 ; 
   reg __420549_420549;
   reg _420550_420550 ; 
   reg __420550_420550;
   reg _420551_420551 ; 
   reg __420551_420551;
   reg _420552_420552 ; 
   reg __420552_420552;
   reg _420553_420553 ; 
   reg __420553_420553;
   reg _420554_420554 ; 
   reg __420554_420554;
   reg _420555_420555 ; 
   reg __420555_420555;
   reg _420556_420556 ; 
   reg __420556_420556;
   reg _420557_420557 ; 
   reg __420557_420557;
   reg _420558_420558 ; 
   reg __420558_420558;
   reg _420559_420559 ; 
   reg __420559_420559;
   reg _420560_420560 ; 
   reg __420560_420560;
   reg _420561_420561 ; 
   reg __420561_420561;
   reg _420562_420562 ; 
   reg __420562_420562;
   reg _420563_420563 ; 
   reg __420563_420563;
   reg _420564_420564 ; 
   reg __420564_420564;
   reg _420565_420565 ; 
   reg __420565_420565;
   reg _420566_420566 ; 
   reg __420566_420566;
   reg _420567_420567 ; 
   reg __420567_420567;
   reg _420568_420568 ; 
   reg __420568_420568;
   reg _420569_420569 ; 
   reg __420569_420569;
   reg _420570_420570 ; 
   reg __420570_420570;
   reg _420571_420571 ; 
   reg __420571_420571;
   reg _420572_420572 ; 
   reg __420572_420572;
   reg _420573_420573 ; 
   reg __420573_420573;
   reg _420574_420574 ; 
   reg __420574_420574;
   reg _420575_420575 ; 
   reg __420575_420575;
   reg _420576_420576 ; 
   reg __420576_420576;
   reg _420577_420577 ; 
   reg __420577_420577;
   reg _420578_420578 ; 
   reg __420578_420578;
   reg _420579_420579 ; 
   reg __420579_420579;
   reg _420580_420580 ; 
   reg __420580_420580;
   reg _420581_420581 ; 
   reg __420581_420581;
   reg _420582_420582 ; 
   reg __420582_420582;
   reg _420583_420583 ; 
   reg __420583_420583;
   reg _420584_420584 ; 
   reg __420584_420584;
   reg _420585_420585 ; 
   reg __420585_420585;
   reg _420586_420586 ; 
   reg __420586_420586;
   reg _420587_420587 ; 
   reg __420587_420587;
   reg _420588_420588 ; 
   reg __420588_420588;
   reg _420589_420589 ; 
   reg __420589_420589;
   reg _420590_420590 ; 
   reg __420590_420590;
   reg _420591_420591 ; 
   reg __420591_420591;
   reg _420592_420592 ; 
   reg __420592_420592;
   reg _420593_420593 ; 
   reg __420593_420593;
   reg _420594_420594 ; 
   reg __420594_420594;
   reg _420595_420595 ; 
   reg __420595_420595;
   reg _420596_420596 ; 
   reg __420596_420596;
   reg _420597_420597 ; 
   reg __420597_420597;
   reg _420598_420598 ; 
   reg __420598_420598;
   reg _420599_420599 ; 
   reg __420599_420599;
   reg _420600_420600 ; 
   reg __420600_420600;
   reg _420601_420601 ; 
   reg __420601_420601;
   reg _420602_420602 ; 
   reg __420602_420602;
   reg _420603_420603 ; 
   reg __420603_420603;
   reg _420604_420604 ; 
   reg __420604_420604;
   reg _420605_420605 ; 
   reg __420605_420605;
   reg _420606_420606 ; 
   reg __420606_420606;
   reg _420607_420607 ; 
   reg __420607_420607;
   reg _420608_420608 ; 
   reg __420608_420608;
   reg _420609_420609 ; 
   reg __420609_420609;
   reg _420610_420610 ; 
   reg __420610_420610;
   reg _420611_420611 ; 
   reg __420611_420611;
   reg _420612_420612 ; 
   reg __420612_420612;
   reg _420613_420613 ; 
   reg __420613_420613;
   reg _420614_420614 ; 
   reg __420614_420614;
   reg _420615_420615 ; 
   reg __420615_420615;
   reg _420616_420616 ; 
   reg __420616_420616;
   reg _420617_420617 ; 
   reg __420617_420617;
   reg _420618_420618 ; 
   reg __420618_420618;
   reg _420619_420619 ; 
   reg __420619_420619;
   reg _420620_420620 ; 
   reg __420620_420620;
   reg _420621_420621 ; 
   reg __420621_420621;
   reg _420622_420622 ; 
   reg __420622_420622;
   reg _420623_420623 ; 
   reg __420623_420623;
   reg _420624_420624 ; 
   reg __420624_420624;
   reg _420625_420625 ; 
   reg __420625_420625;
   reg _420626_420626 ; 
   reg __420626_420626;
   reg _420627_420627 ; 
   reg __420627_420627;
   reg _420628_420628 ; 
   reg __420628_420628;
   reg _420629_420629 ; 
   reg __420629_420629;
   reg _420630_420630 ; 
   reg __420630_420630;
   reg _420631_420631 ; 
   reg __420631_420631;
   reg _420632_420632 ; 
   reg __420632_420632;
   reg _420633_420633 ; 
   reg __420633_420633;
   reg _420634_420634 ; 
   reg __420634_420634;
   reg _420635_420635 ; 
   reg __420635_420635;
   reg _420636_420636 ; 
   reg __420636_420636;
   reg _420637_420637 ; 
   reg __420637_420637;
   reg _420638_420638 ; 
   reg __420638_420638;
   reg _420639_420639 ; 
   reg __420639_420639;
   reg _420640_420640 ; 
   reg __420640_420640;
   reg _420641_420641 ; 
   reg __420641_420641;
   reg _420642_420642 ; 
   reg __420642_420642;
   reg _420643_420643 ; 
   reg __420643_420643;
   reg _420644_420644 ; 
   reg __420644_420644;
   reg _420645_420645 ; 
   reg __420645_420645;
   reg _420646_420646 ; 
   reg __420646_420646;
   reg _420647_420647 ; 
   reg __420647_420647;
   reg _420648_420648 ; 
   reg __420648_420648;
   reg _420649_420649 ; 
   reg __420649_420649;
   reg _420650_420650 ; 
   reg __420650_420650;
   reg _420651_420651 ; 
   reg __420651_420651;
   reg _420652_420652 ; 
   reg __420652_420652;
   reg _420653_420653 ; 
   reg __420653_420653;
   reg _420654_420654 ; 
   reg __420654_420654;
   reg _420655_420655 ; 
   reg __420655_420655;
   reg _420656_420656 ; 
   reg __420656_420656;
   reg _420657_420657 ; 
   reg __420657_420657;
   reg _420658_420658 ; 
   reg __420658_420658;
   reg _420659_420659 ; 
   reg __420659_420659;
   reg _420660_420660 ; 
   reg __420660_420660;
   reg _420661_420661 ; 
   reg __420661_420661;
   reg _420662_420662 ; 
   reg __420662_420662;
   reg _420663_420663 ; 
   reg __420663_420663;
   reg _420664_420664 ; 
   reg __420664_420664;
   reg _420665_420665 ; 
   reg __420665_420665;
   reg _420666_420666 ; 
   reg __420666_420666;
   reg _420667_420667 ; 
   reg __420667_420667;
   reg _420668_420668 ; 
   reg __420668_420668;
   reg _420669_420669 ; 
   reg __420669_420669;
   reg _420670_420670 ; 
   reg __420670_420670;
   reg _420671_420671 ; 
   reg __420671_420671;
   reg _420672_420672 ; 
   reg __420672_420672;
   reg _420673_420673 ; 
   reg __420673_420673;
   reg _420674_420674 ; 
   reg __420674_420674;
   reg _420675_420675 ; 
   reg __420675_420675;
   reg _420676_420676 ; 
   reg __420676_420676;
   reg _420677_420677 ; 
   reg __420677_420677;
   reg _420678_420678 ; 
   reg __420678_420678;
   reg _420679_420679 ; 
   reg __420679_420679;
   reg _420680_420680 ; 
   reg __420680_420680;
   reg _420681_420681 ; 
   reg __420681_420681;
   reg _420682_420682 ; 
   reg __420682_420682;
   reg _420683_420683 ; 
   reg __420683_420683;
   reg _420684_420684 ; 
   reg __420684_420684;
   reg _420685_420685 ; 
   reg __420685_420685;
   reg _420686_420686 ; 
   reg __420686_420686;
   reg _420687_420687 ; 
   reg __420687_420687;
   reg _420688_420688 ; 
   reg __420688_420688;
   reg _420689_420689 ; 
   reg __420689_420689;
   reg _420690_420690 ; 
   reg __420690_420690;
   reg _420691_420691 ; 
   reg __420691_420691;
   reg _420692_420692 ; 
   reg __420692_420692;
   reg _420693_420693 ; 
   reg __420693_420693;
   reg _420694_420694 ; 
   reg __420694_420694;
   reg _420695_420695 ; 
   reg __420695_420695;
   reg _420696_420696 ; 
   reg __420696_420696;
   reg _420697_420697 ; 
   reg __420697_420697;
   reg _420698_420698 ; 
   reg __420698_420698;
   reg _420699_420699 ; 
   reg __420699_420699;
   reg _420700_420700 ; 
   reg __420700_420700;
   reg _420701_420701 ; 
   reg __420701_420701;
   reg _420702_420702 ; 
   reg __420702_420702;
   reg _420703_420703 ; 
   reg __420703_420703;
   reg _420704_420704 ; 
   reg __420704_420704;
   reg _420705_420705 ; 
   reg __420705_420705;
   reg _420706_420706 ; 
   reg __420706_420706;
   reg _420707_420707 ; 
   reg __420707_420707;
   reg _420708_420708 ; 
   reg __420708_420708;
   reg _420709_420709 ; 
   reg __420709_420709;
   reg _420710_420710 ; 
   reg __420710_420710;
   reg _420711_420711 ; 
   reg __420711_420711;
   reg _420712_420712 ; 
   reg __420712_420712;
   reg _420713_420713 ; 
   reg __420713_420713;
   reg _420714_420714 ; 
   reg __420714_420714;
   reg _420715_420715 ; 
   reg __420715_420715;
   reg _420716_420716 ; 
   reg __420716_420716;
   reg _420717_420717 ; 
   reg __420717_420717;
   reg _420718_420718 ; 
   reg __420718_420718;
   reg _420719_420719 ; 
   reg __420719_420719;
   reg _420720_420720 ; 
   reg __420720_420720;
   reg _420721_420721 ; 
   reg __420721_420721;
   reg _420722_420722 ; 
   reg __420722_420722;
   reg _420723_420723 ; 
   reg __420723_420723;
   reg _420724_420724 ; 
   reg __420724_420724;
   reg _420725_420725 ; 
   reg __420725_420725;
   reg _420726_420726 ; 
   reg __420726_420726;
   reg _420727_420727 ; 
   reg __420727_420727;
   reg _420728_420728 ; 
   reg __420728_420728;
   reg _420729_420729 ; 
   reg __420729_420729;
   reg _420730_420730 ; 
   reg __420730_420730;
   reg _420731_420731 ; 
   reg __420731_420731;
   reg _420732_420732 ; 
   reg __420732_420732;
   reg _420733_420733 ; 
   reg __420733_420733;
   reg _420734_420734 ; 
   reg __420734_420734;
   reg _420735_420735 ; 
   reg __420735_420735;
   reg _420736_420736 ; 
   reg __420736_420736;
   reg _420737_420737 ; 
   reg __420737_420737;
   reg _420738_420738 ; 
   reg __420738_420738;
   reg _420739_420739 ; 
   reg __420739_420739;
   reg _420740_420740 ; 
   reg __420740_420740;
   reg _420741_420741 ; 
   reg __420741_420741;
   reg _420742_420742 ; 
   reg __420742_420742;
   reg _420743_420743 ; 
   reg __420743_420743;
   reg _420744_420744 ; 
   reg __420744_420744;
   reg _420745_420745 ; 
   reg __420745_420745;
   reg _420746_420746 ; 
   reg __420746_420746;
   reg _420747_420747 ; 
   reg __420747_420747;
   reg _420748_420748 ; 
   reg __420748_420748;
   reg _420749_420749 ; 
   reg __420749_420749;
   reg _420750_420750 ; 
   reg __420750_420750;
   reg _420751_420751 ; 
   reg __420751_420751;
   reg _420752_420752 ; 
   reg __420752_420752;
   reg _420753_420753 ; 
   reg __420753_420753;
   reg _420754_420754 ; 
   reg __420754_420754;
   reg _420755_420755 ; 
   reg __420755_420755;
   reg _420756_420756 ; 
   reg __420756_420756;
   reg _420757_420757 ; 
   reg __420757_420757;
   reg _420758_420758 ; 
   reg __420758_420758;
   reg _420759_420759 ; 
   reg __420759_420759;
   reg _420760_420760 ; 
   reg __420760_420760;
   reg _420761_420761 ; 
   reg __420761_420761;
   reg _420762_420762 ; 
   reg __420762_420762;
   reg _420763_420763 ; 
   reg __420763_420763;
   reg _420764_420764 ; 
   reg __420764_420764;
   reg _420765_420765 ; 
   reg __420765_420765;
   reg _420766_420766 ; 
   reg __420766_420766;
   reg _420767_420767 ; 
   reg __420767_420767;
   reg _420768_420768 ; 
   reg __420768_420768;
   reg _420769_420769 ; 
   reg __420769_420769;
   reg _420770_420770 ; 
   reg __420770_420770;
   reg _420771_420771 ; 
   reg __420771_420771;
   reg _420772_420772 ; 
   reg __420772_420772;
   reg _420773_420773 ; 
   reg __420773_420773;
   reg _420774_420774 ; 
   reg __420774_420774;
   reg _420775_420775 ; 
   reg __420775_420775;
   reg _420776_420776 ; 
   reg __420776_420776;
   reg _420777_420777 ; 
   reg __420777_420777;
   reg _420778_420778 ; 
   reg __420778_420778;
   reg _420779_420779 ; 
   reg __420779_420779;
   reg _420780_420780 ; 
   reg __420780_420780;
   reg _420781_420781 ; 
   reg __420781_420781;
   reg _420782_420782 ; 
   reg __420782_420782;
   reg _420783_420783 ; 
   reg __420783_420783;
   reg _420784_420784 ; 
   reg __420784_420784;
   reg _420785_420785 ; 
   reg __420785_420785;
   reg _420786_420786 ; 
   reg __420786_420786;
   reg _420787_420787 ; 
   reg __420787_420787;
   reg _420788_420788 ; 
   reg __420788_420788;
   reg _420789_420789 ; 
   reg __420789_420789;
   reg _420790_420790 ; 
   reg __420790_420790;
   reg _420791_420791 ; 
   reg __420791_420791;
   reg _420792_420792 ; 
   reg __420792_420792;
   reg _420793_420793 ; 
   reg __420793_420793;
   reg _420794_420794 ; 
   reg __420794_420794;
   reg _420795_420795 ; 
   reg __420795_420795;
   reg _420796_420796 ; 
   reg __420796_420796;
   reg _420797_420797 ; 
   reg __420797_420797;
   reg _420798_420798 ; 
   reg __420798_420798;
   reg _420799_420799 ; 
   reg __420799_420799;
   reg _420800_420800 ; 
   reg __420800_420800;
   reg _420801_420801 ; 
   reg __420801_420801;
   reg _420802_420802 ; 
   reg __420802_420802;
   reg _420803_420803 ; 
   reg __420803_420803;
   reg _420804_420804 ; 
   reg __420804_420804;
   reg _420805_420805 ; 
   reg __420805_420805;
   reg _420806_420806 ; 
   reg __420806_420806;
   reg _420807_420807 ; 
   reg __420807_420807;
   reg _420808_420808 ; 
   reg __420808_420808;
   reg _420809_420809 ; 
   reg __420809_420809;
   reg _420810_420810 ; 
   reg __420810_420810;
   reg _420811_420811 ; 
   reg __420811_420811;
   reg _420812_420812 ; 
   reg __420812_420812;
   reg _420813_420813 ; 
   reg __420813_420813;
   reg _420814_420814 ; 
   reg __420814_420814;
   reg _420815_420815 ; 
   reg __420815_420815;
   reg _420816_420816 ; 
   reg __420816_420816;
   reg _420817_420817 ; 
   reg __420817_420817;
   reg _420818_420818 ; 
   reg __420818_420818;
   reg _420819_420819 ; 
   reg __420819_420819;
   reg _420820_420820 ; 
   reg __420820_420820;
   reg _420821_420821 ; 
   reg __420821_420821;
   reg _420822_420822 ; 
   reg __420822_420822;
   reg _420823_420823 ; 
   reg __420823_420823;
   reg _420824_420824 ; 
   reg __420824_420824;
   reg _420825_420825 ; 
   reg __420825_420825;
   reg _420826_420826 ; 
   reg __420826_420826;
   reg _420827_420827 ; 
   reg __420827_420827;
   reg _420828_420828 ; 
   reg __420828_420828;
   reg _420829_420829 ; 
   reg __420829_420829;
   reg _420830_420830 ; 
   reg __420830_420830;
   reg _420831_420831 ; 
   reg __420831_420831;
   reg _420832_420832 ; 
   reg __420832_420832;
   reg _420833_420833 ; 
   reg __420833_420833;
   reg _420834_420834 ; 
   reg __420834_420834;
   reg _420835_420835 ; 
   reg __420835_420835;
   reg _420836_420836 ; 
   reg __420836_420836;
   reg _420837_420837 ; 
   reg __420837_420837;
   reg _420838_420838 ; 
   reg __420838_420838;
   reg _420839_420839 ; 
   reg __420839_420839;
   reg _420840_420840 ; 
   reg __420840_420840;
   reg _420841_420841 ; 
   reg __420841_420841;
   reg _420842_420842 ; 
   reg __420842_420842;
   reg _420843_420843 ; 
   reg __420843_420843;
   reg _420844_420844 ; 
   reg __420844_420844;
   reg _420845_420845 ; 
   reg __420845_420845;
   reg _420846_420846 ; 
   reg __420846_420846;
   reg _420847_420847 ; 
   reg __420847_420847;
   reg _420848_420848 ; 
   reg __420848_420848;
   reg _420849_420849 ; 
   reg __420849_420849;
   reg _420850_420850 ; 
   reg __420850_420850;
   reg _420851_420851 ; 
   reg __420851_420851;
   reg _420852_420852 ; 
   reg __420852_420852;
   reg _420853_420853 ; 
   reg __420853_420853;
   reg _420854_420854 ; 
   reg __420854_420854;
   reg _420855_420855 ; 
   reg __420855_420855;
   reg _420856_420856 ; 
   reg __420856_420856;
   reg _420857_420857 ; 
   reg __420857_420857;
   reg _420858_420858 ; 
   reg __420858_420858;
   reg _420859_420859 ; 
   reg __420859_420859;
   reg _420860_420860 ; 
   reg __420860_420860;
   reg _420861_420861 ; 
   reg __420861_420861;
   reg _420862_420862 ; 
   reg __420862_420862;
   reg _420863_420863 ; 
   reg __420863_420863;
   reg _420864_420864 ; 
   reg __420864_420864;
   reg _420865_420865 ; 
   reg __420865_420865;
   reg _420866_420866 ; 
   reg __420866_420866;
   reg _420867_420867 ; 
   reg __420867_420867;
   reg _420868_420868 ; 
   reg __420868_420868;
   reg _420869_420869 ; 
   reg __420869_420869;
   reg _420870_420870 ; 
   reg __420870_420870;
   reg _420871_420871 ; 
   reg __420871_420871;
   reg _420872_420872 ; 
   reg __420872_420872;
   reg _420873_420873 ; 
   reg __420873_420873;
   reg _420874_420874 ; 
   reg __420874_420874;
   reg _420875_420875 ; 
   reg __420875_420875;
   reg _420876_420876 ; 
   reg __420876_420876;
   reg _420877_420877 ; 
   reg __420877_420877;
   reg _420878_420878 ; 
   reg __420878_420878;
   reg _420879_420879 ; 
   reg __420879_420879;
   reg _420880_420880 ; 
   reg __420880_420880;
   reg _420881_420881 ; 
   reg __420881_420881;
   reg _420882_420882 ; 
   reg __420882_420882;
   reg _420883_420883 ; 
   reg __420883_420883;
   reg _420884_420884 ; 
   reg __420884_420884;
   reg _420885_420885 ; 
   reg __420885_420885;
   reg _420886_420886 ; 
   reg __420886_420886;
   reg _420887_420887 ; 
   reg __420887_420887;
   reg _420888_420888 ; 
   reg __420888_420888;
   reg _420889_420889 ; 
   reg __420889_420889;
   reg _420890_420890 ; 
   reg __420890_420890;
   reg _420891_420891 ; 
   reg __420891_420891;
   reg _420892_420892 ; 
   reg __420892_420892;
   reg _420893_420893 ; 
   reg __420893_420893;
   reg _420894_420894 ; 
   reg __420894_420894;
   reg _420895_420895 ; 
   reg __420895_420895;
   reg _420896_420896 ; 
   reg __420896_420896;
   reg _420897_420897 ; 
   reg __420897_420897;
   reg _420898_420898 ; 
   reg __420898_420898;
   reg _420899_420899 ; 
   reg __420899_420899;
   reg _420900_420900 ; 
   reg __420900_420900;
   reg _420901_420901 ; 
   reg __420901_420901;
   reg _420902_420902 ; 
   reg __420902_420902;
   reg _420903_420903 ; 
   reg __420903_420903;
   reg _420904_420904 ; 
   reg __420904_420904;
   reg _420905_420905 ; 
   reg __420905_420905;
   reg _420906_420906 ; 
   reg __420906_420906;
   reg _420907_420907 ; 
   reg __420907_420907;
   reg _420908_420908 ; 
   reg __420908_420908;
   reg _420909_420909 ; 
   reg __420909_420909;
   reg _420910_420910 ; 
   reg __420910_420910;
   reg _420911_420911 ; 
   reg __420911_420911;
   reg _420912_420912 ; 
   reg __420912_420912;
   reg _420913_420913 ; 
   reg __420913_420913;
   reg _420914_420914 ; 
   reg __420914_420914;
   reg _420915_420915 ; 
   reg __420915_420915;
   reg _420916_420916 ; 
   reg __420916_420916;
   reg _420917_420917 ; 
   reg __420917_420917;
   reg _420918_420918 ; 
   reg __420918_420918;
   reg _420919_420919 ; 
   reg __420919_420919;
   reg _420920_420920 ; 
   reg __420920_420920;
   reg _420921_420921 ; 
   reg __420921_420921;
   reg _420922_420922 ; 
   reg __420922_420922;
   reg _420923_420923 ; 
   reg __420923_420923;
   reg _420924_420924 ; 
   reg __420924_420924;
   reg _420925_420925 ; 
   reg __420925_420925;
   reg _420926_420926 ; 
   reg __420926_420926;
   reg _420927_420927 ; 
   reg __420927_420927;
   reg _420928_420928 ; 
   reg __420928_420928;
   reg _420929_420929 ; 
   reg __420929_420929;
   reg _420930_420930 ; 
   reg __420930_420930;
   reg _420931_420931 ; 
   reg __420931_420931;
   reg _420932_420932 ; 
   reg __420932_420932;
   reg _420933_420933 ; 
   reg __420933_420933;
   reg _420934_420934 ; 
   reg __420934_420934;
   reg _420935_420935 ; 
   reg __420935_420935;
   reg _420936_420936 ; 
   reg __420936_420936;
   reg _420937_420937 ; 
   reg __420937_420937;
   reg _420938_420938 ; 
   reg __420938_420938;
   reg _420939_420939 ; 
   reg __420939_420939;
   reg _420940_420940 ; 
   reg __420940_420940;
   reg _420941_420941 ; 
   reg __420941_420941;
   reg _420942_420942 ; 
   reg __420942_420942;
   reg _420943_420943 ; 
   reg __420943_420943;
   reg _420944_420944 ; 
   reg __420944_420944;
   reg _420945_420945 ; 
   reg __420945_420945;
   reg _420946_420946 ; 
   reg __420946_420946;
   reg _420947_420947 ; 
   reg __420947_420947;
   reg _420948_420948 ; 
   reg __420948_420948;
   reg _420949_420949 ; 
   reg __420949_420949;
   reg _420950_420950 ; 
   reg __420950_420950;
   reg _420951_420951 ; 
   reg __420951_420951;
   reg _420952_420952 ; 
   reg __420952_420952;
   reg _420953_420953 ; 
   reg __420953_420953;
   reg _420954_420954 ; 
   reg __420954_420954;
   reg _420955_420955 ; 
   reg __420955_420955;
   reg _420956_420956 ; 
   reg __420956_420956;
   reg _420957_420957 ; 
   reg __420957_420957;
   reg _420958_420958 ; 
   reg __420958_420958;
   reg _420959_420959 ; 
   reg __420959_420959;
   reg _420960_420960 ; 
   reg __420960_420960;
   reg _420961_420961 ; 
   reg __420961_420961;
   reg _420962_420962 ; 
   reg __420962_420962;
   reg _420963_420963 ; 
   reg __420963_420963;
   reg _420964_420964 ; 
   reg __420964_420964;
   reg _420965_420965 ; 
   reg __420965_420965;
   reg _420966_420966 ; 
   reg __420966_420966;
   reg _420967_420967 ; 
   reg __420967_420967;
   reg _420968_420968 ; 
   reg __420968_420968;
   reg _420969_420969 ; 
   reg __420969_420969;
   reg _420970_420970 ; 
   reg __420970_420970;
   reg _420971_420971 ; 
   reg __420971_420971;
   reg _420972_420972 ; 
   reg __420972_420972;
   reg _420973_420973 ; 
   reg __420973_420973;
   reg _420974_420974 ; 
   reg __420974_420974;
   reg _420975_420975 ; 
   reg __420975_420975;
   reg _420976_420976 ; 
   reg __420976_420976;
   reg _420977_420977 ; 
   reg __420977_420977;
   reg _420978_420978 ; 
   reg __420978_420978;
   reg _420979_420979 ; 
   reg __420979_420979;
   reg _420980_420980 ; 
   reg __420980_420980;
   reg _420981_420981 ; 
   reg __420981_420981;
   reg _420982_420982 ; 
   reg __420982_420982;
   reg _420983_420983 ; 
   reg __420983_420983;
   reg _420984_420984 ; 
   reg __420984_420984;
   reg _420985_420985 ; 
   reg __420985_420985;
   reg _420986_420986 ; 
   reg __420986_420986;
   reg _420987_420987 ; 
   reg __420987_420987;
   reg _420988_420988 ; 
   reg __420988_420988;
   reg _420989_420989 ; 
   reg __420989_420989;
   reg _420990_420990 ; 
   reg __420990_420990;
   reg _420991_420991 ; 
   reg __420991_420991;
   reg _420992_420992 ; 
   reg __420992_420992;
   reg _420993_420993 ; 
   reg __420993_420993;
   reg _420994_420994 ; 
   reg __420994_420994;
   reg _420995_420995 ; 
   reg __420995_420995;
   reg _420996_420996 ; 
   reg __420996_420996;
   reg _420997_420997 ; 
   reg __420997_420997;
   reg _420998_420998 ; 
   reg __420998_420998;
   reg _420999_420999 ; 
   reg __420999_420999;
   reg _421000_421000 ; 
   reg __421000_421000;
   reg _421001_421001 ; 
   reg __421001_421001;
   reg _421002_421002 ; 
   reg __421002_421002;
   reg _421003_421003 ; 
   reg __421003_421003;
   reg _421004_421004 ; 
   reg __421004_421004;
   reg _421005_421005 ; 
   reg __421005_421005;
   reg _421006_421006 ; 
   reg __421006_421006;
   reg _421007_421007 ; 
   reg __421007_421007;
   reg _421008_421008 ; 
   reg __421008_421008;
   reg _421009_421009 ; 
   reg __421009_421009;
   reg _421010_421010 ; 
   reg __421010_421010;
   reg _421011_421011 ; 
   reg __421011_421011;
   reg _421012_421012 ; 
   reg __421012_421012;
   reg _421013_421013 ; 
   reg __421013_421013;
   reg _421014_421014 ; 
   reg __421014_421014;
   reg _421015_421015 ; 
   reg __421015_421015;
   reg _421016_421016 ; 
   reg __421016_421016;
   reg _421017_421017 ; 
   reg __421017_421017;
   reg _421018_421018 ; 
   reg __421018_421018;
   reg _421019_421019 ; 
   reg __421019_421019;
   reg _421020_421020 ; 
   reg __421020_421020;
   reg _421021_421021 ; 
   reg __421021_421021;
   reg _421022_421022 ; 
   reg __421022_421022;
   reg _421023_421023 ; 
   reg __421023_421023;
   reg _421024_421024 ; 
   reg __421024_421024;
   reg _421025_421025 ; 
   reg __421025_421025;
   reg _421026_421026 ; 
   reg __421026_421026;
   reg _421027_421027 ; 
   reg __421027_421027;
   reg _421028_421028 ; 
   reg __421028_421028;
   reg _421029_421029 ; 
   reg __421029_421029;
   reg _421030_421030 ; 
   reg __421030_421030;
   reg _421031_421031 ; 
   reg __421031_421031;
   reg _421032_421032 ; 
   reg __421032_421032;
   reg _421033_421033 ; 
   reg __421033_421033;
   reg _421034_421034 ; 
   reg __421034_421034;
   reg _421035_421035 ; 
   reg __421035_421035;
   reg _421036_421036 ; 
   reg __421036_421036;
   reg _421037_421037 ; 
   reg __421037_421037;
   reg _421038_421038 ; 
   reg __421038_421038;
   reg _421039_421039 ; 
   reg __421039_421039;
   reg _421040_421040 ; 
   reg __421040_421040;
   reg _421041_421041 ; 
   reg __421041_421041;
   reg _421042_421042 ; 
   reg __421042_421042;
   reg _421043_421043 ; 
   reg __421043_421043;
   reg _421044_421044 ; 
   reg __421044_421044;
   reg _421045_421045 ; 
   reg __421045_421045;
   reg _421046_421046 ; 
   reg __421046_421046;
   reg _421047_421047 ; 
   reg __421047_421047;
   reg _421048_421048 ; 
   reg __421048_421048;
   reg _421049_421049 ; 
   reg __421049_421049;
   reg _421050_421050 ; 
   reg __421050_421050;
   reg _421051_421051 ; 
   reg __421051_421051;
   reg _421052_421052 ; 
   reg __421052_421052;
   reg _421053_421053 ; 
   reg __421053_421053;
   reg _421054_421054 ; 
   reg __421054_421054;
   reg _421055_421055 ; 
   reg __421055_421055;
   reg _421056_421056 ; 
   reg __421056_421056;
   reg _421057_421057 ; 
   reg __421057_421057;
   reg _421058_421058 ; 
   reg __421058_421058;
   reg _421059_421059 ; 
   reg __421059_421059;
   reg _421060_421060 ; 
   reg __421060_421060;
   reg _421061_421061 ; 
   reg __421061_421061;
   reg _421062_421062 ; 
   reg __421062_421062;
   reg _421063_421063 ; 
   reg __421063_421063;
   reg _421064_421064 ; 
   reg __421064_421064;
   reg _421065_421065 ; 
   reg __421065_421065;
   reg _421066_421066 ; 
   reg __421066_421066;
   reg _421067_421067 ; 
   reg __421067_421067;
   reg _421068_421068 ; 
   reg __421068_421068;
   reg _421069_421069 ; 
   reg __421069_421069;
   reg _421070_421070 ; 
   reg __421070_421070;
   reg _421071_421071 ; 
   reg __421071_421071;
   reg _421072_421072 ; 
   reg __421072_421072;
   reg _421073_421073 ; 
   reg __421073_421073;
   reg _421074_421074 ; 
   reg __421074_421074;
   reg _421075_421075 ; 
   reg __421075_421075;
   reg _421076_421076 ; 
   reg __421076_421076;
   reg _421077_421077 ; 
   reg __421077_421077;
   reg _421078_421078 ; 
   reg __421078_421078;
   reg _421079_421079 ; 
   reg __421079_421079;
   reg _421080_421080 ; 
   reg __421080_421080;
   reg _421081_421081 ; 
   reg __421081_421081;
   reg _421082_421082 ; 
   reg __421082_421082;
   reg _421083_421083 ; 
   reg __421083_421083;
   reg _421084_421084 ; 
   reg __421084_421084;
   reg _421085_421085 ; 
   reg __421085_421085;
   reg _421086_421086 ; 
   reg __421086_421086;
   reg _421087_421087 ; 
   reg __421087_421087;
   reg _421088_421088 ; 
   reg __421088_421088;
   reg _421089_421089 ; 
   reg __421089_421089;
   reg _421090_421090 ; 
   reg __421090_421090;
   reg _421091_421091 ; 
   reg __421091_421091;
   reg _421092_421092 ; 
   reg __421092_421092;
   reg _421093_421093 ; 
   reg __421093_421093;
   reg _421094_421094 ; 
   reg __421094_421094;
   reg _421095_421095 ; 
   reg __421095_421095;
   reg _421096_421096 ; 
   reg __421096_421096;
   reg _421097_421097 ; 
   reg __421097_421097;
   reg _421098_421098 ; 
   reg __421098_421098;
   reg _421099_421099 ; 
   reg __421099_421099;
   reg _421100_421100 ; 
   reg __421100_421100;
   reg _421101_421101 ; 
   reg __421101_421101;
   reg _421102_421102 ; 
   reg __421102_421102;
   reg _421103_421103 ; 
   reg __421103_421103;
   reg _421104_421104 ; 
   reg __421104_421104;
   reg _421105_421105 ; 
   reg __421105_421105;
   reg _421106_421106 ; 
   reg __421106_421106;
   reg _421107_421107 ; 
   reg __421107_421107;
   reg _421108_421108 ; 
   reg __421108_421108;
   reg _421109_421109 ; 
   reg __421109_421109;
   reg _421110_421110 ; 
   reg __421110_421110;
   reg _421111_421111 ; 
   reg __421111_421111;
   reg _421112_421112 ; 
   reg __421112_421112;
   reg _421113_421113 ; 
   reg __421113_421113;
   reg _421114_421114 ; 
   reg __421114_421114;
   reg _421115_421115 ; 
   reg __421115_421115;
   reg _421116_421116 ; 
   reg __421116_421116;
   reg _421117_421117 ; 
   reg __421117_421117;
   reg _421118_421118 ; 
   reg __421118_421118;
   reg _421119_421119 ; 
   reg __421119_421119;
   reg _421120_421120 ; 
   reg __421120_421120;
   reg _421121_421121 ; 
   reg __421121_421121;
   reg _421122_421122 ; 
   reg __421122_421122;
   reg _421123_421123 ; 
   reg __421123_421123;
   reg _421124_421124 ; 
   reg __421124_421124;
   reg _421125_421125 ; 
   reg __421125_421125;
   reg _421126_421126 ; 
   reg __421126_421126;
   reg _421127_421127 ; 
   reg __421127_421127;
   reg _421128_421128 ; 
   reg __421128_421128;
   reg _421129_421129 ; 
   reg __421129_421129;
   reg _421130_421130 ; 
   reg __421130_421130;
   reg _421131_421131 ; 
   reg __421131_421131;
   reg _421132_421132 ; 
   reg __421132_421132;
   reg _421133_421133 ; 
   reg __421133_421133;
   reg _421134_421134 ; 
   reg __421134_421134;
   reg _421135_421135 ; 
   reg __421135_421135;
   reg _421136_421136 ; 
   reg __421136_421136;
   reg _421137_421137 ; 
   reg __421137_421137;
   reg _421138_421138 ; 
   reg __421138_421138;
   reg _421139_421139 ; 
   reg __421139_421139;
   reg _421140_421140 ; 
   reg __421140_421140;
   reg _421141_421141 ; 
   reg __421141_421141;
   reg _421142_421142 ; 
   reg __421142_421142;
   reg _421143_421143 ; 
   reg __421143_421143;
   reg _421144_421144 ; 
   reg __421144_421144;
   reg _421145_421145 ; 
   reg __421145_421145;
   reg _421146_421146 ; 
   reg __421146_421146;
   reg _421147_421147 ; 
   reg __421147_421147;
   reg _421148_421148 ; 
   reg __421148_421148;
   reg _421149_421149 ; 
   reg __421149_421149;
   reg _421150_421150 ; 
   reg __421150_421150;
   reg _421151_421151 ; 
   reg __421151_421151;
   reg _421152_421152 ; 
   reg __421152_421152;
   reg _421153_421153 ; 
   reg __421153_421153;
   reg _421154_421154 ; 
   reg __421154_421154;
   reg _421155_421155 ; 
   reg __421155_421155;
   reg _421156_421156 ; 
   reg __421156_421156;
   reg _421157_421157 ; 
   reg __421157_421157;
   reg _421158_421158 ; 
   reg __421158_421158;
   reg _421159_421159 ; 
   reg __421159_421159;
   reg _421160_421160 ; 
   reg __421160_421160;
   reg _421161_421161 ; 
   reg __421161_421161;
   reg _421162_421162 ; 
   reg __421162_421162;
   reg _421163_421163 ; 
   reg __421163_421163;
   reg _421164_421164 ; 
   reg __421164_421164;
   reg _421165_421165 ; 
   reg __421165_421165;
   reg _421166_421166 ; 
   reg __421166_421166;
   reg _421167_421167 ; 
   reg __421167_421167;
   reg _421168_421168 ; 
   reg __421168_421168;
   reg _421169_421169 ; 
   reg __421169_421169;
   reg _421170_421170 ; 
   reg __421170_421170;
   reg _421171_421171 ; 
   reg __421171_421171;
   reg _421172_421172 ; 
   reg __421172_421172;
   reg _421173_421173 ; 
   reg __421173_421173;
   reg _421174_421174 ; 
   reg __421174_421174;
   reg _421175_421175 ; 
   reg __421175_421175;
   reg _421176_421176 ; 
   reg __421176_421176;
   reg _421177_421177 ; 
   reg __421177_421177;
   reg _421178_421178 ; 
   reg __421178_421178;
   reg _421179_421179 ; 
   reg __421179_421179;
   reg _421180_421180 ; 
   reg __421180_421180;
   reg _421181_421181 ; 
   reg __421181_421181;
   reg _421182_421182 ; 
   reg __421182_421182;
   reg _421183_421183 ; 
   reg __421183_421183;
   reg _421184_421184 ; 
   reg __421184_421184;
   reg _421185_421185 ; 
   reg __421185_421185;
   reg _421186_421186 ; 
   reg __421186_421186;
   reg _421187_421187 ; 
   reg __421187_421187;
   reg _421188_421188 ; 
   reg __421188_421188;
   reg _421189_421189 ; 
   reg __421189_421189;
   reg _421190_421190 ; 
   reg __421190_421190;
   reg _421191_421191 ; 
   reg __421191_421191;
   reg _421192_421192 ; 
   reg __421192_421192;
   reg _421193_421193 ; 
   reg __421193_421193;
   reg _421194_421194 ; 
   reg __421194_421194;
   reg _421195_421195 ; 
   reg __421195_421195;
   reg _421196_421196 ; 
   reg __421196_421196;
   reg _421197_421197 ; 
   reg __421197_421197;
   reg _421198_421198 ; 
   reg __421198_421198;
   reg _421199_421199 ; 
   reg __421199_421199;
   reg _421200_421200 ; 
   reg __421200_421200;
   reg _421201_421201 ; 
   reg __421201_421201;
   reg _421202_421202 ; 
   reg __421202_421202;
   reg _421203_421203 ; 
   reg __421203_421203;
   reg _421204_421204 ; 
   reg __421204_421204;
   reg _421205_421205 ; 
   reg __421205_421205;
   reg _421206_421206 ; 
   reg __421206_421206;
   reg _421207_421207 ; 
   reg __421207_421207;
   reg _421208_421208 ; 
   reg __421208_421208;
   reg _421209_421209 ; 
   reg __421209_421209;
   reg _421210_421210 ; 
   reg __421210_421210;
   reg _421211_421211 ; 
   reg __421211_421211;
   reg _421212_421212 ; 
   reg __421212_421212;
   reg _421213_421213 ; 
   reg __421213_421213;
   reg _421214_421214 ; 
   reg __421214_421214;
   reg _421215_421215 ; 
   reg __421215_421215;
   reg _421216_421216 ; 
   reg __421216_421216;
   reg _421217_421217 ; 
   reg __421217_421217;
   reg _421218_421218 ; 
   reg __421218_421218;
   reg _421219_421219 ; 
   reg __421219_421219;
   reg _421220_421220 ; 
   reg __421220_421220;
   reg _421221_421221 ; 
   reg __421221_421221;
   reg _421222_421222 ; 
   reg __421222_421222;
   reg _421223_421223 ; 
   reg __421223_421223;
   reg _421224_421224 ; 
   reg __421224_421224;
   reg _421225_421225 ; 
   reg __421225_421225;
   reg _421226_421226 ; 
   reg __421226_421226;
   reg _421227_421227 ; 
   reg __421227_421227;
   reg _421228_421228 ; 
   reg __421228_421228;
   reg _421229_421229 ; 
   reg __421229_421229;
   reg _421230_421230 ; 
   reg __421230_421230;
   reg _421231_421231 ; 
   reg __421231_421231;
   reg _421232_421232 ; 
   reg __421232_421232;
   reg _421233_421233 ; 
   reg __421233_421233;
   reg _421234_421234 ; 
   reg __421234_421234;
   reg _421235_421235 ; 
   reg __421235_421235;
   reg _421236_421236 ; 
   reg __421236_421236;
   reg _421237_421237 ; 
   reg __421237_421237;
   reg _421238_421238 ; 
   reg __421238_421238;
   reg _421239_421239 ; 
   reg __421239_421239;
   reg _421240_421240 ; 
   reg __421240_421240;
   reg _421241_421241 ; 
   reg __421241_421241;
   reg _421242_421242 ; 
   reg __421242_421242;
   reg _421243_421243 ; 
   reg __421243_421243;
   reg _421244_421244 ; 
   reg __421244_421244;
   reg _421245_421245 ; 
   reg __421245_421245;
   reg _421246_421246 ; 
   reg __421246_421246;
   reg _421247_421247 ; 
   reg __421247_421247;
   reg _421248_421248 ; 
   reg __421248_421248;
   reg _421249_421249 ; 
   reg __421249_421249;
   reg _421250_421250 ; 
   reg __421250_421250;
   reg _421251_421251 ; 
   reg __421251_421251;
   reg _421252_421252 ; 
   reg __421252_421252;
   reg _421253_421253 ; 
   reg __421253_421253;
   reg _421254_421254 ; 
   reg __421254_421254;
   reg _421255_421255 ; 
   reg __421255_421255;
   reg _421256_421256 ; 
   reg __421256_421256;
   reg _421257_421257 ; 
   reg __421257_421257;
   reg _421258_421258 ; 
   reg __421258_421258;
   reg _421259_421259 ; 
   reg __421259_421259;
   reg _421260_421260 ; 
   reg __421260_421260;
   reg _421261_421261 ; 
   reg __421261_421261;
   reg _421262_421262 ; 
   reg __421262_421262;
   reg _421263_421263 ; 
   reg __421263_421263;
   reg _421264_421264 ; 
   reg __421264_421264;
   reg _421265_421265 ; 
   reg __421265_421265;
   reg _421266_421266 ; 
   reg __421266_421266;
   reg _421267_421267 ; 
   reg __421267_421267;
   reg _421268_421268 ; 
   reg __421268_421268;
   reg _421269_421269 ; 
   reg __421269_421269;
   reg _421270_421270 ; 
   reg __421270_421270;
   reg _421271_421271 ; 
   reg __421271_421271;
   reg _421272_421272 ; 
   reg __421272_421272;
   reg _421273_421273 ; 
   reg __421273_421273;
   reg _421274_421274 ; 
   reg __421274_421274;
   reg _421275_421275 ; 
   reg __421275_421275;
   reg _421276_421276 ; 
   reg __421276_421276;
   reg _421277_421277 ; 
   reg __421277_421277;
   reg _421278_421278 ; 
   reg __421278_421278;
   reg _421279_421279 ; 
   reg __421279_421279;
   reg _421280_421280 ; 
   reg __421280_421280;
   reg _421281_421281 ; 
   reg __421281_421281;
   reg _421282_421282 ; 
   reg __421282_421282;
   reg _421283_421283 ; 
   reg __421283_421283;
   reg _421284_421284 ; 
   reg __421284_421284;
   reg _421285_421285 ; 
   reg __421285_421285;
   reg _421286_421286 ; 
   reg __421286_421286;
   reg _421287_421287 ; 
   reg __421287_421287;
   reg _421288_421288 ; 
   reg __421288_421288;
   reg _421289_421289 ; 
   reg __421289_421289;
   reg _421290_421290 ; 
   reg __421290_421290;
   reg _421291_421291 ; 
   reg __421291_421291;
   reg _421292_421292 ; 
   reg __421292_421292;
   reg _421293_421293 ; 
   reg __421293_421293;
   reg _421294_421294 ; 
   reg __421294_421294;
   reg _421295_421295 ; 
   reg __421295_421295;
   reg _421296_421296 ; 
   reg __421296_421296;
   reg _421297_421297 ; 
   reg __421297_421297;
   reg _421298_421298 ; 
   reg __421298_421298;
   reg _421299_421299 ; 
   reg __421299_421299;
   reg _421300_421300 ; 
   reg __421300_421300;
   reg _421301_421301 ; 
   reg __421301_421301;
   reg _421302_421302 ; 
   reg __421302_421302;
   reg _421303_421303 ; 
   reg __421303_421303;
   reg _421304_421304 ; 
   reg __421304_421304;
   reg _421305_421305 ; 
   reg __421305_421305;
   reg _421306_421306 ; 
   reg __421306_421306;
   reg _421307_421307 ; 
   reg __421307_421307;
   reg _421308_421308 ; 
   reg __421308_421308;
   reg _421309_421309 ; 
   reg __421309_421309;
   reg _421310_421310 ; 
   reg __421310_421310;
   reg _421311_421311 ; 
   reg __421311_421311;
   reg _421312_421312 ; 
   reg __421312_421312;
   reg _421313_421313 ; 
   reg __421313_421313;
   reg _421314_421314 ; 
   reg __421314_421314;
   reg _421315_421315 ; 
   reg __421315_421315;
   reg _421316_421316 ; 
   reg __421316_421316;
   reg _421317_421317 ; 
   reg __421317_421317;
   reg _421318_421318 ; 
   reg __421318_421318;
   reg _421319_421319 ; 
   reg __421319_421319;
   reg _421320_421320 ; 
   reg __421320_421320;
   reg _421321_421321 ; 
   reg __421321_421321;
   reg _421322_421322 ; 
   reg __421322_421322;
   reg _421323_421323 ; 
   reg __421323_421323;
   reg _421324_421324 ; 
   reg __421324_421324;
   reg _421325_421325 ; 
   reg __421325_421325;
   reg _421326_421326 ; 
   reg __421326_421326;
   reg _421327_421327 ; 
   reg __421327_421327;
   reg _421328_421328 ; 
   reg __421328_421328;
   reg _421329_421329 ; 
   reg __421329_421329;
   reg _421330_421330 ; 
   reg __421330_421330;
   reg _421331_421331 ; 
   reg __421331_421331;
   reg _421332_421332 ; 
   reg __421332_421332;
   reg _421333_421333 ; 
   reg __421333_421333;
   reg _421334_421334 ; 
   reg __421334_421334;
   reg _421335_421335 ; 
   reg __421335_421335;
   reg _421336_421336 ; 
   reg __421336_421336;
   reg _421337_421337 ; 
   reg __421337_421337;
   reg _421338_421338 ; 
   reg __421338_421338;
   reg _421339_421339 ; 
   reg __421339_421339;
   reg _421340_421340 ; 
   reg __421340_421340;
   reg _421341_421341 ; 
   reg __421341_421341;
   reg _421342_421342 ; 
   reg __421342_421342;
   reg _421343_421343 ; 
   reg __421343_421343;
   reg _421344_421344 ; 
   reg __421344_421344;
   reg _421345_421345 ; 
   reg __421345_421345;
   reg _421346_421346 ; 
   reg __421346_421346;
   reg _421347_421347 ; 
   reg __421347_421347;
   reg _421348_421348 ; 
   reg __421348_421348;
   reg _421349_421349 ; 
   reg __421349_421349;
   reg _421350_421350 ; 
   reg __421350_421350;
   reg _421351_421351 ; 
   reg __421351_421351;
   reg _421352_421352 ; 
   reg __421352_421352;
   reg _421353_421353 ; 
   reg __421353_421353;
   reg _421354_421354 ; 
   reg __421354_421354;
   reg _421355_421355 ; 
   reg __421355_421355;
   reg _421356_421356 ; 
   reg __421356_421356;
   reg _421357_421357 ; 
   reg __421357_421357;
   reg _421358_421358 ; 
   reg __421358_421358;
   reg _421359_421359 ; 
   reg __421359_421359;
   reg _421360_421360 ; 
   reg __421360_421360;
   reg _421361_421361 ; 
   reg __421361_421361;
   reg _421362_421362 ; 
   reg __421362_421362;
   reg _421363_421363 ; 
   reg __421363_421363;
   reg _421364_421364 ; 
   reg __421364_421364;
   reg _421365_421365 ; 
   reg __421365_421365;
   reg _421366_421366 ; 
   reg __421366_421366;
   reg _421367_421367 ; 
   reg __421367_421367;
   reg _421368_421368 ; 
   reg __421368_421368;
   reg _421369_421369 ; 
   reg __421369_421369;
   reg _421370_421370 ; 
   reg __421370_421370;
   reg _421371_421371 ; 
   reg __421371_421371;
   reg _421372_421372 ; 
   reg __421372_421372;
   reg _421373_421373 ; 
   reg __421373_421373;
   reg _421374_421374 ; 
   reg __421374_421374;
   reg _421375_421375 ; 
   reg __421375_421375;
   reg _421376_421376 ; 
   reg __421376_421376;
   reg _421377_421377 ; 
   reg __421377_421377;
   reg _421378_421378 ; 
   reg __421378_421378;
   reg _421379_421379 ; 
   reg __421379_421379;
   reg _421380_421380 ; 
   reg __421380_421380;
   reg _421381_421381 ; 
   reg __421381_421381;
   reg _421382_421382 ; 
   reg __421382_421382;
   reg _421383_421383 ; 
   reg __421383_421383;
   reg _421384_421384 ; 
   reg __421384_421384;
   reg _421385_421385 ; 
   reg __421385_421385;
   reg _421386_421386 ; 
   reg __421386_421386;
   reg _421387_421387 ; 
   reg __421387_421387;
   reg _421388_421388 ; 
   reg __421388_421388;
   reg _421389_421389 ; 
   reg __421389_421389;
   reg _421390_421390 ; 
   reg __421390_421390;
   reg _421391_421391 ; 
   reg __421391_421391;
   reg _421392_421392 ; 
   reg __421392_421392;
   reg _421393_421393 ; 
   reg __421393_421393;
   reg _421394_421394 ; 
   reg __421394_421394;
   reg _421395_421395 ; 
   reg __421395_421395;
   reg _421396_421396 ; 
   reg __421396_421396;
   reg _421397_421397 ; 
   reg __421397_421397;
   reg _421398_421398 ; 
   reg __421398_421398;
   reg _421399_421399 ; 
   reg __421399_421399;
   reg _421400_421400 ; 
   reg __421400_421400;
   reg _421401_421401 ; 
   reg __421401_421401;
   reg _421402_421402 ; 
   reg __421402_421402;
   reg _421403_421403 ; 
   reg __421403_421403;
   reg _421404_421404 ; 
   reg __421404_421404;
   reg _421405_421405 ; 
   reg __421405_421405;
   reg _421406_421406 ; 
   reg __421406_421406;
   reg _421407_421407 ; 
   reg __421407_421407;
   reg _421408_421408 ; 
   reg __421408_421408;
   reg _421409_421409 ; 
   reg __421409_421409;
   reg _421410_421410 ; 
   reg __421410_421410;
   reg _421411_421411 ; 
   reg __421411_421411;
   reg _421412_421412 ; 
   reg __421412_421412;
   reg _421413_421413 ; 
   reg __421413_421413;
   reg _421414_421414 ; 
   reg __421414_421414;
   reg _421415_421415 ; 
   reg __421415_421415;
   reg _421416_421416 ; 
   reg __421416_421416;
   reg _421417_421417 ; 
   reg __421417_421417;
   reg _421418_421418 ; 
   reg __421418_421418;
   reg _421419_421419 ; 
   reg __421419_421419;
   reg _421420_421420 ; 
   reg __421420_421420;
   reg _421421_421421 ; 
   reg __421421_421421;
   reg _421422_421422 ; 
   reg __421422_421422;
   reg _421423_421423 ; 
   reg __421423_421423;
   reg _421424_421424 ; 
   reg __421424_421424;
   reg _421425_421425 ; 
   reg __421425_421425;
   reg _421426_421426 ; 
   reg __421426_421426;
   reg _421427_421427 ; 
   reg __421427_421427;
   reg _421428_421428 ; 
   reg __421428_421428;
   reg _421429_421429 ; 
   reg __421429_421429;
   reg _421430_421430 ; 
   reg __421430_421430;
   reg _421431_421431 ; 
   reg __421431_421431;
   reg _421432_421432 ; 
   reg __421432_421432;
   reg _421433_421433 ; 
   reg __421433_421433;
   reg _421434_421434 ; 
   reg __421434_421434;
   reg _421435_421435 ; 
   reg __421435_421435;
   reg _421436_421436 ; 
   reg __421436_421436;
   reg _421437_421437 ; 
   reg __421437_421437;
   reg _421438_421438 ; 
   reg __421438_421438;
   reg _421439_421439 ; 
   reg __421439_421439;
   reg _421440_421440 ; 
   reg __421440_421440;
   reg _421441_421441 ; 
   reg __421441_421441;
   reg _421442_421442 ; 
   reg __421442_421442;
   reg _421443_421443 ; 
   reg __421443_421443;
   reg _421444_421444 ; 
   reg __421444_421444;
   reg _421445_421445 ; 
   reg __421445_421445;
   reg _421446_421446 ; 
   reg __421446_421446;
   reg _421447_421447 ; 
   reg __421447_421447;
   reg _421448_421448 ; 
   reg __421448_421448;
   reg _421449_421449 ; 
   reg __421449_421449;
   reg _421450_421450 ; 
   reg __421450_421450;
   reg _421451_421451 ; 
   reg __421451_421451;
   reg _421452_421452 ; 
   reg __421452_421452;
   reg _421453_421453 ; 
   reg __421453_421453;
   reg _421454_421454 ; 
   reg __421454_421454;
   reg _421455_421455 ; 
   reg __421455_421455;
   reg _421456_421456 ; 
   reg __421456_421456;
   reg _421457_421457 ; 
   reg __421457_421457;
   reg _421458_421458 ; 
   reg __421458_421458;
   reg _421459_421459 ; 
   reg __421459_421459;
   reg _421460_421460 ; 
   reg __421460_421460;
   reg _421461_421461 ; 
   reg __421461_421461;
   reg _421462_421462 ; 
   reg __421462_421462;
   reg _421463_421463 ; 
   reg __421463_421463;
   reg _421464_421464 ; 
   reg __421464_421464;
   reg _421465_421465 ; 
   reg __421465_421465;
   reg _421466_421466 ; 
   reg __421466_421466;
   reg _421467_421467 ; 
   reg __421467_421467;
   reg _421468_421468 ; 
   reg __421468_421468;
   reg _421469_421469 ; 
   reg __421469_421469;
   reg _421470_421470 ; 
   reg __421470_421470;
   reg _421471_421471 ; 
   reg __421471_421471;
   reg _421472_421472 ; 
   reg __421472_421472;
   reg _421473_421473 ; 
   reg __421473_421473;
   reg _421474_421474 ; 
   reg __421474_421474;
   reg _421475_421475 ; 
   reg __421475_421475;
   reg _421476_421476 ; 
   reg __421476_421476;
   reg _421477_421477 ; 
   reg __421477_421477;
   reg _421478_421478 ; 
   reg __421478_421478;
   reg _421479_421479 ; 
   reg __421479_421479;
   reg _421480_421480 ; 
   reg __421480_421480;
   reg _421481_421481 ; 
   reg __421481_421481;
   reg _421482_421482 ; 
   reg __421482_421482;
   reg _421483_421483 ; 
   reg __421483_421483;
   reg _421484_421484 ; 
   reg __421484_421484;
   reg _421485_421485 ; 
   reg __421485_421485;
   reg _421486_421486 ; 
   reg __421486_421486;
   reg _421487_421487 ; 
   reg __421487_421487;
   reg _421488_421488 ; 
   reg __421488_421488;
   reg _421489_421489 ; 
   reg __421489_421489;
   reg _421490_421490 ; 
   reg __421490_421490;
   reg _421491_421491 ; 
   reg __421491_421491;
   reg _421492_421492 ; 
   reg __421492_421492;
   reg _421493_421493 ; 
   reg __421493_421493;
   reg _421494_421494 ; 
   reg __421494_421494;
   reg _421495_421495 ; 
   reg __421495_421495;
   reg _421496_421496 ; 
   reg __421496_421496;
   reg _421497_421497 ; 
   reg __421497_421497;
   reg _421498_421498 ; 
   reg __421498_421498;
   reg _421499_421499 ; 
   reg __421499_421499;
   reg _421500_421500 ; 
   reg __421500_421500;
   reg _421501_421501 ; 
   reg __421501_421501;
   reg _421502_421502 ; 
   reg __421502_421502;
   reg _421503_421503 ; 
   reg __421503_421503;
   reg _421504_421504 ; 
   reg __421504_421504;
   reg _421505_421505 ; 
   reg __421505_421505;
   reg _421506_421506 ; 
   reg __421506_421506;
   reg _421507_421507 ; 
   reg __421507_421507;
   reg _421508_421508 ; 
   reg __421508_421508;
   reg _421509_421509 ; 
   reg __421509_421509;
   reg _421510_421510 ; 
   reg __421510_421510;
   reg _421511_421511 ; 
   reg __421511_421511;
   reg _421512_421512 ; 
   reg __421512_421512;
   reg _421513_421513 ; 
   reg __421513_421513;
   reg _421514_421514 ; 
   reg __421514_421514;
   reg _421515_421515 ; 
   reg __421515_421515;
   reg _421516_421516 ; 
   reg __421516_421516;
   reg _421517_421517 ; 
   reg __421517_421517;
   reg _421518_421518 ; 
   reg __421518_421518;
   reg _421519_421519 ; 
   reg __421519_421519;
   reg _421520_421520 ; 
   reg __421520_421520;
   reg _421521_421521 ; 
   reg __421521_421521;
   reg _421522_421522 ; 
   reg __421522_421522;
   reg _421523_421523 ; 
   reg __421523_421523;
   reg _421524_421524 ; 
   reg __421524_421524;
   reg _421525_421525 ; 
   reg __421525_421525;
   reg _421526_421526 ; 
   reg __421526_421526;
   reg _421527_421527 ; 
   reg __421527_421527;
   reg _421528_421528 ; 
   reg __421528_421528;
   reg _421529_421529 ; 
   reg __421529_421529;
   reg _421530_421530 ; 
   reg __421530_421530;
   reg _421531_421531 ; 
   reg __421531_421531;
   reg _421532_421532 ; 
   reg __421532_421532;
   reg _421533_421533 ; 
   reg __421533_421533;
   reg _421534_421534 ; 
   reg __421534_421534;
   reg _421535_421535 ; 
   reg __421535_421535;
   reg _421536_421536 ; 
   reg __421536_421536;
   reg _421537_421537 ; 
   reg __421537_421537;
   reg _421538_421538 ; 
   reg __421538_421538;
   reg _421539_421539 ; 
   reg __421539_421539;
   reg _421540_421540 ; 
   reg __421540_421540;
   reg _421541_421541 ; 
   reg __421541_421541;
   reg _421542_421542 ; 
   reg __421542_421542;
   reg _421543_421543 ; 
   reg __421543_421543;
   reg _421544_421544 ; 
   reg __421544_421544;
   reg _421545_421545 ; 
   reg __421545_421545;
   reg _421546_421546 ; 
   reg __421546_421546;
   reg _421547_421547 ; 
   reg __421547_421547;
   reg _421548_421548 ; 
   reg __421548_421548;
   reg _421549_421549 ; 
   reg __421549_421549;
   reg _421550_421550 ; 
   reg __421550_421550;
   reg _421551_421551 ; 
   reg __421551_421551;
   reg _421552_421552 ; 
   reg __421552_421552;
   reg _421553_421553 ; 
   reg __421553_421553;
   reg _421554_421554 ; 
   reg __421554_421554;
   reg _421555_421555 ; 
   reg __421555_421555;
   reg _421556_421556 ; 
   reg __421556_421556;
   reg _421557_421557 ; 
   reg __421557_421557;
   reg _421558_421558 ; 
   reg __421558_421558;
   reg _421559_421559 ; 
   reg __421559_421559;
   reg _421560_421560 ; 
   reg __421560_421560;
   reg _421561_421561 ; 
   reg __421561_421561;
   reg _421562_421562 ; 
   reg __421562_421562;
   reg _421563_421563 ; 
   reg __421563_421563;
   reg _421564_421564 ; 
   reg __421564_421564;
   reg _421565_421565 ; 
   reg __421565_421565;
   reg _421566_421566 ; 
   reg __421566_421566;
   reg _421567_421567 ; 
   reg __421567_421567;
   reg _421568_421568 ; 
   reg __421568_421568;
   reg _421569_421569 ; 
   reg __421569_421569;
   reg _421570_421570 ; 
   reg __421570_421570;
   reg _421571_421571 ; 
   reg __421571_421571;
   reg _421572_421572 ; 
   reg __421572_421572;
   reg _421573_421573 ; 
   reg __421573_421573;
   reg _421574_421574 ; 
   reg __421574_421574;
   reg _421575_421575 ; 
   reg __421575_421575;
   reg _421576_421576 ; 
   reg __421576_421576;
   reg _421577_421577 ; 
   reg __421577_421577;
   reg _421578_421578 ; 
   reg __421578_421578;
   reg _421579_421579 ; 
   reg __421579_421579;
   reg _421580_421580 ; 
   reg __421580_421580;
   reg _421581_421581 ; 
   reg __421581_421581;
   reg _421582_421582 ; 
   reg __421582_421582;
   reg _421583_421583 ; 
   reg __421583_421583;
   reg _421584_421584 ; 
   reg __421584_421584;
   reg _421585_421585 ; 
   reg __421585_421585;
   reg _421586_421586 ; 
   reg __421586_421586;
   reg _421587_421587 ; 
   reg __421587_421587;
   reg _421588_421588 ; 
   reg __421588_421588;
   reg _421589_421589 ; 
   reg __421589_421589;
   reg _421590_421590 ; 
   reg __421590_421590;
   reg _421591_421591 ; 
   reg __421591_421591;
   reg _421592_421592 ; 
   reg __421592_421592;
   reg _421593_421593 ; 
   reg __421593_421593;
   reg _421594_421594 ; 
   reg __421594_421594;
   reg _421595_421595 ; 
   reg __421595_421595;
   reg _421596_421596 ; 
   reg __421596_421596;
   reg _421597_421597 ; 
   reg __421597_421597;
   reg _421598_421598 ; 
   reg __421598_421598;
   reg _421599_421599 ; 
   reg __421599_421599;
   reg _421600_421600 ; 
   reg __421600_421600;
   reg _421601_421601 ; 
   reg __421601_421601;
   reg _421602_421602 ; 
   reg __421602_421602;
   reg _421603_421603 ; 
   reg __421603_421603;
   reg _421604_421604 ; 
   reg __421604_421604;
   reg _421605_421605 ; 
   reg __421605_421605;
   reg _421606_421606 ; 
   reg __421606_421606;
   reg _421607_421607 ; 
   reg __421607_421607;
   reg _421608_421608 ; 
   reg __421608_421608;
   reg _421609_421609 ; 
   reg __421609_421609;
   reg _421610_421610 ; 
   reg __421610_421610;
   reg _421611_421611 ; 
   reg __421611_421611;
   reg _421612_421612 ; 
   reg __421612_421612;
   reg _421613_421613 ; 
   reg __421613_421613;
   reg _421614_421614 ; 
   reg __421614_421614;
   reg _421615_421615 ; 
   reg __421615_421615;
   reg _421616_421616 ; 
   reg __421616_421616;
   reg _421617_421617 ; 
   reg __421617_421617;
   reg _421618_421618 ; 
   reg __421618_421618;
   reg _421619_421619 ; 
   reg __421619_421619;
   reg _421620_421620 ; 
   reg __421620_421620;
   reg _421621_421621 ; 
   reg __421621_421621;
   reg _421622_421622 ; 
   reg __421622_421622;
   reg _421623_421623 ; 
   reg __421623_421623;
   reg _421624_421624 ; 
   reg __421624_421624;
   reg _421625_421625 ; 
   reg __421625_421625;
   reg _421626_421626 ; 
   reg __421626_421626;
   reg _421627_421627 ; 
   reg __421627_421627;
   reg _421628_421628 ; 
   reg __421628_421628;
   reg _421629_421629 ; 
   reg __421629_421629;
   reg _421630_421630 ; 
   reg __421630_421630;
   reg _421631_421631 ; 
   reg __421631_421631;
   reg _421632_421632 ; 
   reg __421632_421632;
   reg _421633_421633 ; 
   reg __421633_421633;
   reg _421634_421634 ; 
   reg __421634_421634;
   reg _421635_421635 ; 
   reg __421635_421635;
   reg _421636_421636 ; 
   reg __421636_421636;
   reg _421637_421637 ; 
   reg __421637_421637;
   reg _421638_421638 ; 
   reg __421638_421638;
   reg _421639_421639 ; 
   reg __421639_421639;
   reg _421640_421640 ; 
   reg __421640_421640;
   reg _421641_421641 ; 
   reg __421641_421641;
   reg _421642_421642 ; 
   reg __421642_421642;
   reg _421643_421643 ; 
   reg __421643_421643;
   reg _421644_421644 ; 
   reg __421644_421644;
   reg _421645_421645 ; 
   reg __421645_421645;
   reg _421646_421646 ; 
   reg __421646_421646;
   reg _421647_421647 ; 
   reg __421647_421647;
   reg _421648_421648 ; 
   reg __421648_421648;
   reg _421649_421649 ; 
   reg __421649_421649;
   reg _421650_421650 ; 
   reg __421650_421650;
   reg _421651_421651 ; 
   reg __421651_421651;
   reg _421652_421652 ; 
   reg __421652_421652;
   reg _421653_421653 ; 
   reg __421653_421653;
   reg _421654_421654 ; 
   reg __421654_421654;
   reg _421655_421655 ; 
   reg __421655_421655;
   reg _421656_421656 ; 
   reg __421656_421656;
   reg _421657_421657 ; 
   reg __421657_421657;
   reg _421658_421658 ; 
   reg __421658_421658;
   reg _421659_421659 ; 
   reg __421659_421659;
   reg _421660_421660 ; 
   reg __421660_421660;
   reg _421661_421661 ; 
   reg __421661_421661;
   reg _421662_421662 ; 
   reg __421662_421662;
   reg _421663_421663 ; 
   reg __421663_421663;
   reg _421664_421664 ; 
   reg __421664_421664;
   reg _421665_421665 ; 
   reg __421665_421665;
   reg _421666_421666 ; 
   reg __421666_421666;
   reg _421667_421667 ; 
   reg __421667_421667;
   reg _421668_421668 ; 
   reg __421668_421668;
   reg _421669_421669 ; 
   reg __421669_421669;
   reg _421670_421670 ; 
   reg __421670_421670;
   reg _421671_421671 ; 
   reg __421671_421671;
   reg _421672_421672 ; 
   reg __421672_421672;
   reg _421673_421673 ; 
   reg __421673_421673;
   reg _421674_421674 ; 
   reg __421674_421674;
   reg _421675_421675 ; 
   reg __421675_421675;
   reg _421676_421676 ; 
   reg __421676_421676;
   reg _421677_421677 ; 
   reg __421677_421677;
   reg _421678_421678 ; 
   reg __421678_421678;
   reg _421679_421679 ; 
   reg __421679_421679;
   reg _421680_421680 ; 
   reg __421680_421680;
   reg _421681_421681 ; 
   reg __421681_421681;
   reg _421682_421682 ; 
   reg __421682_421682;
   reg _421683_421683 ; 
   reg __421683_421683;
   reg _421684_421684 ; 
   reg __421684_421684;
   reg _421685_421685 ; 
   reg __421685_421685;
   reg _421686_421686 ; 
   reg __421686_421686;
   reg _421687_421687 ; 
   reg __421687_421687;
   reg _421688_421688 ; 
   reg __421688_421688;
   reg _421689_421689 ; 
   reg __421689_421689;
   reg _421690_421690 ; 
   reg __421690_421690;
   reg _421691_421691 ; 
   reg __421691_421691;
   reg _421692_421692 ; 
   reg __421692_421692;
   reg _421693_421693 ; 
   reg __421693_421693;
   reg _421694_421694 ; 
   reg __421694_421694;
   reg _421695_421695 ; 
   reg __421695_421695;
   reg _421696_421696 ; 
   reg __421696_421696;
   reg _421697_421697 ; 
   reg __421697_421697;
   reg _421698_421698 ; 
   reg __421698_421698;
   reg _421699_421699 ; 
   reg __421699_421699;
   reg _421700_421700 ; 
   reg __421700_421700;
   reg _421701_421701 ; 
   reg __421701_421701;
   reg _421702_421702 ; 
   reg __421702_421702;
   reg _421703_421703 ; 
   reg __421703_421703;
   reg _421704_421704 ; 
   reg __421704_421704;
   reg _421705_421705 ; 
   reg __421705_421705;
   reg _421706_421706 ; 
   reg __421706_421706;
   reg _421707_421707 ; 
   reg __421707_421707;
   reg _421708_421708 ; 
   reg __421708_421708;
   reg _421709_421709 ; 
   reg __421709_421709;
   reg _421710_421710 ; 
   reg __421710_421710;
   reg _421711_421711 ; 
   reg __421711_421711;
   reg _421712_421712 ; 
   reg __421712_421712;
   reg _421713_421713 ; 
   reg __421713_421713;
   reg _421714_421714 ; 
   reg __421714_421714;
   reg _421715_421715 ; 
   reg __421715_421715;
   reg _421716_421716 ; 
   reg __421716_421716;
   reg _421717_421717 ; 
   reg __421717_421717;
   reg _421718_421718 ; 
   reg __421718_421718;
   reg _421719_421719 ; 
   reg __421719_421719;
   reg _421720_421720 ; 
   reg __421720_421720;
   reg _421721_421721 ; 
   reg __421721_421721;
   reg _421722_421722 ; 
   reg __421722_421722;
   reg _421723_421723 ; 
   reg __421723_421723;
   reg _421724_421724 ; 
   reg __421724_421724;
   reg _421725_421725 ; 
   reg __421725_421725;
   reg _421726_421726 ; 
   reg __421726_421726;
   reg _421727_421727 ; 
   reg __421727_421727;
   reg _421728_421728 ; 
   reg __421728_421728;
   reg _421729_421729 ; 
   reg __421729_421729;
   reg _421730_421730 ; 
   reg __421730_421730;
   reg _421731_421731 ; 
   reg __421731_421731;
   reg _421732_421732 ; 
   reg __421732_421732;
   reg _421733_421733 ; 
   reg __421733_421733;
   reg _421734_421734 ; 
   reg __421734_421734;
   reg _421735_421735 ; 
   reg __421735_421735;
   reg _421736_421736 ; 
   reg __421736_421736;
   reg _421737_421737 ; 
   reg __421737_421737;
   reg _421738_421738 ; 
   reg __421738_421738;
   reg _421739_421739 ; 
   reg __421739_421739;
   reg _421740_421740 ; 
   reg __421740_421740;
   reg _421741_421741 ; 
   reg __421741_421741;
   reg _421742_421742 ; 
   reg __421742_421742;
   reg _421743_421743 ; 
   reg __421743_421743;
   reg _421744_421744 ; 
   reg __421744_421744;
   reg _421745_421745 ; 
   reg __421745_421745;
   reg _421746_421746 ; 
   reg __421746_421746;
   reg _421747_421747 ; 
   reg __421747_421747;
   reg _421748_421748 ; 
   reg __421748_421748;
   reg _421749_421749 ; 
   reg __421749_421749;
   reg _421750_421750 ; 
   reg __421750_421750;
   reg _421751_421751 ; 
   reg __421751_421751;
   reg _421752_421752 ; 
   reg __421752_421752;
   reg _421753_421753 ; 
   reg __421753_421753;
   reg _421754_421754 ; 
   reg __421754_421754;
   reg _421755_421755 ; 
   reg __421755_421755;
   reg _421756_421756 ; 
   reg __421756_421756;
   reg _421757_421757 ; 
   reg __421757_421757;
   reg _421758_421758 ; 
   reg __421758_421758;
   reg _421759_421759 ; 
   reg __421759_421759;
   reg _421760_421760 ; 
   reg __421760_421760;
   reg _421761_421761 ; 
   reg __421761_421761;
   reg _421762_421762 ; 
   reg __421762_421762;
   reg _421763_421763 ; 
   reg __421763_421763;
   reg _421764_421764 ; 
   reg __421764_421764;
   reg _421765_421765 ; 
   reg __421765_421765;
   reg _421766_421766 ; 
   reg __421766_421766;
   reg _421767_421767 ; 
   reg __421767_421767;
   reg _421768_421768 ; 
   reg __421768_421768;
   reg _421769_421769 ; 
   reg __421769_421769;
   reg _421770_421770 ; 
   reg __421770_421770;
   reg _421771_421771 ; 
   reg __421771_421771;
   reg _421772_421772 ; 
   reg __421772_421772;
   reg _421773_421773 ; 
   reg __421773_421773;
   reg _421774_421774 ; 
   reg __421774_421774;
   reg _421775_421775 ; 
   reg __421775_421775;
   reg _421776_421776 ; 
   reg __421776_421776;
   reg _421777_421777 ; 
   reg __421777_421777;
   reg _421778_421778 ; 
   reg __421778_421778;
   reg _421779_421779 ; 
   reg __421779_421779;
   reg _421780_421780 ; 
   reg __421780_421780;
   reg _421781_421781 ; 
   reg __421781_421781;
   reg _421782_421782 ; 
   reg __421782_421782;
   reg _421783_421783 ; 
   reg __421783_421783;
   reg _421784_421784 ; 
   reg __421784_421784;
   reg _421785_421785 ; 
   reg __421785_421785;
   reg _421786_421786 ; 
   reg __421786_421786;
   reg _421787_421787 ; 
   reg __421787_421787;
   reg _421788_421788 ; 
   reg __421788_421788;
   reg _421789_421789 ; 
   reg __421789_421789;
   reg _421790_421790 ; 
   reg __421790_421790;
   reg _421791_421791 ; 
   reg __421791_421791;
   reg _421792_421792 ; 
   reg __421792_421792;
   reg _421793_421793 ; 
   reg __421793_421793;
   reg _421794_421794 ; 
   reg __421794_421794;
   reg _421795_421795 ; 
   reg __421795_421795;
   reg _421796_421796 ; 
   reg __421796_421796;
   reg _421797_421797 ; 
   reg __421797_421797;
   reg _421798_421798 ; 
   reg __421798_421798;
   reg _421799_421799 ; 
   reg __421799_421799;
   reg _421800_421800 ; 
   reg __421800_421800;
   reg _421801_421801 ; 
   reg __421801_421801;
   reg _421802_421802 ; 
   reg __421802_421802;
   reg _421803_421803 ; 
   reg __421803_421803;
   reg _421804_421804 ; 
   reg __421804_421804;
   reg _421805_421805 ; 
   reg __421805_421805;
   reg _421806_421806 ; 
   reg __421806_421806;
   reg _421807_421807 ; 
   reg __421807_421807;
   reg _421808_421808 ; 
   reg __421808_421808;
   reg _421809_421809 ; 
   reg __421809_421809;
   reg _421810_421810 ; 
   reg __421810_421810;
   reg _421811_421811 ; 
   reg __421811_421811;
   reg _421812_421812 ; 
   reg __421812_421812;
   reg _421813_421813 ; 
   reg __421813_421813;
   reg _421814_421814 ; 
   reg __421814_421814;
   reg _421815_421815 ; 
   reg __421815_421815;
   reg _421816_421816 ; 
   reg __421816_421816;
   reg _421817_421817 ; 
   reg __421817_421817;
   reg _421818_421818 ; 
   reg __421818_421818;
   reg _421819_421819 ; 
   reg __421819_421819;
   reg _421820_421820 ; 
   reg __421820_421820;
   reg _421821_421821 ; 
   reg __421821_421821;
   reg _421822_421822 ; 
   reg __421822_421822;
   reg _421823_421823 ; 
   reg __421823_421823;
   reg _421824_421824 ; 
   reg __421824_421824;
   reg _421825_421825 ; 
   reg __421825_421825;
   reg _421826_421826 ; 
   reg __421826_421826;
   reg _421827_421827 ; 
   reg __421827_421827;
   reg _421828_421828 ; 
   reg __421828_421828;
   reg _421829_421829 ; 
   reg __421829_421829;
   reg _421830_421830 ; 
   reg __421830_421830;
   reg _421831_421831 ; 
   reg __421831_421831;
   reg _421832_421832 ; 
   reg __421832_421832;
   reg _421833_421833 ; 
   reg __421833_421833;
   reg _421834_421834 ; 
   reg __421834_421834;
   reg _421835_421835 ; 
   reg __421835_421835;
   reg _421836_421836 ; 
   reg __421836_421836;
   reg _421837_421837 ; 
   reg __421837_421837;
   reg _421838_421838 ; 
   reg __421838_421838;
   reg _421839_421839 ; 
   reg __421839_421839;
   reg _421840_421840 ; 
   reg __421840_421840;
   reg _421841_421841 ; 
   reg __421841_421841;
   reg _421842_421842 ; 
   reg __421842_421842;
   reg _421843_421843 ; 
   reg __421843_421843;
   reg _421844_421844 ; 
   reg __421844_421844;
   reg _421845_421845 ; 
   reg __421845_421845;
   reg _421846_421846 ; 
   reg __421846_421846;
   reg _421847_421847 ; 
   reg __421847_421847;
   reg _421848_421848 ; 
   reg __421848_421848;
   reg _421849_421849 ; 
   reg __421849_421849;
   reg _421850_421850 ; 
   reg __421850_421850;
   reg _421851_421851 ; 
   reg __421851_421851;
   reg _421852_421852 ; 
   reg __421852_421852;
   reg _421853_421853 ; 
   reg __421853_421853;
   reg _421854_421854 ; 
   reg __421854_421854;
   reg _421855_421855 ; 
   reg __421855_421855;
   reg _421856_421856 ; 
   reg __421856_421856;
   reg _421857_421857 ; 
   reg __421857_421857;
   reg _421858_421858 ; 
   reg __421858_421858;
   reg _421859_421859 ; 
   reg __421859_421859;
   reg _421860_421860 ; 
   reg __421860_421860;
   reg _421861_421861 ; 
   reg __421861_421861;
   reg _421862_421862 ; 
   reg __421862_421862;
   reg _421863_421863 ; 
   reg __421863_421863;
   reg _421864_421864 ; 
   reg __421864_421864;
   reg _421865_421865 ; 
   reg __421865_421865;
   reg _421866_421866 ; 
   reg __421866_421866;
   reg _421867_421867 ; 
   reg __421867_421867;
   reg _421868_421868 ; 
   reg __421868_421868;
   reg _421869_421869 ; 
   reg __421869_421869;
   reg _421870_421870 ; 
   reg __421870_421870;
   reg _421871_421871 ; 
   reg __421871_421871;
   reg _421872_421872 ; 
   reg __421872_421872;
   reg _421873_421873 ; 
   reg __421873_421873;
   reg _421874_421874 ; 
   reg __421874_421874;
   reg _421875_421875 ; 
   reg __421875_421875;
   reg _421876_421876 ; 
   reg __421876_421876;
   reg _421877_421877 ; 
   reg __421877_421877;
   reg _421878_421878 ; 
   reg __421878_421878;
   reg _421879_421879 ; 
   reg __421879_421879;
   reg _421880_421880 ; 
   reg __421880_421880;
   reg _421881_421881 ; 
   reg __421881_421881;
   reg _421882_421882 ; 
   reg __421882_421882;
   reg _421883_421883 ; 
   reg __421883_421883;
   reg _421884_421884 ; 
   reg __421884_421884;
   reg _421885_421885 ; 
   reg __421885_421885;
   reg _421886_421886 ; 
   reg __421886_421886;
   reg _421887_421887 ; 
   reg __421887_421887;
   reg _421888_421888 ; 
   reg __421888_421888;
   reg _421889_421889 ; 
   reg __421889_421889;
   reg _421890_421890 ; 
   reg __421890_421890;
   reg _421891_421891 ; 
   reg __421891_421891;
   reg _421892_421892 ; 
   reg __421892_421892;
   reg _421893_421893 ; 
   reg __421893_421893;
   reg _421894_421894 ; 
   reg __421894_421894;
   reg _421895_421895 ; 
   reg __421895_421895;
   reg _421896_421896 ; 
   reg __421896_421896;
   reg _421897_421897 ; 
   reg __421897_421897;
   reg _421898_421898 ; 
   reg __421898_421898;
   reg _421899_421899 ; 
   reg __421899_421899;
   reg _421900_421900 ; 
   reg __421900_421900;
   reg _421901_421901 ; 
   reg __421901_421901;
   reg _421902_421902 ; 
   reg __421902_421902;
   reg _421903_421903 ; 
   reg __421903_421903;
   reg _421904_421904 ; 
   reg __421904_421904;
   reg _421905_421905 ; 
   reg __421905_421905;
   reg _421906_421906 ; 
   reg __421906_421906;
   reg _421907_421907 ; 
   reg __421907_421907;
   reg _421908_421908 ; 
   reg __421908_421908;
   reg _421909_421909 ; 
   reg __421909_421909;
   reg _421910_421910 ; 
   reg __421910_421910;
   reg _421911_421911 ; 
   reg __421911_421911;
   reg _421912_421912 ; 
   reg __421912_421912;
   reg _421913_421913 ; 
   reg __421913_421913;
   reg _421914_421914 ; 
   reg __421914_421914;
   reg _421915_421915 ; 
   reg __421915_421915;
   reg _421916_421916 ; 
   reg __421916_421916;
   reg _421917_421917 ; 
   reg __421917_421917;
   reg _421918_421918 ; 
   reg __421918_421918;
   reg _421919_421919 ; 
   reg __421919_421919;
   reg _421920_421920 ; 
   reg __421920_421920;
   reg _421921_421921 ; 
   reg __421921_421921;
   reg _421922_421922 ; 
   reg __421922_421922;
   reg _421923_421923 ; 
   reg __421923_421923;
   reg _421924_421924 ; 
   reg __421924_421924;
   reg _421925_421925 ; 
   reg __421925_421925;
   reg _421926_421926 ; 
   reg __421926_421926;
   reg _421927_421927 ; 
   reg __421927_421927;
   reg _421928_421928 ; 
   reg __421928_421928;
   reg _421929_421929 ; 
   reg __421929_421929;
   reg _421930_421930 ; 
   reg __421930_421930;
   reg _421931_421931 ; 
   reg __421931_421931;
   reg _421932_421932 ; 
   reg __421932_421932;
   reg _421933_421933 ; 
   reg __421933_421933;
   reg _421934_421934 ; 
   reg __421934_421934;
   reg _421935_421935 ; 
   reg __421935_421935;
   reg _421936_421936 ; 
   reg __421936_421936;
   reg _421937_421937 ; 
   reg __421937_421937;
   reg _421938_421938 ; 
   reg __421938_421938;
   reg _421939_421939 ; 
   reg __421939_421939;
   reg _421940_421940 ; 
   reg __421940_421940;
   reg _421941_421941 ; 
   reg __421941_421941;
   reg _421942_421942 ; 
   reg __421942_421942;
   reg _421943_421943 ; 
   reg __421943_421943;
   reg _421944_421944 ; 
   reg __421944_421944;
   reg _421945_421945 ; 
   reg __421945_421945;
   reg _421946_421946 ; 
   reg __421946_421946;
   reg _421947_421947 ; 
   reg __421947_421947;
   reg _421948_421948 ; 
   reg __421948_421948;
   reg _421949_421949 ; 
   reg __421949_421949;
   reg _421950_421950 ; 
   reg __421950_421950;
   reg _421951_421951 ; 
   reg __421951_421951;
   reg _421952_421952 ; 
   reg __421952_421952;
   reg _421953_421953 ; 
   reg __421953_421953;
   reg _421954_421954 ; 
   reg __421954_421954;
   reg _421955_421955 ; 
   reg __421955_421955;
   reg _421956_421956 ; 
   reg __421956_421956;
   reg _421957_421957 ; 
   reg __421957_421957;
   reg _421958_421958 ; 
   reg __421958_421958;
   reg _421959_421959 ; 
   reg __421959_421959;
   reg _421960_421960 ; 
   reg __421960_421960;
   reg _421961_421961 ; 
   reg __421961_421961;
   reg _421962_421962 ; 
   reg __421962_421962;
   reg _421963_421963 ; 
   reg __421963_421963;
   reg _421964_421964 ; 
   reg __421964_421964;
   reg _421965_421965 ; 
   reg __421965_421965;
   reg _421966_421966 ; 
   reg __421966_421966;
   reg _421967_421967 ; 
   reg __421967_421967;
   reg _421968_421968 ; 
   reg __421968_421968;
   reg _421969_421969 ; 
   reg __421969_421969;
   reg _421970_421970 ; 
   reg __421970_421970;
   reg _421971_421971 ; 
   reg __421971_421971;
   reg _421972_421972 ; 
   reg __421972_421972;
   reg _421973_421973 ; 
   reg __421973_421973;
   reg _421974_421974 ; 
   reg __421974_421974;
   reg _421975_421975 ; 
   reg __421975_421975;
   reg _421976_421976 ; 
   reg __421976_421976;
   reg _421977_421977 ; 
   reg __421977_421977;
   reg _421978_421978 ; 
   reg __421978_421978;
   reg _421979_421979 ; 
   reg __421979_421979;
   reg _421980_421980 ; 
   reg __421980_421980;
   reg _421981_421981 ; 
   reg __421981_421981;
   reg _421982_421982 ; 
   reg __421982_421982;
   reg _421983_421983 ; 
   reg __421983_421983;
   reg _421984_421984 ; 
   reg __421984_421984;
   reg _421985_421985 ; 
   reg __421985_421985;
   reg _421986_421986 ; 
   reg __421986_421986;
   reg _421987_421987 ; 
   reg __421987_421987;
   reg _421988_421988 ; 
   reg __421988_421988;
   reg _421989_421989 ; 
   reg __421989_421989;
   reg _421990_421990 ; 
   reg __421990_421990;
   reg _421991_421991 ; 
   reg __421991_421991;
   reg _421992_421992 ; 
   reg __421992_421992;
   reg _421993_421993 ; 
   reg __421993_421993;
   reg _421994_421994 ; 
   reg __421994_421994;
   reg _421995_421995 ; 
   reg __421995_421995;
   reg _421996_421996 ; 
   reg __421996_421996;
   reg _421997_421997 ; 
   reg __421997_421997;
   reg _421998_421998 ; 
   reg __421998_421998;
   reg _421999_421999 ; 
   reg __421999_421999;
   reg _422000_422000 ; 
   reg __422000_422000;
   reg _422001_422001 ; 
   reg __422001_422001;
   reg _422002_422002 ; 
   reg __422002_422002;
   reg _422003_422003 ; 
   reg __422003_422003;
   reg _422004_422004 ; 
   reg __422004_422004;
   reg _422005_422005 ; 
   reg __422005_422005;
   reg _422006_422006 ; 
   reg __422006_422006;
   reg _422007_422007 ; 
   reg __422007_422007;
   reg _422008_422008 ; 
   reg __422008_422008;
   reg _422009_422009 ; 
   reg __422009_422009;
   reg _422010_422010 ; 
   reg __422010_422010;
   reg _422011_422011 ; 
   reg __422011_422011;
   reg _422012_422012 ; 
   reg __422012_422012;
   reg _422013_422013 ; 
   reg __422013_422013;
   reg _422014_422014 ; 
   reg __422014_422014;
   reg _422015_422015 ; 
   reg __422015_422015;
   reg _422016_422016 ; 
   reg __422016_422016;
   reg _422017_422017 ; 
   reg __422017_422017;
   reg _422018_422018 ; 
   reg __422018_422018;
   reg _422019_422019 ; 
   reg __422019_422019;
   reg _422020_422020 ; 
   reg __422020_422020;
   reg _422021_422021 ; 
   reg __422021_422021;
   reg _422022_422022 ; 
   reg __422022_422022;
   reg _422023_422023 ; 
   reg __422023_422023;
   reg _422024_422024 ; 
   reg __422024_422024;
   reg _422025_422025 ; 
   reg __422025_422025;
   reg _422026_422026 ; 
   reg __422026_422026;
   reg _422027_422027 ; 
   reg __422027_422027;
   reg _422028_422028 ; 
   reg __422028_422028;
   reg _422029_422029 ; 
   reg __422029_422029;
   reg _422030_422030 ; 
   reg __422030_422030;
   reg _422031_422031 ; 
   reg __422031_422031;
   reg _422032_422032 ; 
   reg __422032_422032;
   reg _422033_422033 ; 
   reg __422033_422033;
   reg _422034_422034 ; 
   reg __422034_422034;
   reg _422035_422035 ; 
   reg __422035_422035;
   reg _422036_422036 ; 
   reg __422036_422036;
   reg _422037_422037 ; 
   reg __422037_422037;
   reg _422038_422038 ; 
   reg __422038_422038;
   reg _422039_422039 ; 
   reg __422039_422039;
   reg _422040_422040 ; 
   reg __422040_422040;
   reg _422041_422041 ; 
   reg __422041_422041;
   reg _422042_422042 ; 
   reg __422042_422042;
   reg _422043_422043 ; 
   reg __422043_422043;
   reg _422044_422044 ; 
   reg __422044_422044;
   reg _422045_422045 ; 
   reg __422045_422045;
   reg _422046_422046 ; 
   reg __422046_422046;
   reg _422047_422047 ; 
   reg __422047_422047;
   reg _422048_422048 ; 
   reg __422048_422048;
   reg _422049_422049 ; 
   reg __422049_422049;
   reg _422050_422050 ; 
   reg __422050_422050;
   reg _422051_422051 ; 
   reg __422051_422051;
   reg _422052_422052 ; 
   reg __422052_422052;
   reg _422053_422053 ; 
   reg __422053_422053;
   reg _422054_422054 ; 
   reg __422054_422054;
   reg _422055_422055 ; 
   reg __422055_422055;
   reg _422056_422056 ; 
   reg __422056_422056;
   reg _422057_422057 ; 
   reg __422057_422057;
   reg _422058_422058 ; 
   reg __422058_422058;
   reg _422059_422059 ; 
   reg __422059_422059;
   reg _422060_422060 ; 
   reg __422060_422060;
   reg _422061_422061 ; 
   reg __422061_422061;
   reg _422062_422062 ; 
   reg __422062_422062;
   reg _422063_422063 ; 
   reg __422063_422063;
   reg _422064_422064 ; 
   reg __422064_422064;
   reg _422065_422065 ; 
   reg __422065_422065;
   reg _422066_422066 ; 
   reg __422066_422066;
   reg _422067_422067 ; 
   reg __422067_422067;
   reg _422068_422068 ; 
   reg __422068_422068;
   reg _422069_422069 ; 
   reg __422069_422069;
   reg _422070_422070 ; 
   reg __422070_422070;
   reg _422071_422071 ; 
   reg __422071_422071;
   reg _422072_422072 ; 
   reg __422072_422072;
   reg _422073_422073 ; 
   reg __422073_422073;
   reg _422074_422074 ; 
   reg __422074_422074;
   reg _422075_422075 ; 
   reg __422075_422075;
   reg _422076_422076 ; 
   reg __422076_422076;
   reg _422077_422077 ; 
   reg __422077_422077;
   reg _422078_422078 ; 
   reg __422078_422078;
   reg _422079_422079 ; 
   reg __422079_422079;
   reg _422080_422080 ; 
   reg __422080_422080;
   reg _422081_422081 ; 
   reg __422081_422081;
   reg _422082_422082 ; 
   reg __422082_422082;
   reg _422083_422083 ; 
   reg __422083_422083;
   reg _422084_422084 ; 
   reg __422084_422084;
   reg _422085_422085 ; 
   reg __422085_422085;
   reg _422086_422086 ; 
   reg __422086_422086;
   reg _422087_422087 ; 
   reg __422087_422087;
   reg _422088_422088 ; 
   reg __422088_422088;
   reg _422089_422089 ; 
   reg __422089_422089;
   reg _422090_422090 ; 
   reg __422090_422090;
   reg _422091_422091 ; 
   reg __422091_422091;
   reg _422092_422092 ; 
   reg __422092_422092;
   reg _422093_422093 ; 
   reg __422093_422093;
   reg _422094_422094 ; 
   reg __422094_422094;
   reg _422095_422095 ; 
   reg __422095_422095;
   reg _422096_422096 ; 
   reg __422096_422096;
   reg _422097_422097 ; 
   reg __422097_422097;
   reg _422098_422098 ; 
   reg __422098_422098;
   reg _422099_422099 ; 
   reg __422099_422099;
   reg _422100_422100 ; 
   reg __422100_422100;
   reg _422101_422101 ; 
   reg __422101_422101;
   reg _422102_422102 ; 
   reg __422102_422102;
   reg _422103_422103 ; 
   reg __422103_422103;
   reg _422104_422104 ; 
   reg __422104_422104;
   reg _422105_422105 ; 
   reg __422105_422105;
   reg _422106_422106 ; 
   reg __422106_422106;
   reg _422107_422107 ; 
   reg __422107_422107;
   reg _422108_422108 ; 
   reg __422108_422108;
   reg _422109_422109 ; 
   reg __422109_422109;
   reg _422110_422110 ; 
   reg __422110_422110;
   reg _422111_422111 ; 
   reg __422111_422111;
   reg _422112_422112 ; 
   reg __422112_422112;
   reg _422113_422113 ; 
   reg __422113_422113;
   reg _422114_422114 ; 
   reg __422114_422114;
   reg _422115_422115 ; 
   reg __422115_422115;
   reg _422116_422116 ; 
   reg __422116_422116;
   reg _422117_422117 ; 
   reg __422117_422117;
   reg _422118_422118 ; 
   reg __422118_422118;
   reg _422119_422119 ; 
   reg __422119_422119;
   reg _422120_422120 ; 
   reg __422120_422120;
   reg _422121_422121 ; 
   reg __422121_422121;
   reg _422122_422122 ; 
   reg __422122_422122;
   reg _422123_422123 ; 
   reg __422123_422123;
   reg _422124_422124 ; 
   reg __422124_422124;
   reg _422125_422125 ; 
   reg __422125_422125;
   reg _422126_422126 ; 
   reg __422126_422126;
   reg _422127_422127 ; 
   reg __422127_422127;
   reg _422128_422128 ; 
   reg __422128_422128;
   reg _422129_422129 ; 
   reg __422129_422129;
   reg _422130_422130 ; 
   reg __422130_422130;
   reg _422131_422131 ; 
   reg __422131_422131;
   reg _422132_422132 ; 
   reg __422132_422132;
   reg _422133_422133 ; 
   reg __422133_422133;
   reg _422134_422134 ; 
   reg __422134_422134;
   reg _422135_422135 ; 
   reg __422135_422135;
   reg _422136_422136 ; 
   reg __422136_422136;
   reg _422137_422137 ; 
   reg __422137_422137;
   reg _422138_422138 ; 
   reg __422138_422138;
   reg _422139_422139 ; 
   reg __422139_422139;
   reg _422140_422140 ; 
   reg __422140_422140;
   reg _422141_422141 ; 
   reg __422141_422141;
   reg _422142_422142 ; 
   reg __422142_422142;
   reg _422143_422143 ; 
   reg __422143_422143;
   reg _422144_422144 ; 
   reg __422144_422144;
   reg _422145_422145 ; 
   reg __422145_422145;
   reg _422146_422146 ; 
   reg __422146_422146;
   reg _422147_422147 ; 
   reg __422147_422147;
   reg _422148_422148 ; 
   reg __422148_422148;
   reg _422149_422149 ; 
   reg __422149_422149;
   reg _422150_422150 ; 
   reg __422150_422150;
   reg _422151_422151 ; 
   reg __422151_422151;
   reg _422152_422152 ; 
   reg __422152_422152;
   reg _422153_422153 ; 
   reg __422153_422153;
   reg _422154_422154 ; 
   reg __422154_422154;
   reg _422155_422155 ; 
   reg __422155_422155;
   reg _422156_422156 ; 
   reg __422156_422156;
   reg _422157_422157 ; 
   reg __422157_422157;
   reg _422158_422158 ; 
   reg __422158_422158;
   reg _422159_422159 ; 
   reg __422159_422159;
   reg _422160_422160 ; 
   reg __422160_422160;
   reg _422161_422161 ; 
   reg __422161_422161;
   reg _422162_422162 ; 
   reg __422162_422162;
   reg _422163_422163 ; 
   reg __422163_422163;
   reg _422164_422164 ; 
   reg __422164_422164;
   reg _422165_422165 ; 
   reg __422165_422165;
   reg _422166_422166 ; 
   reg __422166_422166;
   reg _422167_422167 ; 
   reg __422167_422167;
   reg _422168_422168 ; 
   reg __422168_422168;
   reg _422169_422169 ; 
   reg __422169_422169;
   reg _422170_422170 ; 
   reg __422170_422170;
   reg _422171_422171 ; 
   reg __422171_422171;
   reg _422172_422172 ; 
   reg __422172_422172;
   reg _422173_422173 ; 
   reg __422173_422173;
   reg _422174_422174 ; 
   reg __422174_422174;
   reg _422175_422175 ; 
   reg __422175_422175;
   reg _422176_422176 ; 
   reg __422176_422176;
   reg _422177_422177 ; 
   reg __422177_422177;
   reg _422178_422178 ; 
   reg __422178_422178;
   reg _422179_422179 ; 
   reg __422179_422179;
   reg _422180_422180 ; 
   reg __422180_422180;
   reg _422181_422181 ; 
   reg __422181_422181;
   reg _422182_422182 ; 
   reg __422182_422182;
   reg _422183_422183 ; 
   reg __422183_422183;
   reg _422184_422184 ; 
   reg __422184_422184;
   reg _422185_422185 ; 
   reg __422185_422185;
   reg _422186_422186 ; 
   reg __422186_422186;
   reg _422187_422187 ; 
   reg __422187_422187;
   reg _422188_422188 ; 
   reg __422188_422188;
   reg _422189_422189 ; 
   reg __422189_422189;
   reg _422190_422190 ; 
   reg __422190_422190;
   reg _422191_422191 ; 
   reg __422191_422191;
   reg _422192_422192 ; 
   reg __422192_422192;
   reg _422193_422193 ; 
   reg __422193_422193;
   reg _422194_422194 ; 
   reg __422194_422194;
   reg _422195_422195 ; 
   reg __422195_422195;
   reg _422196_422196 ; 
   reg __422196_422196;
   reg _422197_422197 ; 
   reg __422197_422197;
   reg _422198_422198 ; 
   reg __422198_422198;
   reg _422199_422199 ; 
   reg __422199_422199;
   reg _422200_422200 ; 
   reg __422200_422200;
   reg _422201_422201 ; 
   reg __422201_422201;
   reg _422202_422202 ; 
   reg __422202_422202;
   reg _422203_422203 ; 
   reg __422203_422203;
   reg _422204_422204 ; 
   reg __422204_422204;
   reg _422205_422205 ; 
   reg __422205_422205;
   reg _422206_422206 ; 
   reg __422206_422206;
   reg _422207_422207 ; 
   reg __422207_422207;
   reg _422208_422208 ; 
   reg __422208_422208;
   reg _422209_422209 ; 
   reg __422209_422209;
   reg _422210_422210 ; 
   reg __422210_422210;
   reg _422211_422211 ; 
   reg __422211_422211;
   reg _422212_422212 ; 
   reg __422212_422212;
   reg _422213_422213 ; 
   reg __422213_422213;
   reg _422214_422214 ; 
   reg __422214_422214;
   reg _422215_422215 ; 
   reg __422215_422215;
   reg _422216_422216 ; 
   reg __422216_422216;
   reg _422217_422217 ; 
   reg __422217_422217;
   reg _422218_422218 ; 
   reg __422218_422218;
   reg _422219_422219 ; 
   reg __422219_422219;
   reg _422220_422220 ; 
   reg __422220_422220;
   reg _422221_422221 ; 
   reg __422221_422221;
   reg _422222_422222 ; 
   reg __422222_422222;
   reg _422223_422223 ; 
   reg __422223_422223;
   reg _422224_422224 ; 
   reg __422224_422224;
   reg _422225_422225 ; 
   reg __422225_422225;
   reg _422226_422226 ; 
   reg __422226_422226;
   reg _422227_422227 ; 
   reg __422227_422227;
   reg _422228_422228 ; 
   reg __422228_422228;
   reg _422229_422229 ; 
   reg __422229_422229;
   reg _422230_422230 ; 
   reg __422230_422230;
   reg _422231_422231 ; 
   reg __422231_422231;
   reg _422232_422232 ; 
   reg __422232_422232;
   reg _422233_422233 ; 
   reg __422233_422233;
   reg _422234_422234 ; 
   reg __422234_422234;
   reg _422235_422235 ; 
   reg __422235_422235;
   reg _422236_422236 ; 
   reg __422236_422236;
   reg _422237_422237 ; 
   reg __422237_422237;
   reg _422238_422238 ; 
   reg __422238_422238;
   reg _422239_422239 ; 
   reg __422239_422239;
   reg _422240_422240 ; 
   reg __422240_422240;
   reg _422241_422241 ; 
   reg __422241_422241;
   reg _422242_422242 ; 
   reg __422242_422242;
   reg _422243_422243 ; 
   reg __422243_422243;
   reg _422244_422244 ; 
   reg __422244_422244;
   reg _422245_422245 ; 
   reg __422245_422245;
   reg _422246_422246 ; 
   reg __422246_422246;
   reg _422247_422247 ; 
   reg __422247_422247;
   reg _422248_422248 ; 
   reg __422248_422248;
   reg _422249_422249 ; 
   reg __422249_422249;
   reg _422250_422250 ; 
   reg __422250_422250;
   reg _422251_422251 ; 
   reg __422251_422251;
   reg _422252_422252 ; 
   reg __422252_422252;
   reg _422253_422253 ; 
   reg __422253_422253;
   reg _422254_422254 ; 
   reg __422254_422254;
   reg _422255_422255 ; 
   reg __422255_422255;
   reg _422256_422256 ; 
   reg __422256_422256;
   reg _422257_422257 ; 
   reg __422257_422257;
   reg _422258_422258 ; 
   reg __422258_422258;
   reg _422259_422259 ; 
   reg __422259_422259;
   reg _422260_422260 ; 
   reg __422260_422260;
   reg _422261_422261 ; 
   reg __422261_422261;
   reg _422262_422262 ; 
   reg __422262_422262;
   reg _422263_422263 ; 
   reg __422263_422263;
   reg _422264_422264 ; 
   reg __422264_422264;
   reg _422265_422265 ; 
   reg __422265_422265;
   reg _422266_422266 ; 
   reg __422266_422266;
   reg _422267_422267 ; 
   reg __422267_422267;
   reg _422268_422268 ; 
   reg __422268_422268;
   reg _422269_422269 ; 
   reg __422269_422269;
   reg _422270_422270 ; 
   reg __422270_422270;
   reg _422271_422271 ; 
   reg __422271_422271;
   reg _422272_422272 ; 
   reg __422272_422272;
   reg _422273_422273 ; 
   reg __422273_422273;
   reg _422274_422274 ; 
   reg __422274_422274;
   reg _422275_422275 ; 
   reg __422275_422275;
   reg _422276_422276 ; 
   reg __422276_422276;
   reg _422277_422277 ; 
   reg __422277_422277;
   reg _422278_422278 ; 
   reg __422278_422278;
   reg _422279_422279 ; 
   reg __422279_422279;
   reg _422280_422280 ; 
   reg __422280_422280;
   reg _422281_422281 ; 
   reg __422281_422281;
   reg _422282_422282 ; 
   reg __422282_422282;
   reg _422283_422283 ; 
   reg __422283_422283;
   reg _422284_422284 ; 
   reg __422284_422284;
   reg _422285_422285 ; 
   reg __422285_422285;
   reg _422286_422286 ; 
   reg __422286_422286;
   reg _422287_422287 ; 
   reg __422287_422287;
   reg _422288_422288 ; 
   reg __422288_422288;
   reg _422289_422289 ; 
   reg __422289_422289;
   reg _422290_422290 ; 
   reg __422290_422290;
   reg _422291_422291 ; 
   reg __422291_422291;
   reg _422292_422292 ; 
   reg __422292_422292;
   reg _422293_422293 ; 
   reg __422293_422293;
   reg _422294_422294 ; 
   reg __422294_422294;
   reg _422295_422295 ; 
   reg __422295_422295;
   reg _422296_422296 ; 
   reg __422296_422296;
   reg _422297_422297 ; 
   reg __422297_422297;
   reg _422298_422298 ; 
   reg __422298_422298;
   reg _422299_422299 ; 
   reg __422299_422299;
   reg _422300_422300 ; 
   reg __422300_422300;
   reg _422301_422301 ; 
   reg __422301_422301;
   reg _422302_422302 ; 
   reg __422302_422302;
   reg _422303_422303 ; 
   reg __422303_422303;
   reg _422304_422304 ; 
   reg __422304_422304;
   reg _422305_422305 ; 
   reg __422305_422305;
   reg _422306_422306 ; 
   reg __422306_422306;
   reg _422307_422307 ; 
   reg __422307_422307;
   reg _422308_422308 ; 
   reg __422308_422308;
   reg _422309_422309 ; 
   reg __422309_422309;
   reg _422310_422310 ; 
   reg __422310_422310;
   reg _422311_422311 ; 
   reg __422311_422311;
   reg _422312_422312 ; 
   reg __422312_422312;
   reg _422313_422313 ; 
   reg __422313_422313;
   reg _422314_422314 ; 
   reg __422314_422314;
   reg _422315_422315 ; 
   reg __422315_422315;
   reg _422316_422316 ; 
   reg __422316_422316;
   reg _422317_422317 ; 
   reg __422317_422317;
   reg _422318_422318 ; 
   reg __422318_422318;
   reg _422319_422319 ; 
   reg __422319_422319;
   reg _422320_422320 ; 
   reg __422320_422320;
   reg _422321_422321 ; 
   reg __422321_422321;
   reg _422322_422322 ; 
   reg __422322_422322;
   reg _422323_422323 ; 
   reg __422323_422323;
   reg _422324_422324 ; 
   reg __422324_422324;
   reg _422325_422325 ; 
   reg __422325_422325;
   reg _422326_422326 ; 
   reg __422326_422326;
   reg _422327_422327 ; 
   reg __422327_422327;
   reg _422328_422328 ; 
   reg __422328_422328;
   reg _422329_422329 ; 
   reg __422329_422329;
   reg _422330_422330 ; 
   reg __422330_422330;
   reg _422331_422331 ; 
   reg __422331_422331;
   reg _422332_422332 ; 
   reg __422332_422332;
   reg _422333_422333 ; 
   reg __422333_422333;
   reg _422334_422334 ; 
   reg __422334_422334;
   reg _422335_422335 ; 
   reg __422335_422335;
   reg _422336_422336 ; 
   reg __422336_422336;
   reg _422337_422337 ; 
   reg __422337_422337;
   reg _422338_422338 ; 
   reg __422338_422338;
   reg _422339_422339 ; 
   reg __422339_422339;
   reg _422340_422340 ; 
   reg __422340_422340;
   reg _422341_422341 ; 
   reg __422341_422341;
   reg _422342_422342 ; 
   reg __422342_422342;
   reg _422343_422343 ; 
   reg __422343_422343;
   reg _422344_422344 ; 
   reg __422344_422344;
   reg _422345_422345 ; 
   reg __422345_422345;
   reg _422346_422346 ; 
   reg __422346_422346;
   reg _422347_422347 ; 
   reg __422347_422347;
   reg _422348_422348 ; 
   reg __422348_422348;
   reg _422349_422349 ; 
   reg __422349_422349;
   reg _422350_422350 ; 
   reg __422350_422350;
   reg _422351_422351 ; 
   reg __422351_422351;
   reg _422352_422352 ; 
   reg __422352_422352;
   reg _422353_422353 ; 
   reg __422353_422353;
   reg _422354_422354 ; 
   reg __422354_422354;
   reg _422355_422355 ; 
   reg __422355_422355;
   reg _422356_422356 ; 
   reg __422356_422356;
   reg _422357_422357 ; 
   reg __422357_422357;
   reg _422358_422358 ; 
   reg __422358_422358;
   reg _422359_422359 ; 
   reg __422359_422359;
   reg _422360_422360 ; 
   reg __422360_422360;
   reg _422361_422361 ; 
   reg __422361_422361;
   reg _422362_422362 ; 
   reg __422362_422362;
   reg _422363_422363 ; 
   reg __422363_422363;
   reg _422364_422364 ; 
   reg __422364_422364;
   reg _422365_422365 ; 
   reg __422365_422365;
   reg _422366_422366 ; 
   reg __422366_422366;
   reg _422367_422367 ; 
   reg __422367_422367;
   reg _422368_422368 ; 
   reg __422368_422368;
   reg _422369_422369 ; 
   reg __422369_422369;
   reg _422370_422370 ; 
   reg __422370_422370;
   reg _422371_422371 ; 
   reg __422371_422371;
   reg _422372_422372 ; 
   reg __422372_422372;
   reg _422373_422373 ; 
   reg __422373_422373;
   reg _422374_422374 ; 
   reg __422374_422374;
   reg _422375_422375 ; 
   reg __422375_422375;
   reg _422376_422376 ; 
   reg __422376_422376;
   reg _422377_422377 ; 
   reg __422377_422377;
   reg _422378_422378 ; 
   reg __422378_422378;
   reg _422379_422379 ; 
   reg __422379_422379;
   reg _422380_422380 ; 
   reg __422380_422380;
   reg _422381_422381 ; 
   reg __422381_422381;
   reg _422382_422382 ; 
   reg __422382_422382;
   reg _422383_422383 ; 
   reg __422383_422383;
   reg _422384_422384 ; 
   reg __422384_422384;
   reg _422385_422385 ; 
   reg __422385_422385;
   reg _422386_422386 ; 
   reg __422386_422386;
   reg _422387_422387 ; 
   reg __422387_422387;
   reg _422388_422388 ; 
   reg __422388_422388;
   reg _422389_422389 ; 
   reg __422389_422389;
   reg _422390_422390 ; 
   reg __422390_422390;
   reg _422391_422391 ; 
   reg __422391_422391;
   reg _422392_422392 ; 
   reg __422392_422392;
   reg _422393_422393 ; 
   reg __422393_422393;
   reg _422394_422394 ; 
   reg __422394_422394;
   reg _422395_422395 ; 
   reg __422395_422395;
   reg _422396_422396 ; 
   reg __422396_422396;
   reg _422397_422397 ; 
   reg __422397_422397;
   reg _422398_422398 ; 
   reg __422398_422398;
   reg _422399_422399 ; 
   reg __422399_422399;
   reg _422400_422400 ; 
   reg __422400_422400;
   reg _422401_422401 ; 
   reg __422401_422401;
   reg _422402_422402 ; 
   reg __422402_422402;
   reg _422403_422403 ; 
   reg __422403_422403;
   reg _422404_422404 ; 
   reg __422404_422404;
   reg _422405_422405 ; 
   reg __422405_422405;
   reg _422406_422406 ; 
   reg __422406_422406;
   reg _422407_422407 ; 
   reg __422407_422407;
   reg _422408_422408 ; 
   reg __422408_422408;
   reg _422409_422409 ; 
   reg __422409_422409;
   reg _422410_422410 ; 
   reg __422410_422410;
   reg _422411_422411 ; 
   reg __422411_422411;
   reg _422412_422412 ; 
   reg __422412_422412;
   reg _422413_422413 ; 
   reg __422413_422413;
   reg _422414_422414 ; 
   reg __422414_422414;
   reg _422415_422415 ; 
   reg __422415_422415;
   reg _422416_422416 ; 
   reg __422416_422416;
   reg _422417_422417 ; 
   reg __422417_422417;
   reg _422418_422418 ; 
   reg __422418_422418;
   reg _422419_422419 ; 
   reg __422419_422419;
   reg _422420_422420 ; 
   reg __422420_422420;
   reg _422421_422421 ; 
   reg __422421_422421;
   reg _422422_422422 ; 
   reg __422422_422422;
   reg _422423_422423 ; 
   reg __422423_422423;
   reg _422424_422424 ; 
   reg __422424_422424;
   reg _422425_422425 ; 
   reg __422425_422425;
   reg _422426_422426 ; 
   reg __422426_422426;
   reg _422427_422427 ; 
   reg __422427_422427;
   reg _422428_422428 ; 
   reg __422428_422428;
   reg _422429_422429 ; 
   reg __422429_422429;
   reg _422430_422430 ; 
   reg __422430_422430;
   reg _422431_422431 ; 
   reg __422431_422431;
   reg _422432_422432 ; 
   reg __422432_422432;
   reg _422433_422433 ; 
   reg __422433_422433;
   reg _422434_422434 ; 
   reg __422434_422434;
   reg _422435_422435 ; 
   reg __422435_422435;
   reg _422436_422436 ; 
   reg __422436_422436;
   reg _422437_422437 ; 
   reg __422437_422437;
   reg _422438_422438 ; 
   reg __422438_422438;
   reg _422439_422439 ; 
   reg __422439_422439;
   reg _422440_422440 ; 
   reg __422440_422440;
   reg _422441_422441 ; 
   reg __422441_422441;
   reg _422442_422442 ; 
   reg __422442_422442;
   reg _422443_422443 ; 
   reg __422443_422443;
   reg _422444_422444 ; 
   reg __422444_422444;
   reg _422445_422445 ; 
   reg __422445_422445;
   reg _422446_422446 ; 
   reg __422446_422446;
   reg _422447_422447 ; 
   reg __422447_422447;
   reg _422448_422448 ; 
   reg __422448_422448;
   reg _422449_422449 ; 
   reg __422449_422449;
   reg _422450_422450 ; 
   reg __422450_422450;
   reg _422451_422451 ; 
   reg __422451_422451;
   reg _422452_422452 ; 
   reg __422452_422452;
   reg _422453_422453 ; 
   reg __422453_422453;
   reg _422454_422454 ; 
   reg __422454_422454;
   reg _422455_422455 ; 
   reg __422455_422455;
   reg _422456_422456 ; 
   reg __422456_422456;
   reg _422457_422457 ; 
   reg __422457_422457;
   reg _422458_422458 ; 
   reg __422458_422458;
   reg _422459_422459 ; 
   reg __422459_422459;
   reg _422460_422460 ; 
   reg __422460_422460;
   reg _422461_422461 ; 
   reg __422461_422461;
   reg _422462_422462 ; 
   reg __422462_422462;
   reg _422463_422463 ; 
   reg __422463_422463;
   reg _422464_422464 ; 
   reg __422464_422464;
   reg _422465_422465 ; 
   reg __422465_422465;
   reg _422466_422466 ; 
   reg __422466_422466;
   reg _422467_422467 ; 
   reg __422467_422467;
   reg _422468_422468 ; 
   reg __422468_422468;
   reg _422469_422469 ; 
   reg __422469_422469;
   reg _422470_422470 ; 
   reg __422470_422470;
   reg _422471_422471 ; 
   reg __422471_422471;
   reg _422472_422472 ; 
   reg __422472_422472;
   reg _422473_422473 ; 
   reg __422473_422473;
   reg _422474_422474 ; 
   reg __422474_422474;
   reg _422475_422475 ; 
   reg __422475_422475;
   reg _422476_422476 ; 
   reg __422476_422476;
   reg _422477_422477 ; 
   reg __422477_422477;
   reg _422478_422478 ; 
   reg __422478_422478;
   reg _422479_422479 ; 
   reg __422479_422479;
   reg _422480_422480 ; 
   reg __422480_422480;
   reg _422481_422481 ; 
   reg __422481_422481;
   reg _422482_422482 ; 
   reg __422482_422482;
   reg _422483_422483 ; 
   reg __422483_422483;
   reg _422484_422484 ; 
   reg __422484_422484;
   reg _422485_422485 ; 
   reg __422485_422485;
   reg _422486_422486 ; 
   reg __422486_422486;
   reg _422487_422487 ; 
   reg __422487_422487;
   reg _422488_422488 ; 
   reg __422488_422488;
   reg _422489_422489 ; 
   reg __422489_422489;
   reg _422490_422490 ; 
   reg __422490_422490;
   reg _422491_422491 ; 
   reg __422491_422491;
   reg _422492_422492 ; 
   reg __422492_422492;
   reg _422493_422493 ; 
   reg __422493_422493;
   reg _422494_422494 ; 
   reg __422494_422494;
   reg _422495_422495 ; 
   reg __422495_422495;
   reg _422496_422496 ; 
   reg __422496_422496;
   reg _422497_422497 ; 
   reg __422497_422497;
   reg _422498_422498 ; 
   reg __422498_422498;
   reg _422499_422499 ; 
   reg __422499_422499;
   reg _422500_422500 ; 
   reg __422500_422500;
   reg _422501_422501 ; 
   reg __422501_422501;
   reg _422502_422502 ; 
   reg __422502_422502;
   reg _422503_422503 ; 
   reg __422503_422503;
   reg _422504_422504 ; 
   reg __422504_422504;
   reg _422505_422505 ; 
   reg __422505_422505;
   reg _422506_422506 ; 
   reg __422506_422506;
   reg _422507_422507 ; 
   reg __422507_422507;
   reg _422508_422508 ; 
   reg __422508_422508;
   reg _422509_422509 ; 
   reg __422509_422509;
   reg _422510_422510 ; 
   reg __422510_422510;
   reg _422511_422511 ; 
   reg __422511_422511;
   reg _422512_422512 ; 
   reg __422512_422512;
   reg _422513_422513 ; 
   reg __422513_422513;
   reg _422514_422514 ; 
   reg __422514_422514;
   reg _422515_422515 ; 
   reg __422515_422515;
   reg _422516_422516 ; 
   reg __422516_422516;
   reg _422517_422517 ; 
   reg __422517_422517;
   reg _422518_422518 ; 
   reg __422518_422518;
   reg _422519_422519 ; 
   reg __422519_422519;
   reg _422520_422520 ; 
   reg __422520_422520;
   reg _422521_422521 ; 
   reg __422521_422521;
   reg _422522_422522 ; 
   reg __422522_422522;
   reg _422523_422523 ; 
   reg __422523_422523;
   reg _422524_422524 ; 
   reg __422524_422524;
   reg _422525_422525 ; 
   reg __422525_422525;
   reg _422526_422526 ; 
   reg __422526_422526;
   reg _422527_422527 ; 
   reg __422527_422527;
   reg _422528_422528 ; 
   reg __422528_422528;
   reg _422529_422529 ; 
   reg __422529_422529;
   reg _422530_422530 ; 
   reg __422530_422530;
   reg _422531_422531 ; 
   reg __422531_422531;
   reg _422532_422532 ; 
   reg __422532_422532;
   reg _422533_422533 ; 
   reg __422533_422533;
   reg _422534_422534 ; 
   reg __422534_422534;
   reg _422535_422535 ; 
   reg __422535_422535;
   reg _422536_422536 ; 
   reg __422536_422536;
   reg _422537_422537 ; 
   reg __422537_422537;
   reg _422538_422538 ; 
   reg __422538_422538;
   reg _422539_422539 ; 
   reg __422539_422539;
   reg _422540_422540 ; 
   reg __422540_422540;
   reg _422541_422541 ; 
   reg __422541_422541;
   reg _422542_422542 ; 
   reg __422542_422542;
   reg _422543_422543 ; 
   reg __422543_422543;
   reg _422544_422544 ; 
   reg __422544_422544;
   reg _422545_422545 ; 
   reg __422545_422545;
   reg _422546_422546 ; 
   reg __422546_422546;
   reg _422547_422547 ; 
   reg __422547_422547;
   reg _422548_422548 ; 
   reg __422548_422548;
   reg _422549_422549 ; 
   reg __422549_422549;
   reg _422550_422550 ; 
   reg __422550_422550;
   reg _422551_422551 ; 
   reg __422551_422551;
   reg _422552_422552 ; 
   reg __422552_422552;
   reg _422553_422553 ; 
   reg __422553_422553;
   reg _422554_422554 ; 
   reg __422554_422554;
   reg _422555_422555 ; 
   reg __422555_422555;
   reg _422556_422556 ; 
   reg __422556_422556;
   reg _422557_422557 ; 
   reg __422557_422557;
   reg _422558_422558 ; 
   reg __422558_422558;
   reg _422559_422559 ; 
   reg __422559_422559;
   reg _422560_422560 ; 
   reg __422560_422560;
   reg _422561_422561 ; 
   reg __422561_422561;
   reg _422562_422562 ; 
   reg __422562_422562;
   reg _422563_422563 ; 
   reg __422563_422563;
   reg _422564_422564 ; 
   reg __422564_422564;
   reg _422565_422565 ; 
   reg __422565_422565;
   reg _422566_422566 ; 
   reg __422566_422566;
   reg _422567_422567 ; 
   reg __422567_422567;
   reg _422568_422568 ; 
   reg __422568_422568;
   reg _422569_422569 ; 
   reg __422569_422569;
   reg _422570_422570 ; 
   reg __422570_422570;
   reg _422571_422571 ; 
   reg __422571_422571;
   reg _422572_422572 ; 
   reg __422572_422572;
   reg _422573_422573 ; 
   reg __422573_422573;
   reg _422574_422574 ; 
   reg __422574_422574;
   reg _422575_422575 ; 
   reg __422575_422575;
   reg _422576_422576 ; 
   reg __422576_422576;
   reg _422577_422577 ; 
   reg __422577_422577;
   reg _422578_422578 ; 
   reg __422578_422578;
   reg _422579_422579 ; 
   reg __422579_422579;
   reg _422580_422580 ; 
   reg __422580_422580;
   reg _422581_422581 ; 
   reg __422581_422581;
   reg _422582_422582 ; 
   reg __422582_422582;
   reg _422583_422583 ; 
   reg __422583_422583;
   reg _422584_422584 ; 
   reg __422584_422584;
   reg _422585_422585 ; 
   reg __422585_422585;
   reg _422586_422586 ; 
   reg __422586_422586;
   reg _422587_422587 ; 
   reg __422587_422587;
   reg _422588_422588 ; 
   reg __422588_422588;
   reg _422589_422589 ; 
   reg __422589_422589;
   reg _422590_422590 ; 
   reg __422590_422590;
   reg _422591_422591 ; 
   reg __422591_422591;
   reg _422592_422592 ; 
   reg __422592_422592;
   reg _422593_422593 ; 
   reg __422593_422593;
   reg _422594_422594 ; 
   reg __422594_422594;
   reg _422595_422595 ; 
   reg __422595_422595;
   reg _422596_422596 ; 
   reg __422596_422596;
   reg _422597_422597 ; 
   reg __422597_422597;
   reg _422598_422598 ; 
   reg __422598_422598;
   reg _422599_422599 ; 
   reg __422599_422599;
   reg _422600_422600 ; 
   reg __422600_422600;
   reg _422601_422601 ; 
   reg __422601_422601;
   reg _422602_422602 ; 
   reg __422602_422602;
   reg _422603_422603 ; 
   reg __422603_422603;
   reg _422604_422604 ; 
   reg __422604_422604;
   reg _422605_422605 ; 
   reg __422605_422605;
   reg _422606_422606 ; 
   reg __422606_422606;
   reg _422607_422607 ; 
   reg __422607_422607;
   reg _422608_422608 ; 
   reg __422608_422608;
   reg _422609_422609 ; 
   reg __422609_422609;
   reg _422610_422610 ; 
   reg __422610_422610;
   reg _422611_422611 ; 
   reg __422611_422611;
   reg _422612_422612 ; 
   reg __422612_422612;
   reg _422613_422613 ; 
   reg __422613_422613;
   reg _422614_422614 ; 
   reg __422614_422614;
   reg _422615_422615 ; 
   reg __422615_422615;
   reg _422616_422616 ; 
   reg __422616_422616;
   reg _422617_422617 ; 
   reg __422617_422617;
   reg _422618_422618 ; 
   reg __422618_422618;
   reg _422619_422619 ; 
   reg __422619_422619;
   reg _422620_422620 ; 
   reg __422620_422620;
   reg _422621_422621 ; 
   reg __422621_422621;
   reg _422622_422622 ; 
   reg __422622_422622;
   reg _422623_422623 ; 
   reg __422623_422623;
   reg _422624_422624 ; 
   reg __422624_422624;
   reg _422625_422625 ; 
   reg __422625_422625;
   reg _422626_422626 ; 
   reg __422626_422626;
   reg _422627_422627 ; 
   reg __422627_422627;
   reg _422628_422628 ; 
   reg __422628_422628;
   reg _422629_422629 ; 
   reg __422629_422629;
   reg _422630_422630 ; 
   reg __422630_422630;
   reg _422631_422631 ; 
   reg __422631_422631;
   reg _422632_422632 ; 
   reg __422632_422632;
   reg _422633_422633 ; 
   reg __422633_422633;
   reg _422634_422634 ; 
   reg __422634_422634;
   reg _422635_422635 ; 
   reg __422635_422635;
   reg _422636_422636 ; 
   reg __422636_422636;
   reg _422637_422637 ; 
   reg __422637_422637;
   reg _422638_422638 ; 
   reg __422638_422638;
   reg _422639_422639 ; 
   reg __422639_422639;
   reg _422640_422640 ; 
   reg __422640_422640;
   reg _422641_422641 ; 
   reg __422641_422641;
   reg _422642_422642 ; 
   reg __422642_422642;
   reg _422643_422643 ; 
   reg __422643_422643;
   reg _422644_422644 ; 
   reg __422644_422644;
   reg _422645_422645 ; 
   reg __422645_422645;
   reg _422646_422646 ; 
   reg __422646_422646;
   reg _422647_422647 ; 
   reg __422647_422647;
   reg _422648_422648 ; 
   reg __422648_422648;
   reg _422649_422649 ; 
   reg __422649_422649;
   reg _422650_422650 ; 
   reg __422650_422650;
   reg _422651_422651 ; 
   reg __422651_422651;
   reg _422652_422652 ; 
   reg __422652_422652;
   reg _422653_422653 ; 
   reg __422653_422653;
   reg _422654_422654 ; 
   reg __422654_422654;
   reg _422655_422655 ; 
   reg __422655_422655;
   reg _422656_422656 ; 
   reg __422656_422656;
   reg _422657_422657 ; 
   reg __422657_422657;
   reg _422658_422658 ; 
   reg __422658_422658;
   reg _422659_422659 ; 
   reg __422659_422659;
   reg _422660_422660 ; 
   reg __422660_422660;
   reg _422661_422661 ; 
   reg __422661_422661;
   reg _422662_422662 ; 
   reg __422662_422662;
   reg _422663_422663 ; 
   reg __422663_422663;
   reg _422664_422664 ; 
   reg __422664_422664;
   reg _422665_422665 ; 
   reg __422665_422665;
   reg _422666_422666 ; 
   reg __422666_422666;
   reg _422667_422667 ; 
   reg __422667_422667;
   reg _422668_422668 ; 
   reg __422668_422668;
   reg _422669_422669 ; 
   reg __422669_422669;
   reg _422670_422670 ; 
   reg __422670_422670;
   reg _422671_422671 ; 
   reg __422671_422671;
   reg _422672_422672 ; 
   reg __422672_422672;
   reg _422673_422673 ; 
   reg __422673_422673;
   reg _422674_422674 ; 
   reg __422674_422674;
   reg _422675_422675 ; 
   reg __422675_422675;
   reg _422676_422676 ; 
   reg __422676_422676;
   reg _422677_422677 ; 
   reg __422677_422677;
   reg _422678_422678 ; 
   reg __422678_422678;
   reg _422679_422679 ; 
   reg __422679_422679;
   reg _422680_422680 ; 
   reg __422680_422680;
   reg _422681_422681 ; 
   reg __422681_422681;
   reg _422682_422682 ; 
   reg __422682_422682;
   reg _422683_422683 ; 
   reg __422683_422683;
   reg _422684_422684 ; 
   reg __422684_422684;
   reg _422685_422685 ; 
   reg __422685_422685;
   reg _422686_422686 ; 
   reg __422686_422686;
   reg _422687_422687 ; 
   reg __422687_422687;
   reg _422688_422688 ; 
   reg __422688_422688;
   reg _422689_422689 ; 
   reg __422689_422689;
   reg _422690_422690 ; 
   reg __422690_422690;
   reg _422691_422691 ; 
   reg __422691_422691;
   reg _422692_422692 ; 
   reg __422692_422692;
   reg _422693_422693 ; 
   reg __422693_422693;
   reg _422694_422694 ; 
   reg __422694_422694;
   reg _422695_422695 ; 
   reg __422695_422695;
   reg _422696_422696 ; 
   reg __422696_422696;
   reg _422697_422697 ; 
   reg __422697_422697;
   reg _422698_422698 ; 
   reg __422698_422698;
   reg _422699_422699 ; 
   reg __422699_422699;
   reg _422700_422700 ; 
   reg __422700_422700;
   reg _422701_422701 ; 
   reg __422701_422701;
   reg _422702_422702 ; 
   reg __422702_422702;
   reg _422703_422703 ; 
   reg __422703_422703;
   reg _422704_422704 ; 
   reg __422704_422704;
   reg _422705_422705 ; 
   reg __422705_422705;
   reg _422706_422706 ; 
   reg __422706_422706;
   reg _422707_422707 ; 
   reg __422707_422707;
   reg _422708_422708 ; 
   reg __422708_422708;
   reg _422709_422709 ; 
   reg __422709_422709;
   reg _422710_422710 ; 
   reg __422710_422710;
   reg _422711_422711 ; 
   reg __422711_422711;
   reg _422712_422712 ; 
   reg __422712_422712;
   reg _422713_422713 ; 
   reg __422713_422713;
   reg _422714_422714 ; 
   reg __422714_422714;
   reg _422715_422715 ; 
   reg __422715_422715;
   reg _422716_422716 ; 
   reg __422716_422716;
   reg _422717_422717 ; 
   reg __422717_422717;
   reg _422718_422718 ; 
   reg __422718_422718;
   reg _422719_422719 ; 
   reg __422719_422719;
   reg _422720_422720 ; 
   reg __422720_422720;
   reg _422721_422721 ; 
   reg __422721_422721;
   reg _422722_422722 ; 
   reg __422722_422722;
   reg _422723_422723 ; 
   reg __422723_422723;
   reg _422724_422724 ; 
   reg __422724_422724;
   reg _422725_422725 ; 
   reg __422725_422725;
   reg _422726_422726 ; 
   reg __422726_422726;
   reg _422727_422727 ; 
   reg __422727_422727;
   reg _422728_422728 ; 
   reg __422728_422728;
   reg _422729_422729 ; 
   reg __422729_422729;
   reg _422730_422730 ; 
   reg __422730_422730;
   reg _422731_422731 ; 
   reg __422731_422731;
   reg _422732_422732 ; 
   reg __422732_422732;
   reg _422733_422733 ; 
   reg __422733_422733;
   reg _422734_422734 ; 
   reg __422734_422734;
   reg _422735_422735 ; 
   reg __422735_422735;
   reg _422736_422736 ; 
   reg __422736_422736;
   reg _422737_422737 ; 
   reg __422737_422737;
   reg _422738_422738 ; 
   reg __422738_422738;
   reg _422739_422739 ; 
   reg __422739_422739;
   reg _422740_422740 ; 
   reg __422740_422740;
   reg _422741_422741 ; 
   reg __422741_422741;
   reg _422742_422742 ; 
   reg __422742_422742;
   reg _422743_422743 ; 
   reg __422743_422743;
   reg _422744_422744 ; 
   reg __422744_422744;
   reg _422745_422745 ; 
   reg __422745_422745;
   reg _422746_422746 ; 
   reg __422746_422746;
   reg _422747_422747 ; 
   reg __422747_422747;
   reg _422748_422748 ; 
   reg __422748_422748;
   reg _422749_422749 ; 
   reg __422749_422749;
   reg _422750_422750 ; 
   reg __422750_422750;
   reg _422751_422751 ; 
   reg __422751_422751;
   reg _422752_422752 ; 
   reg __422752_422752;
   reg _422753_422753 ; 
   reg __422753_422753;
   reg _422754_422754 ; 
   reg __422754_422754;
   reg _422755_422755 ; 
   reg __422755_422755;
   reg _422756_422756 ; 
   reg __422756_422756;
   reg _422757_422757 ; 
   reg __422757_422757;
   reg _422758_422758 ; 
   reg __422758_422758;
   reg _422759_422759 ; 
   reg __422759_422759;
   reg _422760_422760 ; 
   reg __422760_422760;
   reg _422761_422761 ; 
   reg __422761_422761;
   reg _422762_422762 ; 
   reg __422762_422762;
   reg _422763_422763 ; 
   reg __422763_422763;
   reg _422764_422764 ; 
   reg __422764_422764;
   reg _422765_422765 ; 
   reg __422765_422765;
   reg _422766_422766 ; 
   reg __422766_422766;
   reg _422767_422767 ; 
   reg __422767_422767;
   reg _422768_422768 ; 
   reg __422768_422768;
   reg _422769_422769 ; 
   reg __422769_422769;
   reg _422770_422770 ; 
   reg __422770_422770;
   reg _422771_422771 ; 
   reg __422771_422771;
   reg _422772_422772 ; 
   reg __422772_422772;
   reg _422773_422773 ; 
   reg __422773_422773;
   reg _422774_422774 ; 
   reg __422774_422774;
   reg _422775_422775 ; 
   reg __422775_422775;
   reg _422776_422776 ; 
   reg __422776_422776;
   reg _422777_422777 ; 
   reg __422777_422777;
   reg _422778_422778 ; 
   reg __422778_422778;
   reg _422779_422779 ; 
   reg __422779_422779;
   reg _422780_422780 ; 
   reg __422780_422780;
   reg _422781_422781 ; 
   reg __422781_422781;
   reg _422782_422782 ; 
   reg __422782_422782;
   reg _422783_422783 ; 
   reg __422783_422783;
   reg _422784_422784 ; 
   reg __422784_422784;
   reg _422785_422785 ; 
   reg __422785_422785;
   reg _422786_422786 ; 
   reg __422786_422786;
   reg _422787_422787 ; 
   reg __422787_422787;
   reg _422788_422788 ; 
   reg __422788_422788;
   reg _422789_422789 ; 
   reg __422789_422789;
   reg _422790_422790 ; 
   reg __422790_422790;
   reg _422791_422791 ; 
   reg __422791_422791;
   reg _422792_422792 ; 
   reg __422792_422792;
   reg _422793_422793 ; 
   reg __422793_422793;
   reg _422794_422794 ; 
   reg __422794_422794;
   reg _422795_422795 ; 
   reg __422795_422795;
   reg _422796_422796 ; 
   reg __422796_422796;
   reg _422797_422797 ; 
   reg __422797_422797;
   reg _422798_422798 ; 
   reg __422798_422798;
   reg _422799_422799 ; 
   reg __422799_422799;
   reg _422800_422800 ; 
   reg __422800_422800;
   reg _422801_422801 ; 
   reg __422801_422801;
   reg _422802_422802 ; 
   reg __422802_422802;
   reg _422803_422803 ; 
   reg __422803_422803;
   reg _422804_422804 ; 
   reg __422804_422804;
   reg _422805_422805 ; 
   reg __422805_422805;
   reg _422806_422806 ; 
   reg __422806_422806;
   reg _422807_422807 ; 
   reg __422807_422807;
   reg _422808_422808 ; 
   reg __422808_422808;
   reg _422809_422809 ; 
   reg __422809_422809;
   reg _422810_422810 ; 
   reg __422810_422810;
   reg _422811_422811 ; 
   reg __422811_422811;
   reg _422812_422812 ; 
   reg __422812_422812;
   reg _422813_422813 ; 
   reg __422813_422813;
   reg _422814_422814 ; 
   reg __422814_422814;
   reg _422815_422815 ; 
   reg __422815_422815;
   reg _422816_422816 ; 
   reg __422816_422816;
   reg _422817_422817 ; 
   reg __422817_422817;
   reg _422818_422818 ; 
   reg __422818_422818;
   reg _422819_422819 ; 
   reg __422819_422819;
   reg _422820_422820 ; 
   reg __422820_422820;
   reg _422821_422821 ; 
   reg __422821_422821;
   reg _422822_422822 ; 
   reg __422822_422822;
   reg _422823_422823 ; 
   reg __422823_422823;
   reg _422824_422824 ; 
   reg __422824_422824;
   reg _422825_422825 ; 
   reg __422825_422825;
   reg _422826_422826 ; 
   reg __422826_422826;
   reg _422827_422827 ; 
   reg __422827_422827;
   reg _422828_422828 ; 
   reg __422828_422828;
   reg _422829_422829 ; 
   reg __422829_422829;
   reg _422830_422830 ; 
   reg __422830_422830;
   reg _422831_422831 ; 
   reg __422831_422831;
   reg _422832_422832 ; 
   reg __422832_422832;
   reg _422833_422833 ; 
   reg __422833_422833;
   reg _422834_422834 ; 
   reg __422834_422834;
   reg _422835_422835 ; 
   reg __422835_422835;
   reg _422836_422836 ; 
   reg __422836_422836;
   reg _422837_422837 ; 
   reg __422837_422837;
   reg _422838_422838 ; 
   reg __422838_422838;
   reg _422839_422839 ; 
   reg __422839_422839;
   reg _422840_422840 ; 
   reg __422840_422840;
   reg _422841_422841 ; 
   reg __422841_422841;
   reg _422842_422842 ; 
   reg __422842_422842;
   reg _422843_422843 ; 
   reg __422843_422843;
   reg _422844_422844 ; 
   reg __422844_422844;
   reg _422845_422845 ; 
   reg __422845_422845;
   reg _422846_422846 ; 
   reg __422846_422846;
   reg _422847_422847 ; 
   reg __422847_422847;
   reg _422848_422848 ; 
   reg __422848_422848;
   reg _422849_422849 ; 
   reg __422849_422849;
   reg _422850_422850 ; 
   reg __422850_422850;
   reg _422851_422851 ; 
   reg __422851_422851;
   reg _422852_422852 ; 
   reg __422852_422852;
   reg _422853_422853 ; 
   reg __422853_422853;
   reg _422854_422854 ; 
   reg __422854_422854;
   reg _422855_422855 ; 
   reg __422855_422855;
   reg _422856_422856 ; 
   reg __422856_422856;
   reg _422857_422857 ; 
   reg __422857_422857;
   reg _422858_422858 ; 
   reg __422858_422858;
   reg _422859_422859 ; 
   reg __422859_422859;
   reg _422860_422860 ; 
   reg __422860_422860;
   reg _422861_422861 ; 
   reg __422861_422861;
   reg _422862_422862 ; 
   reg __422862_422862;
   reg _422863_422863 ; 
   reg __422863_422863;
   reg _422864_422864 ; 
   reg __422864_422864;
   reg _422865_422865 ; 
   reg __422865_422865;
   reg _422866_422866 ; 
   reg __422866_422866;
   reg _422867_422867 ; 
   reg __422867_422867;
   reg _422868_422868 ; 
   reg __422868_422868;
   reg _422869_422869 ; 
   reg __422869_422869;
   reg _422870_422870 ; 
   reg __422870_422870;
   reg _422871_422871 ; 
   reg __422871_422871;
   reg _422872_422872 ; 
   reg __422872_422872;
   reg _422873_422873 ; 
   reg __422873_422873;
   reg _422874_422874 ; 
   reg __422874_422874;
   reg _422875_422875 ; 
   reg __422875_422875;
   reg _422876_422876 ; 
   reg __422876_422876;
   reg _422877_422877 ; 
   reg __422877_422877;
   reg _422878_422878 ; 
   reg __422878_422878;
   reg _422879_422879 ; 
   reg __422879_422879;
   reg _422880_422880 ; 
   reg __422880_422880;
   reg _422881_422881 ; 
   reg __422881_422881;
   reg _422882_422882 ; 
   reg __422882_422882;
   reg _422883_422883 ; 
   reg __422883_422883;
   reg _422884_422884 ; 
   reg __422884_422884;
   reg _422885_422885 ; 
   reg __422885_422885;
   reg _422886_422886 ; 
   reg __422886_422886;
   reg _422887_422887 ; 
   reg __422887_422887;
   reg _422888_422888 ; 
   reg __422888_422888;
   reg _422889_422889 ; 
   reg __422889_422889;
   reg _422890_422890 ; 
   reg __422890_422890;
   reg _422891_422891 ; 
   reg __422891_422891;
   reg _422892_422892 ; 
   reg __422892_422892;
   reg _422893_422893 ; 
   reg __422893_422893;
   reg _422894_422894 ; 
   reg __422894_422894;
   reg _422895_422895 ; 
   reg __422895_422895;
   reg _422896_422896 ; 
   reg __422896_422896;
   reg _422897_422897 ; 
   reg __422897_422897;
   reg _422898_422898 ; 
   reg __422898_422898;
   reg _422899_422899 ; 
   reg __422899_422899;
   reg _422900_422900 ; 
   reg __422900_422900;
   reg _422901_422901 ; 
   reg __422901_422901;
   reg _422902_422902 ; 
   reg __422902_422902;
   reg _422903_422903 ; 
   reg __422903_422903;
   reg _422904_422904 ; 
   reg __422904_422904;
   reg _422905_422905 ; 
   reg __422905_422905;
   reg _422906_422906 ; 
   reg __422906_422906;
   reg _422907_422907 ; 
   reg __422907_422907;
   reg _422908_422908 ; 
   reg __422908_422908;
   reg _422909_422909 ; 
   reg __422909_422909;
   reg _422910_422910 ; 
   reg __422910_422910;
   reg _422911_422911 ; 
   reg __422911_422911;
   reg _422912_422912 ; 
   reg __422912_422912;
   reg _422913_422913 ; 
   reg __422913_422913;
   reg _422914_422914 ; 
   reg __422914_422914;
   reg _422915_422915 ; 
   reg __422915_422915;
   reg _422916_422916 ; 
   reg __422916_422916;
   reg _422917_422917 ; 
   reg __422917_422917;
   reg _422918_422918 ; 
   reg __422918_422918;
   reg _422919_422919 ; 
   reg __422919_422919;
   reg _422920_422920 ; 
   reg __422920_422920;
   reg _422921_422921 ; 
   reg __422921_422921;
   reg _422922_422922 ; 
   reg __422922_422922;
   reg _422923_422923 ; 
   reg __422923_422923;
   reg _422924_422924 ; 
   reg __422924_422924;
   reg _422925_422925 ; 
   reg __422925_422925;
   reg _422926_422926 ; 
   reg __422926_422926;
   reg _422927_422927 ; 
   reg __422927_422927;
   reg _422928_422928 ; 
   reg __422928_422928;
   reg _422929_422929 ; 
   reg __422929_422929;
   reg _422930_422930 ; 
   reg __422930_422930;
   reg _422931_422931 ; 
   reg __422931_422931;
   reg _422932_422932 ; 
   reg __422932_422932;
   reg _422933_422933 ; 
   reg __422933_422933;
   reg _422934_422934 ; 
   reg __422934_422934;
   reg _422935_422935 ; 
   reg __422935_422935;
   reg _422936_422936 ; 
   reg __422936_422936;
   reg _422937_422937 ; 
   reg __422937_422937;
   reg _422938_422938 ; 
   reg __422938_422938;
   reg _422939_422939 ; 
   reg __422939_422939;
   reg _422940_422940 ; 
   reg __422940_422940;
   reg _422941_422941 ; 
   reg __422941_422941;
   reg _422942_422942 ; 
   reg __422942_422942;
   reg _422943_422943 ; 
   reg __422943_422943;
   reg _422944_422944 ; 
   reg __422944_422944;
   reg _422945_422945 ; 
   reg __422945_422945;
   reg _422946_422946 ; 
   reg __422946_422946;
   reg _422947_422947 ; 
   reg __422947_422947;
   reg _422948_422948 ; 
   reg __422948_422948;
   reg _422949_422949 ; 
   reg __422949_422949;
   reg _422950_422950 ; 
   reg __422950_422950;
   reg _422951_422951 ; 
   reg __422951_422951;
   reg _422952_422952 ; 
   reg __422952_422952;
   reg _422953_422953 ; 
   reg __422953_422953;
   reg _422954_422954 ; 
   reg __422954_422954;
   reg _422955_422955 ; 
   reg __422955_422955;
   reg _422956_422956 ; 
   reg __422956_422956;
   reg _422957_422957 ; 
   reg __422957_422957;
   reg _422958_422958 ; 
   reg __422958_422958;
   reg _422959_422959 ; 
   reg __422959_422959;
   reg _422960_422960 ; 
   reg __422960_422960;
   reg _422961_422961 ; 
   reg __422961_422961;
   reg _422962_422962 ; 
   reg __422962_422962;
   reg _422963_422963 ; 
   reg __422963_422963;
   reg _422964_422964 ; 
   reg __422964_422964;
   reg _422965_422965 ; 
   reg __422965_422965;
   reg _422966_422966 ; 
   reg __422966_422966;
   reg _422967_422967 ; 
   reg __422967_422967;
   reg _422968_422968 ; 
   reg __422968_422968;
   reg _422969_422969 ; 
   reg __422969_422969;
   reg _422970_422970 ; 
   reg __422970_422970;
   reg _422971_422971 ; 
   reg __422971_422971;
   reg _422972_422972 ; 
   reg __422972_422972;
   reg _422973_422973 ; 
   reg __422973_422973;
   reg _422974_422974 ; 
   reg __422974_422974;
   reg _422975_422975 ; 
   reg __422975_422975;
   reg _422976_422976 ; 
   reg __422976_422976;
   reg _422977_422977 ; 
   reg __422977_422977;
   reg _422978_422978 ; 
   reg __422978_422978;
   reg _422979_422979 ; 
   reg __422979_422979;
   reg _422980_422980 ; 
   reg __422980_422980;
   reg _422981_422981 ; 
   reg __422981_422981;
   reg _422982_422982 ; 
   reg __422982_422982;
   reg _422983_422983 ; 
   reg __422983_422983;
   reg _422984_422984 ; 
   reg __422984_422984;
   reg _422985_422985 ; 
   reg __422985_422985;
   reg _422986_422986 ; 
   reg __422986_422986;
   reg _422987_422987 ; 
   reg __422987_422987;
   reg _422988_422988 ; 
   reg __422988_422988;
   reg _422989_422989 ; 
   reg __422989_422989;
   reg _422990_422990 ; 
   reg __422990_422990;
   reg _422991_422991 ; 
   reg __422991_422991;
   reg _422992_422992 ; 
   reg __422992_422992;
   reg _422993_422993 ; 
   reg __422993_422993;
   reg _422994_422994 ; 
   reg __422994_422994;
   reg _422995_422995 ; 
   reg __422995_422995;
   reg _422996_422996 ; 
   reg __422996_422996;
   reg _422997_422997 ; 
   reg __422997_422997;
   reg _422998_422998 ; 
   reg __422998_422998;
   reg _422999_422999 ; 
   reg __422999_422999;
   reg _423000_423000 ; 
   reg __423000_423000;
   reg _423001_423001 ; 
   reg __423001_423001;
   reg _423002_423002 ; 
   reg __423002_423002;
   reg _423003_423003 ; 
   reg __423003_423003;
   reg _423004_423004 ; 
   reg __423004_423004;
   reg _423005_423005 ; 
   reg __423005_423005;
   reg _423006_423006 ; 
   reg __423006_423006;
   reg _423007_423007 ; 
   reg __423007_423007;
   reg _423008_423008 ; 
   reg __423008_423008;
   reg _423009_423009 ; 
   reg __423009_423009;
   reg _423010_423010 ; 
   reg __423010_423010;
   reg _423011_423011 ; 
   reg __423011_423011;
   reg _423012_423012 ; 
   reg __423012_423012;
   reg _423013_423013 ; 
   reg __423013_423013;
   reg _423014_423014 ; 
   reg __423014_423014;
   reg _423015_423015 ; 
   reg __423015_423015;
   reg _423016_423016 ; 
   reg __423016_423016;
   reg _423017_423017 ; 
   reg __423017_423017;
   reg _423018_423018 ; 
   reg __423018_423018;
   reg _423019_423019 ; 
   reg __423019_423019;
   reg _423020_423020 ; 
   reg __423020_423020;
   reg _423021_423021 ; 
   reg __423021_423021;
   reg _423022_423022 ; 
   reg __423022_423022;
   reg _423023_423023 ; 
   reg __423023_423023;
   reg _423024_423024 ; 
   reg __423024_423024;
   reg _423025_423025 ; 
   reg __423025_423025;
   reg _423026_423026 ; 
   reg __423026_423026;
   reg _423027_423027 ; 
   reg __423027_423027;
   reg _423028_423028 ; 
   reg __423028_423028;
   reg _423029_423029 ; 
   reg __423029_423029;
   reg _423030_423030 ; 
   reg __423030_423030;
   reg _423031_423031 ; 
   reg __423031_423031;
   reg _423032_423032 ; 
   reg __423032_423032;
   reg _423033_423033 ; 
   reg __423033_423033;
   reg _423034_423034 ; 
   reg __423034_423034;
   reg _423035_423035 ; 
   reg __423035_423035;
   reg _423036_423036 ; 
   reg __423036_423036;
   reg _423037_423037 ; 
   reg __423037_423037;
   reg _423038_423038 ; 
   reg __423038_423038;
   reg _423039_423039 ; 
   reg __423039_423039;
   reg _423040_423040 ; 
   reg __423040_423040;
   reg _423041_423041 ; 
   reg __423041_423041;
   reg _423042_423042 ; 
   reg __423042_423042;
   reg _423043_423043 ; 
   reg __423043_423043;
   reg _423044_423044 ; 
   reg __423044_423044;
   reg _423045_423045 ; 
   reg __423045_423045;
   reg _423046_423046 ; 
   reg __423046_423046;
   reg _423047_423047 ; 
   reg __423047_423047;
   reg _423048_423048 ; 
   reg __423048_423048;
   reg _423049_423049 ; 
   reg __423049_423049;
   reg _423050_423050 ; 
   reg __423050_423050;
   reg _423051_423051 ; 
   reg __423051_423051;
   reg _423052_423052 ; 
   reg __423052_423052;
   reg _423053_423053 ; 
   reg __423053_423053;
   reg _423054_423054 ; 
   reg __423054_423054;
   reg _423055_423055 ; 
   reg __423055_423055;
   reg _423056_423056 ; 
   reg __423056_423056;
   reg _423057_423057 ; 
   reg __423057_423057;
   reg _423058_423058 ; 
   reg __423058_423058;
   reg _423059_423059 ; 
   reg __423059_423059;
   reg _423060_423060 ; 
   reg __423060_423060;
   reg _423061_423061 ; 
   reg __423061_423061;
   reg _423062_423062 ; 
   reg __423062_423062;
   reg _423063_423063 ; 
   reg __423063_423063;
   reg _423064_423064 ; 
   reg __423064_423064;
   reg _423065_423065 ; 
   reg __423065_423065;
   reg _423066_423066 ; 
   reg __423066_423066;
   reg _423067_423067 ; 
   reg __423067_423067;
   reg _423068_423068 ; 
   reg __423068_423068;
   reg _423069_423069 ; 
   reg __423069_423069;
   reg _423070_423070 ; 
   reg __423070_423070;
   reg _423071_423071 ; 
   reg __423071_423071;
   reg _423072_423072 ; 
   reg __423072_423072;
   reg _423073_423073 ; 
   reg __423073_423073;
   reg _423074_423074 ; 
   reg __423074_423074;
   reg _423075_423075 ; 
   reg __423075_423075;
   reg _423076_423076 ; 
   reg __423076_423076;
   reg _423077_423077 ; 
   reg __423077_423077;
   reg _423078_423078 ; 
   reg __423078_423078;
   reg _423079_423079 ; 
   reg __423079_423079;
   reg _423080_423080 ; 
   reg __423080_423080;
   reg _423081_423081 ; 
   reg __423081_423081;
   reg _423082_423082 ; 
   reg __423082_423082;
   reg _423083_423083 ; 
   reg __423083_423083;
   reg _423084_423084 ; 
   reg __423084_423084;
   reg _423085_423085 ; 
   reg __423085_423085;
   reg _423086_423086 ; 
   reg __423086_423086;
   reg _423087_423087 ; 
   reg __423087_423087;
   reg _423088_423088 ; 
   reg __423088_423088;
   reg _423089_423089 ; 
   reg __423089_423089;
   reg _423090_423090 ; 
   reg __423090_423090;
   reg _423091_423091 ; 
   reg __423091_423091;
   reg _423092_423092 ; 
   reg __423092_423092;
   reg _423093_423093 ; 
   reg __423093_423093;
   reg _423094_423094 ; 
   reg __423094_423094;
   reg _423095_423095 ; 
   reg __423095_423095;
   reg _423096_423096 ; 
   reg __423096_423096;
   reg _423097_423097 ; 
   reg __423097_423097;
   reg _423098_423098 ; 
   reg __423098_423098;
   reg _423099_423099 ; 
   reg __423099_423099;
   reg _423100_423100 ; 
   reg __423100_423100;
   reg _423101_423101 ; 
   reg __423101_423101;
   reg _423102_423102 ; 
   reg __423102_423102;
   reg _423103_423103 ; 
   reg __423103_423103;
   reg _423104_423104 ; 
   reg __423104_423104;
   reg _423105_423105 ; 
   reg __423105_423105;
   reg _423106_423106 ; 
   reg __423106_423106;
   reg _423107_423107 ; 
   reg __423107_423107;
   reg _423108_423108 ; 
   reg __423108_423108;
   reg _423109_423109 ; 
   reg __423109_423109;
   reg _423110_423110 ; 
   reg __423110_423110;
   reg _423111_423111 ; 
   reg __423111_423111;
   reg _423112_423112 ; 
   reg __423112_423112;
   reg _423113_423113 ; 
   reg __423113_423113;
   reg _423114_423114 ; 
   reg __423114_423114;
   reg _423115_423115 ; 
   reg __423115_423115;
   reg _423116_423116 ; 
   reg __423116_423116;
   reg _423117_423117 ; 
   reg __423117_423117;
   reg _423118_423118 ; 
   reg __423118_423118;
   reg _423119_423119 ; 
   reg __423119_423119;
   reg _423120_423120 ; 
   reg __423120_423120;
   reg _423121_423121 ; 
   reg __423121_423121;
   reg _423122_423122 ; 
   reg __423122_423122;
   reg _423123_423123 ; 
   reg __423123_423123;
   reg _423124_423124 ; 
   reg __423124_423124;
   reg _423125_423125 ; 
   reg __423125_423125;
   reg _423126_423126 ; 
   reg __423126_423126;
   reg _423127_423127 ; 
   reg __423127_423127;
   reg _423128_423128 ; 
   reg __423128_423128;
   reg _423129_423129 ; 
   reg __423129_423129;
   reg _423130_423130 ; 
   reg __423130_423130;
   reg _423131_423131 ; 
   reg __423131_423131;
   reg _423132_423132 ; 
   reg __423132_423132;
   reg _423133_423133 ; 
   reg __423133_423133;
   reg _423134_423134 ; 
   reg __423134_423134;
   reg _423135_423135 ; 
   reg __423135_423135;
   reg _423136_423136 ; 
   reg __423136_423136;
   reg _423137_423137 ; 
   reg __423137_423137;
   reg _423138_423138 ; 
   reg __423138_423138;
   reg _423139_423139 ; 
   reg __423139_423139;
   reg _423140_423140 ; 
   reg __423140_423140;
   reg _423141_423141 ; 
   reg __423141_423141;
   reg _423142_423142 ; 
   reg __423142_423142;
   reg _423143_423143 ; 
   reg __423143_423143;
   reg _423144_423144 ; 
   reg __423144_423144;
   reg _423145_423145 ; 
   reg __423145_423145;
   reg _423146_423146 ; 
   reg __423146_423146;
   reg _423147_423147 ; 
   reg __423147_423147;
   reg _423148_423148 ; 
   reg __423148_423148;
   reg _423149_423149 ; 
   reg __423149_423149;
   reg _423150_423150 ; 
   reg __423150_423150;
   reg _423151_423151 ; 
   reg __423151_423151;
   reg _423152_423152 ; 
   reg __423152_423152;
   reg _423153_423153 ; 
   reg __423153_423153;
   reg _423154_423154 ; 
   reg __423154_423154;
   reg _423155_423155 ; 
   reg __423155_423155;
   reg _423156_423156 ; 
   reg __423156_423156;
   reg _423157_423157 ; 
   reg __423157_423157;
   reg _423158_423158 ; 
   reg __423158_423158;
   reg _423159_423159 ; 
   reg __423159_423159;
   reg _423160_423160 ; 
   reg __423160_423160;
   reg _423161_423161 ; 
   reg __423161_423161;
   reg _423162_423162 ; 
   reg __423162_423162;
   reg _423163_423163 ; 
   reg __423163_423163;
   reg _423164_423164 ; 
   reg __423164_423164;
   reg _423165_423165 ; 
   reg __423165_423165;
   reg _423166_423166 ; 
   reg __423166_423166;
   reg _423167_423167 ; 
   reg __423167_423167;
   reg _423168_423168 ; 
   reg __423168_423168;
   reg _423169_423169 ; 
   reg __423169_423169;
   reg _423170_423170 ; 
   reg __423170_423170;
   reg _423171_423171 ; 
   reg __423171_423171;
   reg _423172_423172 ; 
   reg __423172_423172;
   reg _423173_423173 ; 
   reg __423173_423173;
   reg _423174_423174 ; 
   reg __423174_423174;
   reg _423175_423175 ; 
   reg __423175_423175;
   reg _423176_423176 ; 
   reg __423176_423176;
   reg _423177_423177 ; 
   reg __423177_423177;
   reg _423178_423178 ; 
   reg __423178_423178;
   reg _423179_423179 ; 
   reg __423179_423179;
   reg _423180_423180 ; 
   reg __423180_423180;
   reg _423181_423181 ; 
   reg __423181_423181;
   reg _423182_423182 ; 
   reg __423182_423182;
   reg _423183_423183 ; 
   reg __423183_423183;
   reg _423184_423184 ; 
   reg __423184_423184;
   reg _423185_423185 ; 
   reg __423185_423185;
   reg _423186_423186 ; 
   reg __423186_423186;
   reg _423187_423187 ; 
   reg __423187_423187;
   reg _423188_423188 ; 
   reg __423188_423188;
   reg _423189_423189 ; 
   reg __423189_423189;
   reg _423190_423190 ; 
   reg __423190_423190;
   reg _423191_423191 ; 
   reg __423191_423191;
   reg _423192_423192 ; 
   reg __423192_423192;
   reg _423193_423193 ; 
   reg __423193_423193;
   reg _423194_423194 ; 
   reg __423194_423194;
   reg _423195_423195 ; 
   reg __423195_423195;
   reg _423196_423196 ; 
   reg __423196_423196;
   reg _423197_423197 ; 
   reg __423197_423197;
   reg _423198_423198 ; 
   reg __423198_423198;
   reg _423199_423199 ; 
   reg __423199_423199;
   reg _423200_423200 ; 
   reg __423200_423200;
   reg _423201_423201 ; 
   reg __423201_423201;
   reg _423202_423202 ; 
   reg __423202_423202;
   reg _423203_423203 ; 
   reg __423203_423203;
   reg _423204_423204 ; 
   reg __423204_423204;
   reg _423205_423205 ; 
   reg __423205_423205;
   reg _423206_423206 ; 
   reg __423206_423206;
   reg _423207_423207 ; 
   reg __423207_423207;
   reg _423208_423208 ; 
   reg __423208_423208;
   reg _423209_423209 ; 
   reg __423209_423209;
   reg _423210_423210 ; 
   reg __423210_423210;
   reg _423211_423211 ; 
   reg __423211_423211;
   reg _423212_423212 ; 
   reg __423212_423212;
   reg _423213_423213 ; 
   reg __423213_423213;
   reg _423214_423214 ; 
   reg __423214_423214;
   reg _423215_423215 ; 
   reg __423215_423215;
   reg _423216_423216 ; 
   reg __423216_423216;
   reg _423217_423217 ; 
   reg __423217_423217;
   reg _423218_423218 ; 
   reg __423218_423218;
   reg _423219_423219 ; 
   reg __423219_423219;
   reg _423220_423220 ; 
   reg __423220_423220;
   reg _423221_423221 ; 
   reg __423221_423221;
   reg _423222_423222 ; 
   reg __423222_423222;
   reg _423223_423223 ; 
   reg __423223_423223;
   reg _423224_423224 ; 
   reg __423224_423224;
   reg _423225_423225 ; 
   reg __423225_423225;
   reg _423226_423226 ; 
   reg __423226_423226;
   reg _423227_423227 ; 
   reg __423227_423227;
   reg _423228_423228 ; 
   reg __423228_423228;
   reg _423229_423229 ; 
   reg __423229_423229;
   reg _423230_423230 ; 
   reg __423230_423230;
   reg _423231_423231 ; 
   reg __423231_423231;
   reg _423232_423232 ; 
   reg __423232_423232;
   reg _423233_423233 ; 
   reg __423233_423233;
   reg _423234_423234 ; 
   reg __423234_423234;
   reg _423235_423235 ; 
   reg __423235_423235;
   reg _423236_423236 ; 
   reg __423236_423236;
   reg _423237_423237 ; 
   reg __423237_423237;
   reg _423238_423238 ; 
   reg __423238_423238;
   reg _423239_423239 ; 
   reg __423239_423239;
   reg _423240_423240 ; 
   reg __423240_423240;
   reg _423241_423241 ; 
   reg __423241_423241;
   reg _423242_423242 ; 
   reg __423242_423242;
   reg _423243_423243 ; 
   reg __423243_423243;
   reg _423244_423244 ; 
   reg __423244_423244;
   reg _423245_423245 ; 
   reg __423245_423245;
   reg _423246_423246 ; 
   reg __423246_423246;
   reg _423247_423247 ; 
   reg __423247_423247;
   reg _423248_423248 ; 
   reg __423248_423248;
   reg _423249_423249 ; 
   reg __423249_423249;
   reg _423250_423250 ; 
   reg __423250_423250;
   reg _423251_423251 ; 
   reg __423251_423251;
   reg _423252_423252 ; 
   reg __423252_423252;
   reg _423253_423253 ; 
   reg __423253_423253;
   reg _423254_423254 ; 
   reg __423254_423254;
   reg _423255_423255 ; 
   reg __423255_423255;
   reg _423256_423256 ; 
   reg __423256_423256;
   reg _423257_423257 ; 
   reg __423257_423257;
   reg _423258_423258 ; 
   reg __423258_423258;
   reg _423259_423259 ; 
   reg __423259_423259;
   reg _423260_423260 ; 
   reg __423260_423260;
   reg _423261_423261 ; 
   reg __423261_423261;
   reg _423262_423262 ; 
   reg __423262_423262;
   reg _423263_423263 ; 
   reg __423263_423263;
   reg _423264_423264 ; 
   reg __423264_423264;
   reg _423265_423265 ; 
   reg __423265_423265;
   reg _423266_423266 ; 
   reg __423266_423266;
   reg _423267_423267 ; 
   reg __423267_423267;
   reg _423268_423268 ; 
   reg __423268_423268;
   reg _423269_423269 ; 
   reg __423269_423269;
   reg _423270_423270 ; 
   reg __423270_423270;
   reg _423271_423271 ; 
   reg __423271_423271;
   reg _423272_423272 ; 
   reg __423272_423272;
   reg _423273_423273 ; 
   reg __423273_423273;
   reg _423274_423274 ; 
   reg __423274_423274;
   reg _423275_423275 ; 
   reg __423275_423275;
   reg _423276_423276 ; 
   reg __423276_423276;
   reg _423277_423277 ; 
   reg __423277_423277;
   reg _423278_423278 ; 
   reg __423278_423278;
   reg _423279_423279 ; 
   reg __423279_423279;
   reg _423280_423280 ; 
   reg __423280_423280;
   reg _423281_423281 ; 
   reg __423281_423281;
   reg _423282_423282 ; 
   reg __423282_423282;
   reg _423283_423283 ; 
   reg __423283_423283;
   reg _423284_423284 ; 
   reg __423284_423284;
   reg _423285_423285 ; 
   reg __423285_423285;
   reg _423286_423286 ; 
   reg __423286_423286;
   reg _423287_423287 ; 
   reg __423287_423287;
   reg _423288_423288 ; 
   reg __423288_423288;
   reg _423289_423289 ; 
   reg __423289_423289;
   reg _423290_423290 ; 
   reg __423290_423290;
   reg _423291_423291 ; 
   reg __423291_423291;
   reg _423292_423292 ; 
   reg __423292_423292;
   reg _423293_423293 ; 
   reg __423293_423293;
   reg _423294_423294 ; 
   reg __423294_423294;
   reg _423295_423295 ; 
   reg __423295_423295;
   reg _423296_423296 ; 
   reg __423296_423296;
   reg _423297_423297 ; 
   reg __423297_423297;
   reg _423298_423298 ; 
   reg __423298_423298;
   reg _423299_423299 ; 
   reg __423299_423299;
   reg _423300_423300 ; 
   reg __423300_423300;
   reg _423301_423301 ; 
   reg __423301_423301;
   reg _423302_423302 ; 
   reg __423302_423302;
   reg _423303_423303 ; 
   reg __423303_423303;
   reg _423304_423304 ; 
   reg __423304_423304;
   reg _423305_423305 ; 
   reg __423305_423305;
   reg _423306_423306 ; 
   reg __423306_423306;
   reg _423307_423307 ; 
   reg __423307_423307;
   reg _423308_423308 ; 
   reg __423308_423308;
   reg _423309_423309 ; 
   reg __423309_423309;
   reg _423310_423310 ; 
   reg __423310_423310;
   reg _423311_423311 ; 
   reg __423311_423311;
   reg _423312_423312 ; 
   reg __423312_423312;
   reg _423313_423313 ; 
   reg __423313_423313;
   reg _423314_423314 ; 
   reg __423314_423314;
   reg _423315_423315 ; 
   reg __423315_423315;
   reg _423316_423316 ; 
   reg __423316_423316;
   reg _423317_423317 ; 
   reg __423317_423317;
   reg _423318_423318 ; 
   reg __423318_423318;
   reg _423319_423319 ; 
   reg __423319_423319;
   reg _423320_423320 ; 
   reg __423320_423320;
   reg _423321_423321 ; 
   reg __423321_423321;
   reg _423322_423322 ; 
   reg __423322_423322;
   reg _423323_423323 ; 
   reg __423323_423323;
   reg _423324_423324 ; 
   reg __423324_423324;
   reg _423325_423325 ; 
   reg __423325_423325;
   reg _423326_423326 ; 
   reg __423326_423326;
   reg _423327_423327 ; 
   reg __423327_423327;
   reg _423328_423328 ; 
   reg __423328_423328;
   reg _423329_423329 ; 
   reg __423329_423329;
   reg _423330_423330 ; 
   reg __423330_423330;
   reg _423331_423331 ; 
   reg __423331_423331;
   reg _423332_423332 ; 
   reg __423332_423332;
   reg _423333_423333 ; 
   reg __423333_423333;
   reg _423334_423334 ; 
   reg __423334_423334;
   reg _423335_423335 ; 
   reg __423335_423335;
   reg _423336_423336 ; 
   reg __423336_423336;
   reg _423337_423337 ; 
   reg __423337_423337;
   reg _423338_423338 ; 
   reg __423338_423338;
   reg _423339_423339 ; 
   reg __423339_423339;
   reg _423340_423340 ; 
   reg __423340_423340;
   reg _423341_423341 ; 
   reg __423341_423341;
   reg _423342_423342 ; 
   reg __423342_423342;
   reg _423343_423343 ; 
   reg __423343_423343;
   reg _423344_423344 ; 
   reg __423344_423344;
   reg _423345_423345 ; 
   reg __423345_423345;
   reg _423346_423346 ; 
   reg __423346_423346;
   reg _423347_423347 ; 
   reg __423347_423347;
   reg _423348_423348 ; 
   reg __423348_423348;
   reg _423349_423349 ; 
   reg __423349_423349;
   reg _423350_423350 ; 
   reg __423350_423350;
   reg _423351_423351 ; 
   reg __423351_423351;
   reg _423352_423352 ; 
   reg __423352_423352;
   reg _423353_423353 ; 
   reg __423353_423353;
   reg _423354_423354 ; 
   reg __423354_423354;
   reg _423355_423355 ; 
   reg __423355_423355;
   reg _423356_423356 ; 
   reg __423356_423356;
   reg _423357_423357 ; 
   reg __423357_423357;
   reg _423358_423358 ; 
   reg __423358_423358;
   reg _423359_423359 ; 
   reg __423359_423359;
   reg _423360_423360 ; 
   reg __423360_423360;
   reg _423361_423361 ; 
   reg __423361_423361;
   reg _423362_423362 ; 
   reg __423362_423362;
   reg _423363_423363 ; 
   reg __423363_423363;
   reg _423364_423364 ; 
   reg __423364_423364;
   reg _423365_423365 ; 
   reg __423365_423365;
   reg _423366_423366 ; 
   reg __423366_423366;
   reg _423367_423367 ; 
   reg __423367_423367;
   reg _423368_423368 ; 
   reg __423368_423368;
   reg _423369_423369 ; 
   reg __423369_423369;
   reg _423370_423370 ; 
   reg __423370_423370;
   reg _423371_423371 ; 
   reg __423371_423371;
   reg _423372_423372 ; 
   reg __423372_423372;
   reg _423373_423373 ; 
   reg __423373_423373;
   reg _423374_423374 ; 
   reg __423374_423374;
   reg _423375_423375 ; 
   reg __423375_423375;
   reg _423376_423376 ; 
   reg __423376_423376;
   reg _423377_423377 ; 
   reg __423377_423377;
   reg _423378_423378 ; 
   reg __423378_423378;
   reg _423379_423379 ; 
   reg __423379_423379;
   reg _423380_423380 ; 
   reg __423380_423380;
   reg _423381_423381 ; 
   reg __423381_423381;
   reg _423382_423382 ; 
   reg __423382_423382;
   reg _423383_423383 ; 
   reg __423383_423383;
   reg _423384_423384 ; 
   reg __423384_423384;
   reg _423385_423385 ; 
   reg __423385_423385;
   reg _423386_423386 ; 
   reg __423386_423386;
   reg _423387_423387 ; 
   reg __423387_423387;
   reg _423388_423388 ; 
   reg __423388_423388;
   reg _423389_423389 ; 
   reg __423389_423389;
   reg _423390_423390 ; 
   reg __423390_423390;
   reg _423391_423391 ; 
   reg __423391_423391;
   reg _423392_423392 ; 
   reg __423392_423392;
   reg _423393_423393 ; 
   reg __423393_423393;
   reg _423394_423394 ; 
   reg __423394_423394;
   reg _423395_423395 ; 
   reg __423395_423395;
   reg _423396_423396 ; 
   reg __423396_423396;
   reg _423397_423397 ; 
   reg __423397_423397;
   reg _423398_423398 ; 
   reg __423398_423398;
   reg _423399_423399 ; 
   reg __423399_423399;
   reg _423400_423400 ; 
   reg __423400_423400;
   reg _423401_423401 ; 
   reg __423401_423401;
   reg _423402_423402 ; 
   reg __423402_423402;
   reg _423403_423403 ; 
   reg __423403_423403;
   reg _423404_423404 ; 
   reg __423404_423404;
   reg _423405_423405 ; 
   reg __423405_423405;
   reg _423406_423406 ; 
   reg __423406_423406;
   reg _423407_423407 ; 
   reg __423407_423407;
   reg _423408_423408 ; 
   reg __423408_423408;
   reg _423409_423409 ; 
   reg __423409_423409;
   reg _423410_423410 ; 
   reg __423410_423410;
   reg _423411_423411 ; 
   reg __423411_423411;
   reg _423412_423412 ; 
   reg __423412_423412;
   reg _423413_423413 ; 
   reg __423413_423413;
   reg _423414_423414 ; 
   reg __423414_423414;
   reg _423415_423415 ; 
   reg __423415_423415;
   reg _423416_423416 ; 
   reg __423416_423416;
   reg _423417_423417 ; 
   reg __423417_423417;
   reg _423418_423418 ; 
   reg __423418_423418;
   reg _423419_423419 ; 
   reg __423419_423419;
   reg _423420_423420 ; 
   reg __423420_423420;
   reg _423421_423421 ; 
   reg __423421_423421;
   reg _423422_423422 ; 
   reg __423422_423422;
   reg _423423_423423 ; 
   reg __423423_423423;
   reg _423424_423424 ; 
   reg __423424_423424;
   reg _423425_423425 ; 
   reg __423425_423425;
   reg _423426_423426 ; 
   reg __423426_423426;
   reg _423427_423427 ; 
   reg __423427_423427;
   reg _423428_423428 ; 
   reg __423428_423428;
   reg _423429_423429 ; 
   reg __423429_423429;
   reg _423430_423430 ; 
   reg __423430_423430;
   reg _423431_423431 ; 
   reg __423431_423431;
   reg _423432_423432 ; 
   reg __423432_423432;
   reg _423433_423433 ; 
   reg __423433_423433;
   reg _423434_423434 ; 
   reg __423434_423434;
   reg _423435_423435 ; 
   reg __423435_423435;
   reg _423436_423436 ; 
   reg __423436_423436;
   reg _423437_423437 ; 
   reg __423437_423437;
   reg _423438_423438 ; 
   reg __423438_423438;
   reg _423439_423439 ; 
   reg __423439_423439;
   reg _423440_423440 ; 
   reg __423440_423440;
   reg _423441_423441 ; 
   reg __423441_423441;
   reg _423442_423442 ; 
   reg __423442_423442;
   reg _423443_423443 ; 
   reg __423443_423443;
   reg _423444_423444 ; 
   reg __423444_423444;
   reg _423445_423445 ; 
   reg __423445_423445;
   reg _423446_423446 ; 
   reg __423446_423446;
   reg _423447_423447 ; 
   reg __423447_423447;
   reg _423448_423448 ; 
   reg __423448_423448;
   reg _423449_423449 ; 
   reg __423449_423449;
   reg _423450_423450 ; 
   reg __423450_423450;
   reg _423451_423451 ; 
   reg __423451_423451;
   reg _423452_423452 ; 
   reg __423452_423452;
   reg _423453_423453 ; 
   reg __423453_423453;
   reg _423454_423454 ; 
   reg __423454_423454;
   reg _423455_423455 ; 
   reg __423455_423455;
   reg _423456_423456 ; 
   reg __423456_423456;
   reg _423457_423457 ; 
   reg __423457_423457;
   reg _423458_423458 ; 
   reg __423458_423458;
   reg _423459_423459 ; 
   reg __423459_423459;
   reg _423460_423460 ; 
   reg __423460_423460;
   reg _423461_423461 ; 
   reg __423461_423461;
   reg _423462_423462 ; 
   reg __423462_423462;
   reg _423463_423463 ; 
   reg __423463_423463;
   reg _423464_423464 ; 
   reg __423464_423464;
   reg _423465_423465 ; 
   reg __423465_423465;
   reg _423466_423466 ; 
   reg __423466_423466;
   reg _423467_423467 ; 
   reg __423467_423467;
   reg _423468_423468 ; 
   reg __423468_423468;
   reg _423469_423469 ; 
   reg __423469_423469;
   reg _423470_423470 ; 
   reg __423470_423470;
   reg _423471_423471 ; 
   reg __423471_423471;
   reg _423472_423472 ; 
   reg __423472_423472;
   reg _423473_423473 ; 
   reg __423473_423473;
   reg _423474_423474 ; 
   reg __423474_423474;
   reg _423475_423475 ; 
   reg __423475_423475;
   reg _423476_423476 ; 
   reg __423476_423476;
   reg _423477_423477 ; 
   reg __423477_423477;
   reg _423478_423478 ; 
   reg __423478_423478;
   reg _423479_423479 ; 
   reg __423479_423479;
   reg _423480_423480 ; 
   reg __423480_423480;
   reg _423481_423481 ; 
   reg __423481_423481;
   reg _423482_423482 ; 
   reg __423482_423482;
   reg _423483_423483 ; 
   reg __423483_423483;
   reg _423484_423484 ; 
   reg __423484_423484;
   reg _423485_423485 ; 
   reg __423485_423485;
   reg _423486_423486 ; 
   reg __423486_423486;
   reg _423487_423487 ; 
   reg __423487_423487;
   reg _423488_423488 ; 
   reg __423488_423488;
   reg _423489_423489 ; 
   reg __423489_423489;
   reg _423490_423490 ; 
   reg __423490_423490;
   reg _423491_423491 ; 
   reg __423491_423491;
   reg _423492_423492 ; 
   reg __423492_423492;
   reg _423493_423493 ; 
   reg __423493_423493;
   reg _423494_423494 ; 
   reg __423494_423494;
   reg _423495_423495 ; 
   reg __423495_423495;
   reg _423496_423496 ; 
   reg __423496_423496;
   reg _423497_423497 ; 
   reg __423497_423497;
   reg _423498_423498 ; 
   reg __423498_423498;
   reg _423499_423499 ; 
   reg __423499_423499;
   reg _423500_423500 ; 
   reg __423500_423500;
   reg _423501_423501 ; 
   reg __423501_423501;
   reg _423502_423502 ; 
   reg __423502_423502;
   reg _423503_423503 ; 
   reg __423503_423503;
   reg _423504_423504 ; 
   reg __423504_423504;
   reg _423505_423505 ; 
   reg __423505_423505;
   reg _423506_423506 ; 
   reg __423506_423506;
   reg _423507_423507 ; 
   reg __423507_423507;
   reg _423508_423508 ; 
   reg __423508_423508;
   reg _423509_423509 ; 
   reg __423509_423509;
   reg _423510_423510 ; 
   reg __423510_423510;
   reg _423511_423511 ; 
   reg __423511_423511;
   reg _423512_423512 ; 
   reg __423512_423512;
   reg _423513_423513 ; 
   reg __423513_423513;
   reg _423514_423514 ; 
   reg __423514_423514;
   reg _423515_423515 ; 
   reg __423515_423515;
   reg _423516_423516 ; 
   reg __423516_423516;
   reg _423517_423517 ; 
   reg __423517_423517;
   reg _423518_423518 ; 
   reg __423518_423518;
   reg _423519_423519 ; 
   reg __423519_423519;
   reg _423520_423520 ; 
   reg __423520_423520;
   reg _423521_423521 ; 
   reg __423521_423521;
   reg _423522_423522 ; 
   reg __423522_423522;
   reg _423523_423523 ; 
   reg __423523_423523;
   reg _423524_423524 ; 
   reg __423524_423524;
   reg _423525_423525 ; 
   reg __423525_423525;
   reg _423526_423526 ; 
   reg __423526_423526;
   reg _423527_423527 ; 
   reg __423527_423527;
   reg _423528_423528 ; 
   reg __423528_423528;
   reg _423529_423529 ; 
   reg __423529_423529;
   reg _423530_423530 ; 
   reg __423530_423530;
   reg _423531_423531 ; 
   reg __423531_423531;
   reg _423532_423532 ; 
   reg __423532_423532;
   reg _423533_423533 ; 
   reg __423533_423533;
   reg _423534_423534 ; 
   reg __423534_423534;
   reg _423535_423535 ; 
   reg __423535_423535;
   reg _423536_423536 ; 
   reg __423536_423536;
   reg _423537_423537 ; 
   reg __423537_423537;
   reg _423538_423538 ; 
   reg __423538_423538;
   reg _423539_423539 ; 
   reg __423539_423539;
   reg _423540_423540 ; 
   reg __423540_423540;
   reg _423541_423541 ; 
   reg __423541_423541;
   reg _423542_423542 ; 
   reg __423542_423542;
   reg _423543_423543 ; 
   reg __423543_423543;
   reg _423544_423544 ; 
   reg __423544_423544;
   reg _423545_423545 ; 
   reg __423545_423545;
   reg _423546_423546 ; 
   reg __423546_423546;
   reg _423547_423547 ; 
   reg __423547_423547;
   reg _423548_423548 ; 
   reg __423548_423548;
   reg _423549_423549 ; 
   reg __423549_423549;
   reg _423550_423550 ; 
   reg __423550_423550;
   reg _423551_423551 ; 
   reg __423551_423551;
   reg _423552_423552 ; 
   reg __423552_423552;
   reg _423553_423553 ; 
   reg __423553_423553;
   reg _423554_423554 ; 
   reg __423554_423554;
   reg _423555_423555 ; 
   reg __423555_423555;
   reg _423556_423556 ; 
   reg __423556_423556;
   reg _423557_423557 ; 
   reg __423557_423557;
   reg _423558_423558 ; 
   reg __423558_423558;
   reg _423559_423559 ; 
   reg __423559_423559;
   reg _423560_423560 ; 
   reg __423560_423560;
   reg _423561_423561 ; 
   reg __423561_423561;
   reg _423562_423562 ; 
   reg __423562_423562;
   reg _423563_423563 ; 
   reg __423563_423563;
   reg _423564_423564 ; 
   reg __423564_423564;
   reg _423565_423565 ; 
   reg __423565_423565;
   reg _423566_423566 ; 
   reg __423566_423566;
   reg _423567_423567 ; 
   reg __423567_423567;
   reg _423568_423568 ; 
   reg __423568_423568;
   reg _423569_423569 ; 
   reg __423569_423569;
   reg _423570_423570 ; 
   reg __423570_423570;
   reg _423571_423571 ; 
   reg __423571_423571;
   reg _423572_423572 ; 
   reg __423572_423572;
   reg _423573_423573 ; 
   reg __423573_423573;
   reg _423574_423574 ; 
   reg __423574_423574;
   reg _423575_423575 ; 
   reg __423575_423575;
   reg _423576_423576 ; 
   reg __423576_423576;
   reg _423577_423577 ; 
   reg __423577_423577;
   reg _423578_423578 ; 
   reg __423578_423578;
   reg _423579_423579 ; 
   reg __423579_423579;
   reg _423580_423580 ; 
   reg __423580_423580;
   reg _423581_423581 ; 
   reg __423581_423581;
   reg _423582_423582 ; 
   reg __423582_423582;
   reg _423583_423583 ; 
   reg __423583_423583;
   reg _423584_423584 ; 
   reg __423584_423584;
   reg _423585_423585 ; 
   reg __423585_423585;
   reg _423586_423586 ; 
   reg __423586_423586;
   reg _423587_423587 ; 
   reg __423587_423587;
   reg _423588_423588 ; 
   reg __423588_423588;
   reg _423589_423589 ; 
   reg __423589_423589;
   reg _423590_423590 ; 
   reg __423590_423590;
   reg _423591_423591 ; 
   reg __423591_423591;
   reg _423592_423592 ; 
   reg __423592_423592;
   reg _423593_423593 ; 
   reg __423593_423593;
   reg _423594_423594 ; 
   reg __423594_423594;
   reg _423595_423595 ; 
   reg __423595_423595;
   reg _423596_423596 ; 
   reg __423596_423596;
   reg _423597_423597 ; 
   reg __423597_423597;
   reg _423598_423598 ; 
   reg __423598_423598;
   reg _423599_423599 ; 
   reg __423599_423599;
   reg _423600_423600 ; 
   reg __423600_423600;
   reg _423601_423601 ; 
   reg __423601_423601;
   reg _423602_423602 ; 
   reg __423602_423602;
   reg _423603_423603 ; 
   reg __423603_423603;
   reg _423604_423604 ; 
   reg __423604_423604;
   reg _423605_423605 ; 
   reg __423605_423605;
   reg _423606_423606 ; 
   reg __423606_423606;
   reg _423607_423607 ; 
   reg __423607_423607;
   reg _423608_423608 ; 
   reg __423608_423608;
   reg _423609_423609 ; 
   reg __423609_423609;
   reg _423610_423610 ; 
   reg __423610_423610;
   reg _423611_423611 ; 
   reg __423611_423611;
   reg _423612_423612 ; 
   reg __423612_423612;
   reg _423613_423613 ; 
   reg __423613_423613;
   reg _423614_423614 ; 
   reg __423614_423614;
   reg _423615_423615 ; 
   reg __423615_423615;
   reg _423616_423616 ; 
   reg __423616_423616;
   reg _423617_423617 ; 
   reg __423617_423617;
   reg _423618_423618 ; 
   reg __423618_423618;
   reg _423619_423619 ; 
   reg __423619_423619;
   reg _423620_423620 ; 
   reg __423620_423620;
   reg _423621_423621 ; 
   reg __423621_423621;
   reg _423622_423622 ; 
   reg __423622_423622;
   reg _423623_423623 ; 
   reg __423623_423623;
   reg _423624_423624 ; 
   reg __423624_423624;
   reg _423625_423625 ; 
   reg __423625_423625;
   reg _423626_423626 ; 
   reg __423626_423626;
   reg _423627_423627 ; 
   reg __423627_423627;
   reg _423628_423628 ; 
   reg __423628_423628;
   reg _423629_423629 ; 
   reg __423629_423629;
   reg _423630_423630 ; 
   reg __423630_423630;
   reg _423631_423631 ; 
   reg __423631_423631;
   reg _423632_423632 ; 
   reg __423632_423632;
   reg _423633_423633 ; 
   reg __423633_423633;
   reg _423634_423634 ; 
   reg __423634_423634;
   reg _423635_423635 ; 
   reg __423635_423635;
   reg _423636_423636 ; 
   reg __423636_423636;
   reg _423637_423637 ; 
   reg __423637_423637;
   reg _423638_423638 ; 
   reg __423638_423638;
   reg _423639_423639 ; 
   reg __423639_423639;
   reg _423640_423640 ; 
   reg __423640_423640;
   reg _423641_423641 ; 
   reg __423641_423641;
   reg _423642_423642 ; 
   reg __423642_423642;
   reg _423643_423643 ; 
   reg __423643_423643;
   reg _423644_423644 ; 
   reg __423644_423644;
   reg _423645_423645 ; 
   reg __423645_423645;
   reg _423646_423646 ; 
   reg __423646_423646;
   reg _423647_423647 ; 
   reg __423647_423647;
   reg _423648_423648 ; 
   reg __423648_423648;
   reg _423649_423649 ; 
   reg __423649_423649;
   reg _423650_423650 ; 
   reg __423650_423650;
   reg _423651_423651 ; 
   reg __423651_423651;
   reg _423652_423652 ; 
   reg __423652_423652;
   reg _423653_423653 ; 
   reg __423653_423653;
   reg _423654_423654 ; 
   reg __423654_423654;
   reg _423655_423655 ; 
   reg __423655_423655;
   reg _423656_423656 ; 
   reg __423656_423656;
   reg _423657_423657 ; 
   reg __423657_423657;
   reg _423658_423658 ; 
   reg __423658_423658;
   reg _423659_423659 ; 
   reg __423659_423659;
   reg _423660_423660 ; 
   reg __423660_423660;
   reg _423661_423661 ; 
   reg __423661_423661;
   reg _423662_423662 ; 
   reg __423662_423662;
   reg _423663_423663 ; 
   reg __423663_423663;
   reg _423664_423664 ; 
   reg __423664_423664;
   reg _423665_423665 ; 
   reg __423665_423665;
   reg _423666_423666 ; 
   reg __423666_423666;
   reg _423667_423667 ; 
   reg __423667_423667;
   reg _423668_423668 ; 
   reg __423668_423668;
   reg _423669_423669 ; 
   reg __423669_423669;
   reg _423670_423670 ; 
   reg __423670_423670;
   reg _423671_423671 ; 
   reg __423671_423671;
   reg _423672_423672 ; 
   reg __423672_423672;
   reg _423673_423673 ; 
   reg __423673_423673;
   reg _423674_423674 ; 
   reg __423674_423674;
   reg _423675_423675 ; 
   reg __423675_423675;
   reg _423676_423676 ; 
   reg __423676_423676;
   reg _423677_423677 ; 
   reg __423677_423677;
   reg _423678_423678 ; 
   reg __423678_423678;
   reg _423679_423679 ; 
   reg __423679_423679;
   reg _423680_423680 ; 
   reg __423680_423680;
   reg _423681_423681 ; 
   reg __423681_423681;
   reg _423682_423682 ; 
   reg __423682_423682;
   reg _423683_423683 ; 
   reg __423683_423683;
   reg _423684_423684 ; 
   reg __423684_423684;
   reg _423685_423685 ; 
   reg __423685_423685;
   reg _423686_423686 ; 
   reg __423686_423686;
   reg _423687_423687 ; 
   reg __423687_423687;
   reg _423688_423688 ; 
   reg __423688_423688;
   reg _423689_423689 ; 
   reg __423689_423689;
   reg _423690_423690 ; 
   reg __423690_423690;
   reg _423691_423691 ; 
   reg __423691_423691;
   reg _423692_423692 ; 
   reg __423692_423692;
   reg _423693_423693 ; 
   reg __423693_423693;
   reg _423694_423694 ; 
   reg __423694_423694;
   reg _423695_423695 ; 
   reg __423695_423695;
   reg _423696_423696 ; 
   reg __423696_423696;
   reg _423697_423697 ; 
   reg __423697_423697;
   reg _423698_423698 ; 
   reg __423698_423698;
   reg _423699_423699 ; 
   reg __423699_423699;
   reg _423700_423700 ; 
   reg __423700_423700;
   reg _423701_423701 ; 
   reg __423701_423701;
   reg _423702_423702 ; 
   reg __423702_423702;
   reg _423703_423703 ; 
   reg __423703_423703;
   reg _423704_423704 ; 
   reg __423704_423704;
   reg _423705_423705 ; 
   reg __423705_423705;
   reg _423706_423706 ; 
   reg __423706_423706;
   reg _423707_423707 ; 
   reg __423707_423707;
   reg _423708_423708 ; 
   reg __423708_423708;
   reg _423709_423709 ; 
   reg __423709_423709;
   reg _423710_423710 ; 
   reg __423710_423710;
   reg _423711_423711 ; 
   reg __423711_423711;
   reg _423712_423712 ; 
   reg __423712_423712;
   reg _423713_423713 ; 
   reg __423713_423713;
   reg _423714_423714 ; 
   reg __423714_423714;
   reg _423715_423715 ; 
   reg __423715_423715;
   reg _423716_423716 ; 
   reg __423716_423716;
   reg _423717_423717 ; 
   reg __423717_423717;
   reg _423718_423718 ; 
   reg __423718_423718;
   reg _423719_423719 ; 
   reg __423719_423719;
   reg _423720_423720 ; 
   reg __423720_423720;
   reg _423721_423721 ; 
   reg __423721_423721;
   reg _423722_423722 ; 
   reg __423722_423722;
   reg _423723_423723 ; 
   reg __423723_423723;
   reg _423724_423724 ; 
   reg __423724_423724;
   reg _423725_423725 ; 
   reg __423725_423725;
   reg _423726_423726 ; 
   reg __423726_423726;
   reg _423727_423727 ; 
   reg __423727_423727;
   reg _423728_423728 ; 
   reg __423728_423728;
   reg _423729_423729 ; 
   reg __423729_423729;
   reg _423730_423730 ; 
   reg __423730_423730;
   reg _423731_423731 ; 
   reg __423731_423731;
   reg _423732_423732 ; 
   reg __423732_423732;
   reg _423733_423733 ; 
   reg __423733_423733;
   reg _423734_423734 ; 
   reg __423734_423734;
   reg _423735_423735 ; 
   reg __423735_423735;
   reg _423736_423736 ; 
   reg __423736_423736;
   reg _423737_423737 ; 
   reg __423737_423737;
   reg _423738_423738 ; 
   reg __423738_423738;
   reg _423739_423739 ; 
   reg __423739_423739;
   reg _423740_423740 ; 
   reg __423740_423740;
   reg _423741_423741 ; 
   reg __423741_423741;
   reg _423742_423742 ; 
   reg __423742_423742;
   reg _423743_423743 ; 
   reg __423743_423743;
   reg _423744_423744 ; 
   reg __423744_423744;
   reg _423745_423745 ; 
   reg __423745_423745;
   reg _423746_423746 ; 
   reg __423746_423746;
   reg _423747_423747 ; 
   reg __423747_423747;
   reg _423748_423748 ; 
   reg __423748_423748;
   reg _423749_423749 ; 
   reg __423749_423749;
   reg _423750_423750 ; 
   reg __423750_423750;
   reg _423751_423751 ; 
   reg __423751_423751;
   reg _423752_423752 ; 
   reg __423752_423752;
   reg _423753_423753 ; 
   reg __423753_423753;
   reg _423754_423754 ; 
   reg __423754_423754;
   reg _423755_423755 ; 
   reg __423755_423755;
   reg _423756_423756 ; 
   reg __423756_423756;
   reg _423757_423757 ; 
   reg __423757_423757;
   reg _423758_423758 ; 
   reg __423758_423758;
   reg _423759_423759 ; 
   reg __423759_423759;
   reg _423760_423760 ; 
   reg __423760_423760;
   reg _423761_423761 ; 
   reg __423761_423761;
   reg _423762_423762 ; 
   reg __423762_423762;
   reg _423763_423763 ; 
   reg __423763_423763;
   reg _423764_423764 ; 
   reg __423764_423764;
   reg _423765_423765 ; 
   reg __423765_423765;
   reg _423766_423766 ; 
   reg __423766_423766;
   reg _423767_423767 ; 
   reg __423767_423767;
   reg _423768_423768 ; 
   reg __423768_423768;
   reg _423769_423769 ; 
   reg __423769_423769;
   reg _423770_423770 ; 
   reg __423770_423770;
   reg _423771_423771 ; 
   reg __423771_423771;
   reg _423772_423772 ; 
   reg __423772_423772;
   reg _423773_423773 ; 
   reg __423773_423773;
   reg _423774_423774 ; 
   reg __423774_423774;
   reg _423775_423775 ; 
   reg __423775_423775;
   reg _423776_423776 ; 
   reg __423776_423776;
   reg _423777_423777 ; 
   reg __423777_423777;
   reg _423778_423778 ; 
   reg __423778_423778;
   reg _423779_423779 ; 
   reg __423779_423779;
   reg _423780_423780 ; 
   reg __423780_423780;
   reg _423781_423781 ; 
   reg __423781_423781;
   reg _423782_423782 ; 
   reg __423782_423782;
   reg _423783_423783 ; 
   reg __423783_423783;
   reg _423784_423784 ; 
   reg __423784_423784;
   reg _423785_423785 ; 
   reg __423785_423785;
   reg _423786_423786 ; 
   reg __423786_423786;
   reg _423787_423787 ; 
   reg __423787_423787;
   reg _423788_423788 ; 
   reg __423788_423788;
   reg _423789_423789 ; 
   reg __423789_423789;
   reg _423790_423790 ; 
   reg __423790_423790;
   reg _423791_423791 ; 
   reg __423791_423791;
   reg _423792_423792 ; 
   reg __423792_423792;
   reg _423793_423793 ; 
   reg __423793_423793;
   reg _423794_423794 ; 
   reg __423794_423794;
   reg _423795_423795 ; 
   reg __423795_423795;
   reg _423796_423796 ; 
   reg __423796_423796;
   reg _423797_423797 ; 
   reg __423797_423797;
   reg _423798_423798 ; 
   reg __423798_423798;
   reg _423799_423799 ; 
   reg __423799_423799;
   reg _423800_423800 ; 
   reg __423800_423800;
   reg _423801_423801 ; 
   reg __423801_423801;
   reg _423802_423802 ; 
   reg __423802_423802;
   reg _423803_423803 ; 
   reg __423803_423803;
   reg _423804_423804 ; 
   reg __423804_423804;
   reg _423805_423805 ; 
   reg __423805_423805;
   reg _423806_423806 ; 
   reg __423806_423806;
   reg _423807_423807 ; 
   reg __423807_423807;
   reg _423808_423808 ; 
   reg __423808_423808;
   reg _423809_423809 ; 
   reg __423809_423809;
   reg _423810_423810 ; 
   reg __423810_423810;
   reg _423811_423811 ; 
   reg __423811_423811;
   reg _423812_423812 ; 
   reg __423812_423812;
   reg _423813_423813 ; 
   reg __423813_423813;
   reg _423814_423814 ; 
   reg __423814_423814;
   reg _423815_423815 ; 
   reg __423815_423815;
   reg _423816_423816 ; 
   reg __423816_423816;
   reg _423817_423817 ; 
   reg __423817_423817;
   reg _423818_423818 ; 
   reg __423818_423818;
   reg _423819_423819 ; 
   reg __423819_423819;
   reg _423820_423820 ; 
   reg __423820_423820;
   reg _423821_423821 ; 
   reg __423821_423821;
   reg _423822_423822 ; 
   reg __423822_423822;
   reg _423823_423823 ; 
   reg __423823_423823;
   reg _423824_423824 ; 
   reg __423824_423824;
   reg _423825_423825 ; 
   reg __423825_423825;
   reg _423826_423826 ; 
   reg __423826_423826;
   reg _423827_423827 ; 
   reg __423827_423827;
   reg _423828_423828 ; 
   reg __423828_423828;
   reg _423829_423829 ; 
   reg __423829_423829;
   reg _423830_423830 ; 
   reg __423830_423830;
   reg _423831_423831 ; 
   reg __423831_423831;
   reg _423832_423832 ; 
   reg __423832_423832;
   reg _423833_423833 ; 
   reg __423833_423833;
   reg _423834_423834 ; 
   reg __423834_423834;
   reg _423835_423835 ; 
   reg __423835_423835;
   reg _423836_423836 ; 
   reg __423836_423836;
   reg _423837_423837 ; 
   reg __423837_423837;
   reg _423838_423838 ; 
   reg __423838_423838;
   reg _423839_423839 ; 
   reg __423839_423839;
   reg _423840_423840 ; 
   reg __423840_423840;
   reg _423841_423841 ; 
   reg __423841_423841;
   reg _423842_423842 ; 
   reg __423842_423842;
   reg _423843_423843 ; 
   reg __423843_423843;
   reg _423844_423844 ; 
   reg __423844_423844;
   reg _423845_423845 ; 
   reg __423845_423845;
   reg _423846_423846 ; 
   reg __423846_423846;
   reg _423847_423847 ; 
   reg __423847_423847;
   reg _423848_423848 ; 
   reg __423848_423848;
   reg _423849_423849 ; 
   reg __423849_423849;
   reg _423850_423850 ; 
   reg __423850_423850;
   reg _423851_423851 ; 
   reg __423851_423851;
   reg _423852_423852 ; 
   reg __423852_423852;
   reg _423853_423853 ; 
   reg __423853_423853;
   reg _423854_423854 ; 
   reg __423854_423854;
   reg _423855_423855 ; 
   reg __423855_423855;
   reg _423856_423856 ; 
   reg __423856_423856;
   reg _423857_423857 ; 
   reg __423857_423857;
   reg _423858_423858 ; 
   reg __423858_423858;
   reg _423859_423859 ; 
   reg __423859_423859;
   reg _423860_423860 ; 
   reg __423860_423860;
   reg _423861_423861 ; 
   reg __423861_423861;
   reg _423862_423862 ; 
   reg __423862_423862;
   reg _423863_423863 ; 
   reg __423863_423863;
   reg _423864_423864 ; 
   reg __423864_423864;
   reg _423865_423865 ; 
   reg __423865_423865;
   reg _423866_423866 ; 
   reg __423866_423866;
   reg _423867_423867 ; 
   reg __423867_423867;
   reg _423868_423868 ; 
   reg __423868_423868;
   reg _423869_423869 ; 
   reg __423869_423869;
   reg _423870_423870 ; 
   reg __423870_423870;
   reg _423871_423871 ; 
   reg __423871_423871;
   reg _423872_423872 ; 
   reg __423872_423872;
   reg _423873_423873 ; 
   reg __423873_423873;
   reg _423874_423874 ; 
   reg __423874_423874;
   reg _423875_423875 ; 
   reg __423875_423875;
   reg _423876_423876 ; 
   reg __423876_423876;
   reg _423877_423877 ; 
   reg __423877_423877;
   reg _423878_423878 ; 
   reg __423878_423878;
   reg _423879_423879 ; 
   reg __423879_423879;
   reg _423880_423880 ; 
   reg __423880_423880;
   reg _423881_423881 ; 
   reg __423881_423881;
   reg _423882_423882 ; 
   reg __423882_423882;
   reg _423883_423883 ; 
   reg __423883_423883;
   reg _423884_423884 ; 
   reg __423884_423884;
   reg _423885_423885 ; 
   reg __423885_423885;
   reg _423886_423886 ; 
   reg __423886_423886;
   reg _423887_423887 ; 
   reg __423887_423887;
   reg _423888_423888 ; 
   reg __423888_423888;
   reg _423889_423889 ; 
   reg __423889_423889;
   reg _423890_423890 ; 
   reg __423890_423890;
   reg _423891_423891 ; 
   reg __423891_423891;
   reg _423892_423892 ; 
   reg __423892_423892;
   reg _423893_423893 ; 
   reg __423893_423893;
   reg _423894_423894 ; 
   reg __423894_423894;
   reg _423895_423895 ; 
   reg __423895_423895;
   reg _423896_423896 ; 
   reg __423896_423896;
   reg _423897_423897 ; 
   reg __423897_423897;
   reg _423898_423898 ; 
   reg __423898_423898;
   reg _423899_423899 ; 
   reg __423899_423899;
   reg _423900_423900 ; 
   reg __423900_423900;
   reg _423901_423901 ; 
   reg __423901_423901;
   reg _423902_423902 ; 
   reg __423902_423902;
   reg _423903_423903 ; 
   reg __423903_423903;
   reg _423904_423904 ; 
   reg __423904_423904;
   reg _423905_423905 ; 
   reg __423905_423905;
   reg _423906_423906 ; 
   reg __423906_423906;
   reg _423907_423907 ; 
   reg __423907_423907;
   reg _423908_423908 ; 
   reg __423908_423908;
   reg _423909_423909 ; 
   reg __423909_423909;
   reg _423910_423910 ; 
   reg __423910_423910;
   reg _423911_423911 ; 
   reg __423911_423911;
   reg _423912_423912 ; 
   reg __423912_423912;
   reg _423913_423913 ; 
   reg __423913_423913;
   reg _423914_423914 ; 
   reg __423914_423914;
   reg _423915_423915 ; 
   reg __423915_423915;
   reg _423916_423916 ; 
   reg __423916_423916;
   reg _423917_423917 ; 
   reg __423917_423917;
   reg _423918_423918 ; 
   reg __423918_423918;
   reg _423919_423919 ; 
   reg __423919_423919;
   reg _423920_423920 ; 
   reg __423920_423920;
   reg _423921_423921 ; 
   reg __423921_423921;
   reg _423922_423922 ; 
   reg __423922_423922;
   reg _423923_423923 ; 
   reg __423923_423923;
   reg _423924_423924 ; 
   reg __423924_423924;
   reg _423925_423925 ; 
   reg __423925_423925;
   reg _423926_423926 ; 
   reg __423926_423926;
   reg _423927_423927 ; 
   reg __423927_423927;
   reg _423928_423928 ; 
   reg __423928_423928;
   reg _423929_423929 ; 
   reg __423929_423929;
   reg _423930_423930 ; 
   reg __423930_423930;
   reg _423931_423931 ; 
   reg __423931_423931;
   reg _423932_423932 ; 
   reg __423932_423932;
   reg _423933_423933 ; 
   reg __423933_423933;
   reg _423934_423934 ; 
   reg __423934_423934;
   reg _423935_423935 ; 
   reg __423935_423935;
   reg _423936_423936 ; 
   reg __423936_423936;
   reg _423937_423937 ; 
   reg __423937_423937;
   reg _423938_423938 ; 
   reg __423938_423938;
   reg _423939_423939 ; 
   reg __423939_423939;
   reg _423940_423940 ; 
   reg __423940_423940;
   reg _423941_423941 ; 
   reg __423941_423941;
   reg _423942_423942 ; 
   reg __423942_423942;
   reg _423943_423943 ; 
   reg __423943_423943;
   reg _423944_423944 ; 
   reg __423944_423944;
   reg _423945_423945 ; 
   reg __423945_423945;
   reg _423946_423946 ; 
   reg __423946_423946;
   reg _423947_423947 ; 
   reg __423947_423947;
   reg _423948_423948 ; 
   reg __423948_423948;
   reg _423949_423949 ; 
   reg __423949_423949;
   reg _423950_423950 ; 
   reg __423950_423950;
   reg _423951_423951 ; 
   reg __423951_423951;
   reg _423952_423952 ; 
   reg __423952_423952;
   reg _423953_423953 ; 
   reg __423953_423953;
   reg _423954_423954 ; 
   reg __423954_423954;
   reg _423955_423955 ; 
   reg __423955_423955;
   reg _423956_423956 ; 
   reg __423956_423956;
   reg _423957_423957 ; 
   reg __423957_423957;
   reg _423958_423958 ; 
   reg __423958_423958;
   reg _423959_423959 ; 
   reg __423959_423959;
   reg _423960_423960 ; 
   reg __423960_423960;
   reg _423961_423961 ; 
   reg __423961_423961;
   reg _423962_423962 ; 
   reg __423962_423962;
   reg _423963_423963 ; 
   reg __423963_423963;
   reg _423964_423964 ; 
   reg __423964_423964;
   reg _423965_423965 ; 
   reg __423965_423965;
   reg _423966_423966 ; 
   reg __423966_423966;
   reg _423967_423967 ; 
   reg __423967_423967;
   reg _423968_423968 ; 
   reg __423968_423968;
   reg _423969_423969 ; 
   reg __423969_423969;
   reg _423970_423970 ; 
   reg __423970_423970;
   reg _423971_423971 ; 
   reg __423971_423971;
   reg _423972_423972 ; 
   reg __423972_423972;
   reg _423973_423973 ; 
   reg __423973_423973;
   reg _423974_423974 ; 
   reg __423974_423974;
   reg _423975_423975 ; 
   reg __423975_423975;
   reg _423976_423976 ; 
   reg __423976_423976;
   reg _423977_423977 ; 
   reg __423977_423977;
   reg _423978_423978 ; 
   reg __423978_423978;
   reg _423979_423979 ; 
   reg __423979_423979;
   reg _423980_423980 ; 
   reg __423980_423980;
   reg _423981_423981 ; 
   reg __423981_423981;
   reg _423982_423982 ; 
   reg __423982_423982;
   reg _423983_423983 ; 
   reg __423983_423983;
   reg _423984_423984 ; 
   reg __423984_423984;
   reg _423985_423985 ; 
   reg __423985_423985;
   reg _423986_423986 ; 
   reg __423986_423986;
   reg _423987_423987 ; 
   reg __423987_423987;
   reg _423988_423988 ; 
   reg __423988_423988;
   reg _423989_423989 ; 
   reg __423989_423989;
   reg _423990_423990 ; 
   reg __423990_423990;
   reg _423991_423991 ; 
   reg __423991_423991;
   reg _423992_423992 ; 
   reg __423992_423992;
   reg _423993_423993 ; 
   reg __423993_423993;
   reg _423994_423994 ; 
   reg __423994_423994;
   reg _423995_423995 ; 
   reg __423995_423995;
   reg _423996_423996 ; 
   reg __423996_423996;
   reg _423997_423997 ; 
   reg __423997_423997;
   reg _423998_423998 ; 
   reg __423998_423998;
   reg _423999_423999 ; 
   reg __423999_423999;
   reg _424000_424000 ; 
   reg __424000_424000;
   reg _424001_424001 ; 
   reg __424001_424001;
   reg _424002_424002 ; 
   reg __424002_424002;
   reg _424003_424003 ; 
   reg __424003_424003;
   reg _424004_424004 ; 
   reg __424004_424004;
   reg _424005_424005 ; 
   reg __424005_424005;
   reg _424006_424006 ; 
   reg __424006_424006;
   reg _424007_424007 ; 
   reg __424007_424007;
   reg _424008_424008 ; 
   reg __424008_424008;
   reg _424009_424009 ; 
   reg __424009_424009;
   reg _424010_424010 ; 
   reg __424010_424010;
   reg _424011_424011 ; 
   reg __424011_424011;
   reg _424012_424012 ; 
   reg __424012_424012;
   reg _424013_424013 ; 
   reg __424013_424013;
   reg _424014_424014 ; 
   reg __424014_424014;
   reg _424015_424015 ; 
   reg __424015_424015;
   reg _424016_424016 ; 
   reg __424016_424016;
   reg _424017_424017 ; 
   reg __424017_424017;
   reg _424018_424018 ; 
   reg __424018_424018;
   reg _424019_424019 ; 
   reg __424019_424019;
   reg _424020_424020 ; 
   reg __424020_424020;
   reg _424021_424021 ; 
   reg __424021_424021;
   reg _424022_424022 ; 
   reg __424022_424022;
   reg _424023_424023 ; 
   reg __424023_424023;
   reg _424024_424024 ; 
   reg __424024_424024;
   reg _424025_424025 ; 
   reg __424025_424025;
   reg _424026_424026 ; 
   reg __424026_424026;
   reg _424027_424027 ; 
   reg __424027_424027;
   reg _424028_424028 ; 
   reg __424028_424028;
   reg _424029_424029 ; 
   reg __424029_424029;
   reg _424030_424030 ; 
   reg __424030_424030;
   reg _424031_424031 ; 
   reg __424031_424031;
   reg _424032_424032 ; 
   reg __424032_424032;
   reg _424033_424033 ; 
   reg __424033_424033;
   reg _424034_424034 ; 
   reg __424034_424034;
   reg _424035_424035 ; 
   reg __424035_424035;
   reg _424036_424036 ; 
   reg __424036_424036;
   reg _424037_424037 ; 
   reg __424037_424037;
   reg _424038_424038 ; 
   reg __424038_424038;
   reg _424039_424039 ; 
   reg __424039_424039;
   reg _424040_424040 ; 
   reg __424040_424040;
   reg _424041_424041 ; 
   reg __424041_424041;
   reg _424042_424042 ; 
   reg __424042_424042;
   reg _424043_424043 ; 
   reg __424043_424043;
   reg _424044_424044 ; 
   reg __424044_424044;
   reg _424045_424045 ; 
   reg __424045_424045;
   reg _424046_424046 ; 
   reg __424046_424046;
   reg _424047_424047 ; 
   reg __424047_424047;
   reg _424048_424048 ; 
   reg __424048_424048;
   reg _424049_424049 ; 
   reg __424049_424049;
   reg _424050_424050 ; 
   reg __424050_424050;
   reg _424051_424051 ; 
   reg __424051_424051;
   reg _424052_424052 ; 
   reg __424052_424052;
   reg _424053_424053 ; 
   reg __424053_424053;
   reg _424054_424054 ; 
   reg __424054_424054;
   reg _424055_424055 ; 
   reg __424055_424055;
   reg _424056_424056 ; 
   reg __424056_424056;
   reg _424057_424057 ; 
   reg __424057_424057;
   reg _424058_424058 ; 
   reg __424058_424058;
   reg _424059_424059 ; 
   reg __424059_424059;
   reg _424060_424060 ; 
   reg __424060_424060;
   reg _424061_424061 ; 
   reg __424061_424061;
   reg _424062_424062 ; 
   reg __424062_424062;
   reg _424063_424063 ; 
   reg __424063_424063;
   reg _424064_424064 ; 
   reg __424064_424064;
   reg _424065_424065 ; 
   reg __424065_424065;
   reg _424066_424066 ; 
   reg __424066_424066;
   reg _424067_424067 ; 
   reg __424067_424067;
   reg _424068_424068 ; 
   reg __424068_424068;
   reg _424069_424069 ; 
   reg __424069_424069;
   reg _424070_424070 ; 
   reg __424070_424070;
   reg _424071_424071 ; 
   reg __424071_424071;
   reg _424072_424072 ; 
   reg __424072_424072;
   reg _424073_424073 ; 
   reg __424073_424073;
   reg _424074_424074 ; 
   reg __424074_424074;
   reg _424075_424075 ; 
   reg __424075_424075;
   reg _424076_424076 ; 
   reg __424076_424076;
   reg _424077_424077 ; 
   reg __424077_424077;
   reg _424078_424078 ; 
   reg __424078_424078;
   reg _424079_424079 ; 
   reg __424079_424079;
   reg _424080_424080 ; 
   reg __424080_424080;
   reg _424081_424081 ; 
   reg __424081_424081;
   reg _424082_424082 ; 
   reg __424082_424082;
   reg _424083_424083 ; 
   reg __424083_424083;
   reg _424084_424084 ; 
   reg __424084_424084;
   reg _424085_424085 ; 
   reg __424085_424085;
   reg _424086_424086 ; 
   reg __424086_424086;
   reg _424087_424087 ; 
   reg __424087_424087;
   reg _424088_424088 ; 
   reg __424088_424088;
   reg _424089_424089 ; 
   reg __424089_424089;
   reg _424090_424090 ; 
   reg __424090_424090;
   reg _424091_424091 ; 
   reg __424091_424091;
   reg _424092_424092 ; 
   reg __424092_424092;
   reg _424093_424093 ; 
   reg __424093_424093;
   reg _424094_424094 ; 
   reg __424094_424094;
   reg _424095_424095 ; 
   reg __424095_424095;
   reg _424096_424096 ; 
   reg __424096_424096;
   reg _424097_424097 ; 
   reg __424097_424097;
   reg _424098_424098 ; 
   reg __424098_424098;
   reg _424099_424099 ; 
   reg __424099_424099;
   reg _424100_424100 ; 
   reg __424100_424100;
   reg _424101_424101 ; 
   reg __424101_424101;
   reg _424102_424102 ; 
   reg __424102_424102;
   reg _424103_424103 ; 
   reg __424103_424103;
   reg _424104_424104 ; 
   reg __424104_424104;
   reg _424105_424105 ; 
   reg __424105_424105;
   reg _424106_424106 ; 
   reg __424106_424106;
   reg _424107_424107 ; 
   reg __424107_424107;
   reg _424108_424108 ; 
   reg __424108_424108;
   reg _424109_424109 ; 
   reg __424109_424109;
   reg _424110_424110 ; 
   reg __424110_424110;
   reg _424111_424111 ; 
   reg __424111_424111;
   reg _424112_424112 ; 
   reg __424112_424112;
   reg _424113_424113 ; 
   reg __424113_424113;
   reg _424114_424114 ; 
   reg __424114_424114;
   reg _424115_424115 ; 
   reg __424115_424115;
   reg _424116_424116 ; 
   reg __424116_424116;
   reg _424117_424117 ; 
   reg __424117_424117;
   reg _424118_424118 ; 
   reg __424118_424118;
   reg _424119_424119 ; 
   reg __424119_424119;
   reg _424120_424120 ; 
   reg __424120_424120;
   reg _424121_424121 ; 
   reg __424121_424121;
   reg _424122_424122 ; 
   reg __424122_424122;
   reg _424123_424123 ; 
   reg __424123_424123;
   reg _424124_424124 ; 
   reg __424124_424124;
   reg _424125_424125 ; 
   reg __424125_424125;
   reg _424126_424126 ; 
   reg __424126_424126;
   reg _424127_424127 ; 
   reg __424127_424127;
   reg _424128_424128 ; 
   reg __424128_424128;
   reg _424129_424129 ; 
   reg __424129_424129;
   reg _424130_424130 ; 
   reg __424130_424130;
   reg _424131_424131 ; 
   reg __424131_424131;
   reg _424132_424132 ; 
   reg __424132_424132;
   reg _424133_424133 ; 
   reg __424133_424133;
   reg _424134_424134 ; 
   reg __424134_424134;
   reg _424135_424135 ; 
   reg __424135_424135;
   reg _424136_424136 ; 
   reg __424136_424136;
   reg _424137_424137 ; 
   reg __424137_424137;
   reg _424138_424138 ; 
   reg __424138_424138;
   reg _424139_424139 ; 
   reg __424139_424139;
   reg _424140_424140 ; 
   reg __424140_424140;
   reg _424141_424141 ; 
   reg __424141_424141;
   reg _424142_424142 ; 
   reg __424142_424142;
   reg _424143_424143 ; 
   reg __424143_424143;
   reg _424144_424144 ; 
   reg __424144_424144;
   reg _424145_424145 ; 
   reg __424145_424145;
   reg _424146_424146 ; 
   reg __424146_424146;
   reg _424147_424147 ; 
   reg __424147_424147;
   reg _424148_424148 ; 
   reg __424148_424148;
   reg _424149_424149 ; 
   reg __424149_424149;
   reg _424150_424150 ; 
   reg __424150_424150;
   reg _424151_424151 ; 
   reg __424151_424151;
   reg _424152_424152 ; 
   reg __424152_424152;
   reg _424153_424153 ; 
   reg __424153_424153;
   reg _424154_424154 ; 
   reg __424154_424154;
   reg _424155_424155 ; 
   reg __424155_424155;
   reg _424156_424156 ; 
   reg __424156_424156;
   reg _424157_424157 ; 
   reg __424157_424157;
   reg _424158_424158 ; 
   reg __424158_424158;
   reg _424159_424159 ; 
   reg __424159_424159;
   reg _424160_424160 ; 
   reg __424160_424160;
   reg _424161_424161 ; 
   reg __424161_424161;
   reg _424162_424162 ; 
   reg __424162_424162;
   reg _424163_424163 ; 
   reg __424163_424163;
   reg _424164_424164 ; 
   reg __424164_424164;
   reg _424165_424165 ; 
   reg __424165_424165;
   reg _424166_424166 ; 
   reg __424166_424166;
   reg _424167_424167 ; 
   reg __424167_424167;
   reg _424168_424168 ; 
   reg __424168_424168;
   reg _424169_424169 ; 
   reg __424169_424169;
   reg _424170_424170 ; 
   reg __424170_424170;
   reg _424171_424171 ; 
   reg __424171_424171;
   reg _424172_424172 ; 
   reg __424172_424172;
   reg _424173_424173 ; 
   reg __424173_424173;
   reg _424174_424174 ; 
   reg __424174_424174;
   reg _424175_424175 ; 
   reg __424175_424175;
   reg _424176_424176 ; 
   reg __424176_424176;
   reg _424177_424177 ; 
   reg __424177_424177;
   reg _424178_424178 ; 
   reg __424178_424178;
   reg _424179_424179 ; 
   reg __424179_424179;
   reg _424180_424180 ; 
   reg __424180_424180;
   reg _424181_424181 ; 
   reg __424181_424181;
   reg _424182_424182 ; 
   reg __424182_424182;
   reg _424183_424183 ; 
   reg __424183_424183;
   reg _424184_424184 ; 
   reg __424184_424184;
   reg _424185_424185 ; 
   reg __424185_424185;
   reg _424186_424186 ; 
   reg __424186_424186;
   reg _424187_424187 ; 
   reg __424187_424187;
   reg _424188_424188 ; 
   reg __424188_424188;
   reg _424189_424189 ; 
   reg __424189_424189;
   reg _424190_424190 ; 
   reg __424190_424190;
   reg _424191_424191 ; 
   reg __424191_424191;
   reg _424192_424192 ; 
   reg __424192_424192;
   reg _424193_424193 ; 
   reg __424193_424193;
   reg _424194_424194 ; 
   reg __424194_424194;
   reg _424195_424195 ; 
   reg __424195_424195;
   reg _424196_424196 ; 
   reg __424196_424196;
   reg _424197_424197 ; 
   reg __424197_424197;
   reg _424198_424198 ; 
   reg __424198_424198;
   reg _424199_424199 ; 
   reg __424199_424199;
   reg _424200_424200 ; 
   reg __424200_424200;
   reg _424201_424201 ; 
   reg __424201_424201;
   reg _424202_424202 ; 
   reg __424202_424202;
   reg _424203_424203 ; 
   reg __424203_424203;
   reg _424204_424204 ; 
   reg __424204_424204;
   reg _424205_424205 ; 
   reg __424205_424205;
   reg _424206_424206 ; 
   reg __424206_424206;
   reg _424207_424207 ; 
   reg __424207_424207;
   reg _424208_424208 ; 
   reg __424208_424208;
   reg _424209_424209 ; 
   reg __424209_424209;
   reg _424210_424210 ; 
   reg __424210_424210;
   reg _424211_424211 ; 
   reg __424211_424211;
   reg _424212_424212 ; 
   reg __424212_424212;
   reg _424213_424213 ; 
   reg __424213_424213;
   reg _424214_424214 ; 
   reg __424214_424214;
   reg _424215_424215 ; 
   reg __424215_424215;
   reg _424216_424216 ; 
   reg __424216_424216;
   reg _424217_424217 ; 
   reg __424217_424217;
   reg _424218_424218 ; 
   reg __424218_424218;
   reg _424219_424219 ; 
   reg __424219_424219;
   reg _424220_424220 ; 
   reg __424220_424220;
   reg _424221_424221 ; 
   reg __424221_424221;
   reg _424222_424222 ; 
   reg __424222_424222;
   reg _424223_424223 ; 
   reg __424223_424223;
   reg _424224_424224 ; 
   reg __424224_424224;
   reg _424225_424225 ; 
   reg __424225_424225;
   reg _424226_424226 ; 
   reg __424226_424226;
   reg _424227_424227 ; 
   reg __424227_424227;
   reg _424228_424228 ; 
   reg __424228_424228;
   reg _424229_424229 ; 
   reg __424229_424229;
   reg _424230_424230 ; 
   reg __424230_424230;
   reg _424231_424231 ; 
   reg __424231_424231;
   reg _424232_424232 ; 
   reg __424232_424232;
   reg _424233_424233 ; 
   reg __424233_424233;
   reg _424234_424234 ; 
   reg __424234_424234;
   reg _424235_424235 ; 
   reg __424235_424235;
   reg _424236_424236 ; 
   reg __424236_424236;
   reg _424237_424237 ; 
   reg __424237_424237;
   reg _424238_424238 ; 
   reg __424238_424238;
   reg _424239_424239 ; 
   reg __424239_424239;
   reg _424240_424240 ; 
   reg __424240_424240;
   reg _424241_424241 ; 
   reg __424241_424241;
   reg _424242_424242 ; 
   reg __424242_424242;
   reg _424243_424243 ; 
   reg __424243_424243;
   reg _424244_424244 ; 
   reg __424244_424244;
   reg _424245_424245 ; 
   reg __424245_424245;
   reg _424246_424246 ; 
   reg __424246_424246;
   reg _424247_424247 ; 
   reg __424247_424247;
   reg _424248_424248 ; 
   reg __424248_424248;
   reg _424249_424249 ; 
   reg __424249_424249;
   reg _424250_424250 ; 
   reg __424250_424250;
   reg _424251_424251 ; 
   reg __424251_424251;
   reg _424252_424252 ; 
   reg __424252_424252;
   reg _424253_424253 ; 
   reg __424253_424253;
   reg _424254_424254 ; 
   reg __424254_424254;
   reg _424255_424255 ; 
   reg __424255_424255;
   reg _424256_424256 ; 
   reg __424256_424256;
   reg _424257_424257 ; 
   reg __424257_424257;
   reg _424258_424258 ; 
   reg __424258_424258;
   reg _424259_424259 ; 
   reg __424259_424259;
   reg _424260_424260 ; 
   reg __424260_424260;
   reg _424261_424261 ; 
   reg __424261_424261;
   reg _424262_424262 ; 
   reg __424262_424262;
   reg _424263_424263 ; 
   reg __424263_424263;
   reg _424264_424264 ; 
   reg __424264_424264;
   reg _424265_424265 ; 
   reg __424265_424265;
   reg _424266_424266 ; 
   reg __424266_424266;
   reg _424267_424267 ; 
   reg __424267_424267;
   reg _424268_424268 ; 
   reg __424268_424268;
   reg _424269_424269 ; 
   reg __424269_424269;
   reg _424270_424270 ; 
   reg __424270_424270;
   reg _424271_424271 ; 
   reg __424271_424271;
   reg _424272_424272 ; 
   reg __424272_424272;
   reg _424273_424273 ; 
   reg __424273_424273;
   reg _424274_424274 ; 
   reg __424274_424274;
   reg _424275_424275 ; 
   reg __424275_424275;
   reg _424276_424276 ; 
   reg __424276_424276;
   reg _424277_424277 ; 
   reg __424277_424277;
   reg _424278_424278 ; 
   reg __424278_424278;
   reg _424279_424279 ; 
   reg __424279_424279;
   reg _424280_424280 ; 
   reg __424280_424280;
   reg _424281_424281 ; 
   reg __424281_424281;
   reg _424282_424282 ; 
   reg __424282_424282;
   reg _424283_424283 ; 
   reg __424283_424283;
   reg _424284_424284 ; 
   reg __424284_424284;
   reg _424285_424285 ; 
   reg __424285_424285;
   reg _424286_424286 ; 
   reg __424286_424286;
   reg _424287_424287 ; 
   reg __424287_424287;
   reg _424288_424288 ; 
   reg __424288_424288;
   reg _424289_424289 ; 
   reg __424289_424289;
   reg _424290_424290 ; 
   reg __424290_424290;
   reg _424291_424291 ; 
   reg __424291_424291;
   reg _424292_424292 ; 
   reg __424292_424292;
   reg _424293_424293 ; 
   reg __424293_424293;
   reg _424294_424294 ; 
   reg __424294_424294;
   reg _424295_424295 ; 
   reg __424295_424295;
   reg _424296_424296 ; 
   reg __424296_424296;
   reg _424297_424297 ; 
   reg __424297_424297;
   reg _424298_424298 ; 
   reg __424298_424298;
   reg _424299_424299 ; 
   reg __424299_424299;
   reg _424300_424300 ; 
   reg __424300_424300;
   reg _424301_424301 ; 
   reg __424301_424301;
   reg _424302_424302 ; 
   reg __424302_424302;
   reg _424303_424303 ; 
   reg __424303_424303;
   reg _424304_424304 ; 
   reg __424304_424304;
   reg _424305_424305 ; 
   reg __424305_424305;
   reg _424306_424306 ; 
   reg __424306_424306;
   reg _424307_424307 ; 
   reg __424307_424307;
   reg _424308_424308 ; 
   reg __424308_424308;
   reg _424309_424309 ; 
   reg __424309_424309;
   reg _424310_424310 ; 
   reg __424310_424310;
   reg _424311_424311 ; 
   reg __424311_424311;
   reg _424312_424312 ; 
   reg __424312_424312;
   reg _424313_424313 ; 
   reg __424313_424313;
   reg _424314_424314 ; 
   reg __424314_424314;
   reg _424315_424315 ; 
   reg __424315_424315;
   reg _424316_424316 ; 
   reg __424316_424316;
   reg _424317_424317 ; 
   reg __424317_424317;
   reg _424318_424318 ; 
   reg __424318_424318;
   reg _424319_424319 ; 
   reg __424319_424319;
   reg _424320_424320 ; 
   reg __424320_424320;
   reg _424321_424321 ; 
   reg __424321_424321;
   reg _424322_424322 ; 
   reg __424322_424322;
   reg _424323_424323 ; 
   reg __424323_424323;
   reg _424324_424324 ; 
   reg __424324_424324;
   reg _424325_424325 ; 
   reg __424325_424325;
   reg _424326_424326 ; 
   reg __424326_424326;
   reg _424327_424327 ; 
   reg __424327_424327;
   reg _424328_424328 ; 
   reg __424328_424328;
   reg _424329_424329 ; 
   reg __424329_424329;
   reg _424330_424330 ; 
   reg __424330_424330;
   reg _424331_424331 ; 
   reg __424331_424331;
   reg _424332_424332 ; 
   reg __424332_424332;
   reg _424333_424333 ; 
   reg __424333_424333;
   reg _424334_424334 ; 
   reg __424334_424334;
   reg _424335_424335 ; 
   reg __424335_424335;
   reg _424336_424336 ; 
   reg __424336_424336;
   reg _424337_424337 ; 
   reg __424337_424337;
   reg _424338_424338 ; 
   reg __424338_424338;
   reg _424339_424339 ; 
   reg __424339_424339;
   reg _424340_424340 ; 
   reg __424340_424340;
   reg _424341_424341 ; 
   reg __424341_424341;
   reg _424342_424342 ; 
   reg __424342_424342;
   reg _424343_424343 ; 
   reg __424343_424343;
   reg _424344_424344 ; 
   reg __424344_424344;
   reg _424345_424345 ; 
   reg __424345_424345;
   reg _424346_424346 ; 
   reg __424346_424346;
   reg _424347_424347 ; 
   reg __424347_424347;
   reg _424348_424348 ; 
   reg __424348_424348;
   reg _424349_424349 ; 
   reg __424349_424349;
   reg _424350_424350 ; 
   reg __424350_424350;
   reg _424351_424351 ; 
   reg __424351_424351;
   reg _424352_424352 ; 
   reg __424352_424352;
   reg _424353_424353 ; 
   reg __424353_424353;
   reg _424354_424354 ; 
   reg __424354_424354;
   reg _424355_424355 ; 
   reg __424355_424355;
   reg _424356_424356 ; 
   reg __424356_424356;
   reg _424357_424357 ; 
   reg __424357_424357;
   reg _424358_424358 ; 
   reg __424358_424358;
   reg _424359_424359 ; 
   reg __424359_424359;
   reg _424360_424360 ; 
   reg __424360_424360;
   reg _424361_424361 ; 
   reg __424361_424361;
   reg _424362_424362 ; 
   reg __424362_424362;
   reg _424363_424363 ; 
   reg __424363_424363;
   reg _424364_424364 ; 
   reg __424364_424364;
   reg _424365_424365 ; 
   reg __424365_424365;
   reg _424366_424366 ; 
   reg __424366_424366;
   reg _424367_424367 ; 
   reg __424367_424367;
   reg _424368_424368 ; 
   reg __424368_424368;
   reg _424369_424369 ; 
   reg __424369_424369;
   reg _424370_424370 ; 
   reg __424370_424370;
   reg _424371_424371 ; 
   reg __424371_424371;
   reg _424372_424372 ; 
   reg __424372_424372;
   reg _424373_424373 ; 
   reg __424373_424373;
   reg _424374_424374 ; 
   reg __424374_424374;
   reg _424375_424375 ; 
   reg __424375_424375;
   reg _424376_424376 ; 
   reg __424376_424376;
   reg _424377_424377 ; 
   reg __424377_424377;
   reg _424378_424378 ; 
   reg __424378_424378;
   reg _424379_424379 ; 
   reg __424379_424379;
   reg _424380_424380 ; 
   reg __424380_424380;
   reg _424381_424381 ; 
   reg __424381_424381;
   reg _424382_424382 ; 
   reg __424382_424382;
   reg _424383_424383 ; 
   reg __424383_424383;
   reg _424384_424384 ; 
   reg __424384_424384;
   reg _424385_424385 ; 
   reg __424385_424385;
   reg _424386_424386 ; 
   reg __424386_424386;
   reg _424387_424387 ; 
   reg __424387_424387;
   reg _424388_424388 ; 
   reg __424388_424388;
   reg _424389_424389 ; 
   reg __424389_424389;
   reg _424390_424390 ; 
   reg __424390_424390;
   reg _424391_424391 ; 
   reg __424391_424391;
   reg _424392_424392 ; 
   reg __424392_424392;
   reg _424393_424393 ; 
   reg __424393_424393;
   reg _424394_424394 ; 
   reg __424394_424394;
   reg _424395_424395 ; 
   reg __424395_424395;
   reg _424396_424396 ; 
   reg __424396_424396;
   reg _424397_424397 ; 
   reg __424397_424397;
   reg _424398_424398 ; 
   reg __424398_424398;
   reg _424399_424399 ; 
   reg __424399_424399;
   reg _424400_424400 ; 
   reg __424400_424400;
   reg _424401_424401 ; 
   reg __424401_424401;
   reg _424402_424402 ; 
   reg __424402_424402;
   reg _424403_424403 ; 
   reg __424403_424403;
   reg _424404_424404 ; 
   reg __424404_424404;
   reg _424405_424405 ; 
   reg __424405_424405;
   reg _424406_424406 ; 
   reg __424406_424406;
   reg _424407_424407 ; 
   reg __424407_424407;
   reg _424408_424408 ; 
   reg __424408_424408;
   reg _424409_424409 ; 
   reg __424409_424409;
   reg _424410_424410 ; 
   reg __424410_424410;
   reg _424411_424411 ; 
   reg __424411_424411;
   reg _424412_424412 ; 
   reg __424412_424412;
   reg _424413_424413 ; 
   reg __424413_424413;
   reg _424414_424414 ; 
   reg __424414_424414;
   reg _424415_424415 ; 
   reg __424415_424415;
   reg _424416_424416 ; 
   reg __424416_424416;
   reg _424417_424417 ; 
   reg __424417_424417;
   reg _424418_424418 ; 
   reg __424418_424418;
   reg _424419_424419 ; 
   reg __424419_424419;
   reg _424420_424420 ; 
   reg __424420_424420;
   reg _424421_424421 ; 
   reg __424421_424421;
   reg _424422_424422 ; 
   reg __424422_424422;
   reg _424423_424423 ; 
   reg __424423_424423;
   reg _424424_424424 ; 
   reg __424424_424424;
   reg _424425_424425 ; 
   reg __424425_424425;
   reg _424426_424426 ; 
   reg __424426_424426;
   reg _424427_424427 ; 
   reg __424427_424427;
   reg _424428_424428 ; 
   reg __424428_424428;
   reg _424429_424429 ; 
   reg __424429_424429;
   reg _424430_424430 ; 
   reg __424430_424430;
   reg _424431_424431 ; 
   reg __424431_424431;
   reg _424432_424432 ; 
   reg __424432_424432;
   reg _424433_424433 ; 
   reg __424433_424433;
   reg _424434_424434 ; 
   reg __424434_424434;
   reg _424435_424435 ; 
   reg __424435_424435;
   reg _424436_424436 ; 
   reg __424436_424436;
   reg _424437_424437 ; 
   reg __424437_424437;
   reg _424438_424438 ; 
   reg __424438_424438;
   reg _424439_424439 ; 
   reg __424439_424439;
   reg _424440_424440 ; 
   reg __424440_424440;
   reg _424441_424441 ; 
   reg __424441_424441;
   reg _424442_424442 ; 
   reg __424442_424442;
   reg _424443_424443 ; 
   reg __424443_424443;
   reg _424444_424444 ; 
   reg __424444_424444;
   reg _424445_424445 ; 
   reg __424445_424445;
   reg _424446_424446 ; 
   reg __424446_424446;
   reg _424447_424447 ; 
   reg __424447_424447;
   reg _424448_424448 ; 
   reg __424448_424448;
   reg _424449_424449 ; 
   reg __424449_424449;
   reg _424450_424450 ; 
   reg __424450_424450;
   reg _424451_424451 ; 
   reg __424451_424451;
   reg _424452_424452 ; 
   reg __424452_424452;
   reg _424453_424453 ; 
   reg __424453_424453;
   reg _424454_424454 ; 
   reg __424454_424454;
   reg _424455_424455 ; 
   reg __424455_424455;
   reg _424456_424456 ; 
   reg __424456_424456;
   reg _424457_424457 ; 
   reg __424457_424457;
   reg _424458_424458 ; 
   reg __424458_424458;
   reg _424459_424459 ; 
   reg __424459_424459;
   reg _424460_424460 ; 
   reg __424460_424460;
   reg _424461_424461 ; 
   reg __424461_424461;
   reg _424462_424462 ; 
   reg __424462_424462;
   reg _424463_424463 ; 
   reg __424463_424463;
   reg _424464_424464 ; 
   reg __424464_424464;
   reg _424465_424465 ; 
   reg __424465_424465;
   reg _424466_424466 ; 
   reg __424466_424466;
   reg _424467_424467 ; 
   reg __424467_424467;
   reg _424468_424468 ; 
   reg __424468_424468;
   reg _424469_424469 ; 
   reg __424469_424469;
   reg _424470_424470 ; 
   reg __424470_424470;
   reg _424471_424471 ; 
   reg __424471_424471;
   reg _424472_424472 ; 
   reg __424472_424472;
   reg _424473_424473 ; 
   reg __424473_424473;
   reg _424474_424474 ; 
   reg __424474_424474;
   reg _424475_424475 ; 
   reg __424475_424475;
   reg _424476_424476 ; 
   reg __424476_424476;
   reg _424477_424477 ; 
   reg __424477_424477;
   reg _424478_424478 ; 
   reg __424478_424478;
   reg _424479_424479 ; 
   reg __424479_424479;
   reg _424480_424480 ; 
   reg __424480_424480;
   reg _424481_424481 ; 
   reg __424481_424481;
   reg _424482_424482 ; 
   reg __424482_424482;
   reg _424483_424483 ; 
   reg __424483_424483;
   reg _424484_424484 ; 
   reg __424484_424484;
   reg _424485_424485 ; 
   reg __424485_424485;
   reg _424486_424486 ; 
   reg __424486_424486;
   reg _424487_424487 ; 
   reg __424487_424487;
   reg _424488_424488 ; 
   reg __424488_424488;
   reg _424489_424489 ; 
   reg __424489_424489;
   reg _424490_424490 ; 
   reg __424490_424490;
   reg _424491_424491 ; 
   reg __424491_424491;
   reg _424492_424492 ; 
   reg __424492_424492;
   reg _424493_424493 ; 
   reg __424493_424493;
   reg _424494_424494 ; 
   reg __424494_424494;
   reg _424495_424495 ; 
   reg __424495_424495;
   reg _424496_424496 ; 
   reg __424496_424496;
   reg _424497_424497 ; 
   reg __424497_424497;
   reg _424498_424498 ; 
   reg __424498_424498;
   reg _424499_424499 ; 
   reg __424499_424499;
   reg _424500_424500 ; 
   reg __424500_424500;
   reg _424501_424501 ; 
   reg __424501_424501;
   reg _424502_424502 ; 
   reg __424502_424502;
   reg _424503_424503 ; 
   reg __424503_424503;
   reg _424504_424504 ; 
   reg __424504_424504;
   reg _424505_424505 ; 
   reg __424505_424505;
   reg _424506_424506 ; 
   reg __424506_424506;
   reg _424507_424507 ; 
   reg __424507_424507;
   reg _424508_424508 ; 
   reg __424508_424508;
   reg _424509_424509 ; 
   reg __424509_424509;
   reg _424510_424510 ; 
   reg __424510_424510;
   reg _424511_424511 ; 
   reg __424511_424511;
   reg _424512_424512 ; 
   reg __424512_424512;
   reg _424513_424513 ; 
   reg __424513_424513;
   reg _424514_424514 ; 
   reg __424514_424514;
   reg _424515_424515 ; 
   reg __424515_424515;
   reg _424516_424516 ; 
   reg __424516_424516;
   reg _424517_424517 ; 
   reg __424517_424517;
   reg _424518_424518 ; 
   reg __424518_424518;
   reg _424519_424519 ; 
   reg __424519_424519;
   reg _424520_424520 ; 
   reg __424520_424520;
   reg _424521_424521 ; 
   reg __424521_424521;
   reg _424522_424522 ; 
   reg __424522_424522;
   reg _424523_424523 ; 
   reg __424523_424523;
   reg _424524_424524 ; 
   reg __424524_424524;
   reg _424525_424525 ; 
   reg __424525_424525;
   reg _424526_424526 ; 
   reg __424526_424526;
   reg _424527_424527 ; 
   reg __424527_424527;
   reg _424528_424528 ; 
   reg __424528_424528;
   reg _424529_424529 ; 
   reg __424529_424529;
   reg _424530_424530 ; 
   reg __424530_424530;
   reg _424531_424531 ; 
   reg __424531_424531;
   reg _424532_424532 ; 
   reg __424532_424532;
   reg _424533_424533 ; 
   reg __424533_424533;
   reg _424534_424534 ; 
   reg __424534_424534;
   reg _424535_424535 ; 
   reg __424535_424535;
   reg _424536_424536 ; 
   reg __424536_424536;
   reg _424537_424537 ; 
   reg __424537_424537;
   reg _424538_424538 ; 
   reg __424538_424538;
   reg _424539_424539 ; 
   reg __424539_424539;
   reg _424540_424540 ; 
   reg __424540_424540;
   reg _424541_424541 ; 
   reg __424541_424541;
   reg _424542_424542 ; 
   reg __424542_424542;
   reg _424543_424543 ; 
   reg __424543_424543;
   reg _424544_424544 ; 
   reg __424544_424544;
   reg _424545_424545 ; 
   reg __424545_424545;
   reg _424546_424546 ; 
   reg __424546_424546;
   reg _424547_424547 ; 
   reg __424547_424547;
   reg _424548_424548 ; 
   reg __424548_424548;
   reg _424549_424549 ; 
   reg __424549_424549;
   reg _424550_424550 ; 
   reg __424550_424550;
   reg _424551_424551 ; 
   reg __424551_424551;
   reg _424552_424552 ; 
   reg __424552_424552;
   reg _424553_424553 ; 
   reg __424553_424553;
   reg _424554_424554 ; 
   reg __424554_424554;
   reg _424555_424555 ; 
   reg __424555_424555;
   reg _424556_424556 ; 
   reg __424556_424556;
   reg _424557_424557 ; 
   reg __424557_424557;
   reg _424558_424558 ; 
   reg __424558_424558;
   reg _424559_424559 ; 
   reg __424559_424559;
   reg _424560_424560 ; 
   reg __424560_424560;
   reg _424561_424561 ; 
   reg __424561_424561;
   reg _424562_424562 ; 
   reg __424562_424562;
   reg _424563_424563 ; 
   reg __424563_424563;
   reg _424564_424564 ; 
   reg __424564_424564;
   reg _424565_424565 ; 
   reg __424565_424565;
   reg _424566_424566 ; 
   reg __424566_424566;
   reg _424567_424567 ; 
   reg __424567_424567;
   reg _424568_424568 ; 
   reg __424568_424568;
   reg _424569_424569 ; 
   reg __424569_424569;
   reg _424570_424570 ; 
   reg __424570_424570;
   reg _424571_424571 ; 
   reg __424571_424571;
   reg _424572_424572 ; 
   reg __424572_424572;
   reg _424573_424573 ; 
   reg __424573_424573;
   reg _424574_424574 ; 
   reg __424574_424574;
   reg _424575_424575 ; 
   reg __424575_424575;
   reg _424576_424576 ; 
   reg __424576_424576;
   reg _424577_424577 ; 
   reg __424577_424577;
   reg _424578_424578 ; 
   reg __424578_424578;
   reg _424579_424579 ; 
   reg __424579_424579;
   reg _424580_424580 ; 
   reg __424580_424580;
   reg _424581_424581 ; 
   reg __424581_424581;
   reg _424582_424582 ; 
   reg __424582_424582;
   reg _424583_424583 ; 
   reg __424583_424583;
   reg _424584_424584 ; 
   reg __424584_424584;
   reg _424585_424585 ; 
   reg __424585_424585;
   reg _424586_424586 ; 
   reg __424586_424586;
   reg _424587_424587 ; 
   reg __424587_424587;
   reg _424588_424588 ; 
   reg __424588_424588;
   reg _424589_424589 ; 
   reg __424589_424589;
   reg _424590_424590 ; 
   reg __424590_424590;
   reg _424591_424591 ; 
   reg __424591_424591;
   reg _424592_424592 ; 
   reg __424592_424592;
   reg _424593_424593 ; 
   reg __424593_424593;
   reg _424594_424594 ; 
   reg __424594_424594;
   reg _424595_424595 ; 
   reg __424595_424595;
   reg _424596_424596 ; 
   reg __424596_424596;
   reg _424597_424597 ; 
   reg __424597_424597;
   reg _424598_424598 ; 
   reg __424598_424598;
   reg _424599_424599 ; 
   reg __424599_424599;
   reg _424600_424600 ; 
   reg __424600_424600;
   reg _424601_424601 ; 
   reg __424601_424601;
   reg _424602_424602 ; 
   reg __424602_424602;
   reg _424603_424603 ; 
   reg __424603_424603;
   reg _424604_424604 ; 
   reg __424604_424604;
   reg _424605_424605 ; 
   reg __424605_424605;
   reg _424606_424606 ; 
   reg __424606_424606;
   reg _424607_424607 ; 
   reg __424607_424607;
   reg _424608_424608 ; 
   reg __424608_424608;
   reg _424609_424609 ; 
   reg __424609_424609;
   reg _424610_424610 ; 
   reg __424610_424610;
   reg _424611_424611 ; 
   reg __424611_424611;
   reg _424612_424612 ; 
   reg __424612_424612;
   reg _424613_424613 ; 
   reg __424613_424613;
   reg _424614_424614 ; 
   reg __424614_424614;
   reg _424615_424615 ; 
   reg __424615_424615;
   reg _424616_424616 ; 
   reg __424616_424616;
   reg _424617_424617 ; 
   reg __424617_424617;
   reg _424618_424618 ; 
   reg __424618_424618;
   reg _424619_424619 ; 
   reg __424619_424619;
   reg _424620_424620 ; 
   reg __424620_424620;
   reg _424621_424621 ; 
   reg __424621_424621;
   reg _424622_424622 ; 
   reg __424622_424622;
   reg _424623_424623 ; 
   reg __424623_424623;
   reg _424624_424624 ; 
   reg __424624_424624;
   reg _424625_424625 ; 
   reg __424625_424625;
   reg _424626_424626 ; 
   reg __424626_424626;
   reg _424627_424627 ; 
   reg __424627_424627;
   reg _424628_424628 ; 
   reg __424628_424628;
   reg _424629_424629 ; 
   reg __424629_424629;
   reg _424630_424630 ; 
   reg __424630_424630;
   reg _424631_424631 ; 
   reg __424631_424631;
   reg _424632_424632 ; 
   reg __424632_424632;
   reg _424633_424633 ; 
   reg __424633_424633;
   reg _424634_424634 ; 
   reg __424634_424634;
   reg _424635_424635 ; 
   reg __424635_424635;
   reg _424636_424636 ; 
   reg __424636_424636;
   reg _424637_424637 ; 
   reg __424637_424637;
   reg _424638_424638 ; 
   reg __424638_424638;
   reg _424639_424639 ; 
   reg __424639_424639;
   reg _424640_424640 ; 
   reg __424640_424640;
   reg _424641_424641 ; 
   reg __424641_424641;
   reg _424642_424642 ; 
   reg __424642_424642;
   reg _424643_424643 ; 
   reg __424643_424643;
   reg _424644_424644 ; 
   reg __424644_424644;
   reg _424645_424645 ; 
   reg __424645_424645;
   reg _424646_424646 ; 
   reg __424646_424646;
   reg _424647_424647 ; 
   reg __424647_424647;
   reg _424648_424648 ; 
   reg __424648_424648;
   reg _424649_424649 ; 
   reg __424649_424649;
   reg _424650_424650 ; 
   reg __424650_424650;
   reg _424651_424651 ; 
   reg __424651_424651;
   reg _424652_424652 ; 
   reg __424652_424652;
   reg _424653_424653 ; 
   reg __424653_424653;
   reg _424654_424654 ; 
   reg __424654_424654;
   reg _424655_424655 ; 
   reg __424655_424655;
   reg _424656_424656 ; 
   reg __424656_424656;
   reg _424657_424657 ; 
   reg __424657_424657;
   reg _424658_424658 ; 
   reg __424658_424658;
   reg _424659_424659 ; 
   reg __424659_424659;
   reg _424660_424660 ; 
   reg __424660_424660;
   reg _424661_424661 ; 
   reg __424661_424661;
   reg _424662_424662 ; 
   reg __424662_424662;
   reg _424663_424663 ; 
   reg __424663_424663;
   reg _424664_424664 ; 
   reg __424664_424664;
   reg _424665_424665 ; 
   reg __424665_424665;
   reg _424666_424666 ; 
   reg __424666_424666;
   reg _424667_424667 ; 
   reg __424667_424667;
   reg _424668_424668 ; 
   reg __424668_424668;
   reg _424669_424669 ; 
   reg __424669_424669;
   reg _424670_424670 ; 
   reg __424670_424670;
   reg _424671_424671 ; 
   reg __424671_424671;
   reg _424672_424672 ; 
   reg __424672_424672;
   reg _424673_424673 ; 
   reg __424673_424673;
   reg _424674_424674 ; 
   reg __424674_424674;
   reg _424675_424675 ; 
   reg __424675_424675;
   reg _424676_424676 ; 
   reg __424676_424676;
   reg _424677_424677 ; 
   reg __424677_424677;
   reg _424678_424678 ; 
   reg __424678_424678;
   reg _424679_424679 ; 
   reg __424679_424679;
   reg _424680_424680 ; 
   reg __424680_424680;
   reg _424681_424681 ; 
   reg __424681_424681;
   reg _424682_424682 ; 
   reg __424682_424682;
   reg _424683_424683 ; 
   reg __424683_424683;
   reg _424684_424684 ; 
   reg __424684_424684;
   reg _424685_424685 ; 
   reg __424685_424685;
   reg _424686_424686 ; 
   reg __424686_424686;
   reg _424687_424687 ; 
   reg __424687_424687;
   reg _424688_424688 ; 
   reg __424688_424688;
   reg _424689_424689 ; 
   reg __424689_424689;
   reg _424690_424690 ; 
   reg __424690_424690;
   reg _424691_424691 ; 
   reg __424691_424691;
   reg _424692_424692 ; 
   reg __424692_424692;
   reg _424693_424693 ; 
   reg __424693_424693;
   reg _424694_424694 ; 
   reg __424694_424694;
   reg _424695_424695 ; 
   reg __424695_424695;
   reg _424696_424696 ; 
   reg __424696_424696;
   reg _424697_424697 ; 
   reg __424697_424697;
   reg _424698_424698 ; 
   reg __424698_424698;
   reg _424699_424699 ; 
   reg __424699_424699;
   reg _424700_424700 ; 
   reg __424700_424700;
   reg _424701_424701 ; 
   reg __424701_424701;
   reg _424702_424702 ; 
   reg __424702_424702;
   reg _424703_424703 ; 
   reg __424703_424703;
   reg _424704_424704 ; 
   reg __424704_424704;
   reg _424705_424705 ; 
   reg __424705_424705;
   reg _424706_424706 ; 
   reg __424706_424706;
   reg _424707_424707 ; 
   reg __424707_424707;
   reg _424708_424708 ; 
   reg __424708_424708;
   reg _424709_424709 ; 
   reg __424709_424709;
   reg _424710_424710 ; 
   reg __424710_424710;
   reg _424711_424711 ; 
   reg __424711_424711;
   reg _424712_424712 ; 
   reg __424712_424712;
   reg _424713_424713 ; 
   reg __424713_424713;
   reg _424714_424714 ; 
   reg __424714_424714;
   reg _424715_424715 ; 
   reg __424715_424715;
   reg _424716_424716 ; 
   reg __424716_424716;
   reg _424717_424717 ; 
   reg __424717_424717;
   reg _424718_424718 ; 
   reg __424718_424718;
   reg _424719_424719 ; 
   reg __424719_424719;
   reg _424720_424720 ; 
   reg __424720_424720;
   reg _424721_424721 ; 
   reg __424721_424721;
   reg _424722_424722 ; 
   reg __424722_424722;
   reg _424723_424723 ; 
   reg __424723_424723;
   reg _424724_424724 ; 
   reg __424724_424724;
   reg _424725_424725 ; 
   reg __424725_424725;
   reg _424726_424726 ; 
   reg __424726_424726;
   reg _424727_424727 ; 
   reg __424727_424727;
   reg _424728_424728 ; 
   reg __424728_424728;
   reg _424729_424729 ; 
   reg __424729_424729;
   reg _424730_424730 ; 
   reg __424730_424730;
   reg _424731_424731 ; 
   reg __424731_424731;
   reg _424732_424732 ; 
   reg __424732_424732;
   reg _424733_424733 ; 
   reg __424733_424733;
   reg _424734_424734 ; 
   reg __424734_424734;
   reg _424735_424735 ; 
   reg __424735_424735;
   reg _424736_424736 ; 
   reg __424736_424736;
   reg _424737_424737 ; 
   reg __424737_424737;
   reg _424738_424738 ; 
   reg __424738_424738;
   reg _424739_424739 ; 
   reg __424739_424739;
   reg _424740_424740 ; 
   reg __424740_424740;
   reg _424741_424741 ; 
   reg __424741_424741;
   reg _424742_424742 ; 
   reg __424742_424742;
   reg _424743_424743 ; 
   reg __424743_424743;
   reg _424744_424744 ; 
   reg __424744_424744;
   reg _424745_424745 ; 
   reg __424745_424745;
   reg _424746_424746 ; 
   reg __424746_424746;
   reg _424747_424747 ; 
   reg __424747_424747;
   reg _424748_424748 ; 
   reg __424748_424748;
   reg _424749_424749 ; 
   reg __424749_424749;
   reg _424750_424750 ; 
   reg __424750_424750;
   reg _424751_424751 ; 
   reg __424751_424751;
   reg _424752_424752 ; 
   reg __424752_424752;
   reg _424753_424753 ; 
   reg __424753_424753;
   reg _424754_424754 ; 
   reg __424754_424754;
   reg _424755_424755 ; 
   reg __424755_424755;
   reg _424756_424756 ; 
   reg __424756_424756;
   reg _424757_424757 ; 
   reg __424757_424757;
   reg _424758_424758 ; 
   reg __424758_424758;
   reg _424759_424759 ; 
   reg __424759_424759;
   reg _424760_424760 ; 
   reg __424760_424760;
   reg _424761_424761 ; 
   reg __424761_424761;
   reg _424762_424762 ; 
   reg __424762_424762;
   reg _424763_424763 ; 
   reg __424763_424763;
   reg _424764_424764 ; 
   reg __424764_424764;
   reg _424765_424765 ; 
   reg __424765_424765;
   reg _424766_424766 ; 
   reg __424766_424766;
   reg _424767_424767 ; 
   reg __424767_424767;
   reg _424768_424768 ; 
   reg __424768_424768;
   reg _424769_424769 ; 
   reg __424769_424769;
   reg _424770_424770 ; 
   reg __424770_424770;
   reg _424771_424771 ; 
   reg __424771_424771;
   reg _424772_424772 ; 
   reg __424772_424772;
   reg _424773_424773 ; 
   reg __424773_424773;
   reg _424774_424774 ; 
   reg __424774_424774;
   reg _424775_424775 ; 
   reg __424775_424775;
   reg _424776_424776 ; 
   reg __424776_424776;
   reg _424777_424777 ; 
   reg __424777_424777;
   reg _424778_424778 ; 
   reg __424778_424778;
   reg _424779_424779 ; 
   reg __424779_424779;
   reg _424780_424780 ; 
   reg __424780_424780;
   reg _424781_424781 ; 
   reg __424781_424781;
   reg _424782_424782 ; 
   reg __424782_424782;
   reg _424783_424783 ; 
   reg __424783_424783;
   reg _424784_424784 ; 
   reg __424784_424784;
   reg _424785_424785 ; 
   reg __424785_424785;
   reg _424786_424786 ; 
   reg __424786_424786;
   reg _424787_424787 ; 
   reg __424787_424787;
   reg _424788_424788 ; 
   reg __424788_424788;
   reg _424789_424789 ; 
   reg __424789_424789;
   reg _424790_424790 ; 
   reg __424790_424790;
   reg _424791_424791 ; 
   reg __424791_424791;
   reg _424792_424792 ; 
   reg __424792_424792;
   reg _424793_424793 ; 
   reg __424793_424793;
   reg _424794_424794 ; 
   reg __424794_424794;
   reg _424795_424795 ; 
   reg __424795_424795;
   reg _424796_424796 ; 
   reg __424796_424796;
   reg _424797_424797 ; 
   reg __424797_424797;
   reg _424798_424798 ; 
   reg __424798_424798;
   reg _424799_424799 ; 
   reg __424799_424799;
   reg _424800_424800 ; 
   reg __424800_424800;
   reg _424801_424801 ; 
   reg __424801_424801;
   reg _424802_424802 ; 
   reg __424802_424802;
   reg _424803_424803 ; 
   reg __424803_424803;
   reg _424804_424804 ; 
   reg __424804_424804;
   reg _424805_424805 ; 
   reg __424805_424805;
   reg _424806_424806 ; 
   reg __424806_424806;
   reg _424807_424807 ; 
   reg __424807_424807;
   reg _424808_424808 ; 
   reg __424808_424808;
   reg _424809_424809 ; 
   reg __424809_424809;
   reg _424810_424810 ; 
   reg __424810_424810;
   reg _424811_424811 ; 
   reg __424811_424811;
   reg _424812_424812 ; 
   reg __424812_424812;
   reg _424813_424813 ; 
   reg __424813_424813;
   reg _424814_424814 ; 
   reg __424814_424814;
   reg _424815_424815 ; 
   reg __424815_424815;
   reg _424816_424816 ; 
   reg __424816_424816;
   reg _424817_424817 ; 
   reg __424817_424817;
   reg _424818_424818 ; 
   reg __424818_424818;
   reg _424819_424819 ; 
   reg __424819_424819;
   reg _424820_424820 ; 
   reg __424820_424820;
   reg _424821_424821 ; 
   reg __424821_424821;
   reg _424822_424822 ; 
   reg __424822_424822;
   reg _424823_424823 ; 
   reg __424823_424823;
   reg _424824_424824 ; 
   reg __424824_424824;
   reg _424825_424825 ; 
   reg __424825_424825;
   reg _424826_424826 ; 
   reg __424826_424826;
   reg _424827_424827 ; 
   reg __424827_424827;
   reg _424828_424828 ; 
   reg __424828_424828;
   reg _424829_424829 ; 
   reg __424829_424829;
   reg _424830_424830 ; 
   reg __424830_424830;
   reg _424831_424831 ; 
   reg __424831_424831;
   reg _424832_424832 ; 
   reg __424832_424832;
   reg _424833_424833 ; 
   reg __424833_424833;
   reg _424834_424834 ; 
   reg __424834_424834;
   reg _424835_424835 ; 
   reg __424835_424835;
   reg _424836_424836 ; 
   reg __424836_424836;
   reg _424837_424837 ; 
   reg __424837_424837;
   reg _424838_424838 ; 
   reg __424838_424838;
   reg _424839_424839 ; 
   reg __424839_424839;
   reg _424840_424840 ; 
   reg __424840_424840;
   reg _424841_424841 ; 
   reg __424841_424841;
   reg _424842_424842 ; 
   reg __424842_424842;
   reg _424843_424843 ; 
   reg __424843_424843;
   reg _424844_424844 ; 
   reg __424844_424844;
   reg _424845_424845 ; 
   reg __424845_424845;
   reg _424846_424846 ; 
   reg __424846_424846;
   reg _424847_424847 ; 
   reg __424847_424847;
   reg _424848_424848 ; 
   reg __424848_424848;
   reg _424849_424849 ; 
   reg __424849_424849;
   reg _424850_424850 ; 
   reg __424850_424850;
   reg _424851_424851 ; 
   reg __424851_424851;
   reg _424852_424852 ; 
   reg __424852_424852;
   reg _424853_424853 ; 
   reg __424853_424853;
   reg _424854_424854 ; 
   reg __424854_424854;
   reg _424855_424855 ; 
   reg __424855_424855;
   reg _424856_424856 ; 
   reg __424856_424856;
   reg _424857_424857 ; 
   reg __424857_424857;
   reg _424858_424858 ; 
   reg __424858_424858;
   reg _424859_424859 ; 
   reg __424859_424859;
   reg _424860_424860 ; 
   reg __424860_424860;
   reg _424861_424861 ; 
   reg __424861_424861;
   reg _424862_424862 ; 
   reg __424862_424862;
   reg _424863_424863 ; 
   reg __424863_424863;
   reg _424864_424864 ; 
   reg __424864_424864;
   reg _424865_424865 ; 
   reg __424865_424865;
   reg _424866_424866 ; 
   reg __424866_424866;
   reg _424867_424867 ; 
   reg __424867_424867;
   reg _424868_424868 ; 
   reg __424868_424868;
   reg _424869_424869 ; 
   reg __424869_424869;
   reg _424870_424870 ; 
   reg __424870_424870;
   reg _424871_424871 ; 
   reg __424871_424871;
   reg _424872_424872 ; 
   reg __424872_424872;
   reg _424873_424873 ; 
   reg __424873_424873;
   reg _424874_424874 ; 
   reg __424874_424874;
   reg _424875_424875 ; 
   reg __424875_424875;
   reg _424876_424876 ; 
   reg __424876_424876;
   reg _424877_424877 ; 
   reg __424877_424877;
   reg _424878_424878 ; 
   reg __424878_424878;
   reg _424879_424879 ; 
   reg __424879_424879;
   reg _424880_424880 ; 
   reg __424880_424880;
   reg _424881_424881 ; 
   reg __424881_424881;
   reg _424882_424882 ; 
   reg __424882_424882;
   reg _424883_424883 ; 
   reg __424883_424883;
   reg _424884_424884 ; 
   reg __424884_424884;
   reg _424885_424885 ; 
   reg __424885_424885;
   reg _424886_424886 ; 
   reg __424886_424886;
   reg _424887_424887 ; 
   reg __424887_424887;
   reg _424888_424888 ; 
   reg __424888_424888;
   reg _424889_424889 ; 
   reg __424889_424889;
   reg _424890_424890 ; 
   reg __424890_424890;
   reg _424891_424891 ; 
   reg __424891_424891;
   reg _424892_424892 ; 
   reg __424892_424892;
   reg _424893_424893 ; 
   reg __424893_424893;
   reg _424894_424894 ; 
   reg __424894_424894;
   reg _424895_424895 ; 
   reg __424895_424895;
   reg _424896_424896 ; 
   reg __424896_424896;
   reg _424897_424897 ; 
   reg __424897_424897;
   reg _424898_424898 ; 
   reg __424898_424898;
   reg _424899_424899 ; 
   reg __424899_424899;
   reg _424900_424900 ; 
   reg __424900_424900;
   reg _424901_424901 ; 
   reg __424901_424901;
   reg _424902_424902 ; 
   reg __424902_424902;
   reg _424903_424903 ; 
   reg __424903_424903;
   reg _424904_424904 ; 
   reg __424904_424904;
   reg _424905_424905 ; 
   reg __424905_424905;
   reg _424906_424906 ; 
   reg __424906_424906;
   reg _424907_424907 ; 
   reg __424907_424907;
   reg _424908_424908 ; 
   reg __424908_424908;
   reg _424909_424909 ; 
   reg __424909_424909;
   reg _424910_424910 ; 
   reg __424910_424910;
   reg _424911_424911 ; 
   reg __424911_424911;
   reg _424912_424912 ; 
   reg __424912_424912;
   reg _424913_424913 ; 
   reg __424913_424913;
   reg _424914_424914 ; 
   reg __424914_424914;
   reg _424915_424915 ; 
   reg __424915_424915;
   reg _424916_424916 ; 
   reg __424916_424916;
   reg _424917_424917 ; 
   reg __424917_424917;
   reg _424918_424918 ; 
   reg __424918_424918;
   reg _424919_424919 ; 
   reg __424919_424919;
   reg _424920_424920 ; 
   reg __424920_424920;
   reg _424921_424921 ; 
   reg __424921_424921;
   reg _424922_424922 ; 
   reg __424922_424922;
   reg _424923_424923 ; 
   reg __424923_424923;
   reg _424924_424924 ; 
   reg __424924_424924;
   reg _424925_424925 ; 
   reg __424925_424925;
   reg _424926_424926 ; 
   reg __424926_424926;
   reg _424927_424927 ; 
   reg __424927_424927;
   reg _424928_424928 ; 
   reg __424928_424928;
   reg _424929_424929 ; 
   reg __424929_424929;
   reg _424930_424930 ; 
   reg __424930_424930;
   reg _424931_424931 ; 
   reg __424931_424931;
   reg _424932_424932 ; 
   reg __424932_424932;
   reg _424933_424933 ; 
   reg __424933_424933;
   reg _424934_424934 ; 
   reg __424934_424934;
   reg _424935_424935 ; 
   reg __424935_424935;
   reg _424936_424936 ; 
   reg __424936_424936;
   reg _424937_424937 ; 
   reg __424937_424937;
   reg _424938_424938 ; 
   reg __424938_424938;
   reg _424939_424939 ; 
   reg __424939_424939;
   reg _424940_424940 ; 
   reg __424940_424940;
   reg _424941_424941 ; 
   reg __424941_424941;
   reg _424942_424942 ; 
   reg __424942_424942;
   reg _424943_424943 ; 
   reg __424943_424943;
   reg _424944_424944 ; 
   reg __424944_424944;
   reg _424945_424945 ; 
   reg __424945_424945;
   reg _424946_424946 ; 
   reg __424946_424946;
   reg _424947_424947 ; 
   reg __424947_424947;
   reg _424948_424948 ; 
   reg __424948_424948;
   reg _424949_424949 ; 
   reg __424949_424949;
   reg _424950_424950 ; 
   reg __424950_424950;
   reg _424951_424951 ; 
   reg __424951_424951;
   reg _424952_424952 ; 
   reg __424952_424952;
   reg _424953_424953 ; 
   reg __424953_424953;
   reg _424954_424954 ; 
   reg __424954_424954;
   reg _424955_424955 ; 
   reg __424955_424955;
   reg _424956_424956 ; 
   reg __424956_424956;
   reg _424957_424957 ; 
   reg __424957_424957;
   reg _424958_424958 ; 
   reg __424958_424958;
   reg _424959_424959 ; 
   reg __424959_424959;
   reg _424960_424960 ; 
   reg __424960_424960;
   reg _424961_424961 ; 
   reg __424961_424961;
   reg _424962_424962 ; 
   reg __424962_424962;
   reg _424963_424963 ; 
   reg __424963_424963;
   reg _424964_424964 ; 
   reg __424964_424964;
   reg _424965_424965 ; 
   reg __424965_424965;
   reg _424966_424966 ; 
   reg __424966_424966;
   reg _424967_424967 ; 
   reg __424967_424967;
   reg _424968_424968 ; 
   reg __424968_424968;
   reg _424969_424969 ; 
   reg __424969_424969;
   reg _424970_424970 ; 
   reg __424970_424970;
   reg _424971_424971 ; 
   reg __424971_424971;
   reg _424972_424972 ; 
   reg __424972_424972;
   reg _424973_424973 ; 
   reg __424973_424973;
   reg _424974_424974 ; 
   reg __424974_424974;
   reg _424975_424975 ; 
   reg __424975_424975;
   reg _424976_424976 ; 
   reg __424976_424976;
   reg _424977_424977 ; 
   reg __424977_424977;
   reg _424978_424978 ; 
   reg __424978_424978;
   reg _424979_424979 ; 
   reg __424979_424979;
   reg _424980_424980 ; 
   reg __424980_424980;
   reg _424981_424981 ; 
   reg __424981_424981;
   reg _424982_424982 ; 
   reg __424982_424982;
   reg _424983_424983 ; 
   reg __424983_424983;
   reg _424984_424984 ; 
   reg __424984_424984;
   reg _424985_424985 ; 
   reg __424985_424985;
   reg _424986_424986 ; 
   reg __424986_424986;
   reg _424987_424987 ; 
   reg __424987_424987;
   reg _424988_424988 ; 
   reg __424988_424988;
   reg _424989_424989 ; 
   reg __424989_424989;
   reg _424990_424990 ; 
   reg __424990_424990;
   reg _424991_424991 ; 
   reg __424991_424991;
   reg _424992_424992 ; 
   reg __424992_424992;
   reg _424993_424993 ; 
   reg __424993_424993;
   reg _424994_424994 ; 
   reg __424994_424994;
   reg _424995_424995 ; 
   reg __424995_424995;
   reg _424996_424996 ; 
   reg __424996_424996;
   reg _424997_424997 ; 
   reg __424997_424997;
   reg _424998_424998 ; 
   reg __424998_424998;
   reg _424999_424999 ; 
   reg __424999_424999;
   reg _425000_425000 ; 
   reg __425000_425000;
   reg _425001_425001 ; 
   reg __425001_425001;
   reg _425002_425002 ; 
   reg __425002_425002;
   reg _425003_425003 ; 
   reg __425003_425003;
   reg _425004_425004 ; 
   reg __425004_425004;
   reg _425005_425005 ; 
   reg __425005_425005;
   reg _425006_425006 ; 
   reg __425006_425006;
   reg _425007_425007 ; 
   reg __425007_425007;
   reg _425008_425008 ; 
   reg __425008_425008;
   reg _425009_425009 ; 
   reg __425009_425009;
   reg _425010_425010 ; 
   reg __425010_425010;
   reg _425011_425011 ; 
   reg __425011_425011;
   reg _425012_425012 ; 
   reg __425012_425012;
   reg _425013_425013 ; 
   reg __425013_425013;
   reg _425014_425014 ; 
   reg __425014_425014;
   reg _425015_425015 ; 
   reg __425015_425015;
   reg _425016_425016 ; 
   reg __425016_425016;
   reg _425017_425017 ; 
   reg __425017_425017;
   reg _425018_425018 ; 
   reg __425018_425018;
   reg _425019_425019 ; 
   reg __425019_425019;
   reg _425020_425020 ; 
   reg __425020_425020;
   reg _425021_425021 ; 
   reg __425021_425021;
   reg _425022_425022 ; 
   reg __425022_425022;
   reg _425023_425023 ; 
   reg __425023_425023;
   reg _425024_425024 ; 
   reg __425024_425024;
   reg _425025_425025 ; 
   reg __425025_425025;
   reg _425026_425026 ; 
   reg __425026_425026;
   reg _425027_425027 ; 
   reg __425027_425027;
   reg _425028_425028 ; 
   reg __425028_425028;
   reg _425029_425029 ; 
   reg __425029_425029;
   reg _425030_425030 ; 
   reg __425030_425030;
   reg _425031_425031 ; 
   reg __425031_425031;
   reg _425032_425032 ; 
   reg __425032_425032;
   reg _425033_425033 ; 
   reg __425033_425033;
   reg _425034_425034 ; 
   reg __425034_425034;
   reg _425035_425035 ; 
   reg __425035_425035;
   reg _425036_425036 ; 
   reg __425036_425036;
   reg _425037_425037 ; 
   reg __425037_425037;
   reg _425038_425038 ; 
   reg __425038_425038;
   reg _425039_425039 ; 
   reg __425039_425039;
   reg _425040_425040 ; 
   reg __425040_425040;
   reg _425041_425041 ; 
   reg __425041_425041;
   reg _425042_425042 ; 
   reg __425042_425042;
   reg _425043_425043 ; 
   reg __425043_425043;
   reg _425044_425044 ; 
   reg __425044_425044;
   reg _425045_425045 ; 
   reg __425045_425045;
   reg _425046_425046 ; 
   reg __425046_425046;
   reg _425047_425047 ; 
   reg __425047_425047;
   reg _425048_425048 ; 
   reg __425048_425048;
   reg _425049_425049 ; 
   reg __425049_425049;
   reg _425050_425050 ; 
   reg __425050_425050;
   reg _425051_425051 ; 
   reg __425051_425051;
   reg _425052_425052 ; 
   reg __425052_425052;
   reg _425053_425053 ; 
   reg __425053_425053;
   reg _425054_425054 ; 
   reg __425054_425054;
   reg _425055_425055 ; 
   reg __425055_425055;
   reg _425056_425056 ; 
   reg __425056_425056;
   reg _425057_425057 ; 
   reg __425057_425057;
   reg _425058_425058 ; 
   reg __425058_425058;
   reg _425059_425059 ; 
   reg __425059_425059;
   reg _425060_425060 ; 
   reg __425060_425060;
   reg _425061_425061 ; 
   reg __425061_425061;
   reg _425062_425062 ; 
   reg __425062_425062;
   reg _425063_425063 ; 
   reg __425063_425063;
   reg _425064_425064 ; 
   reg __425064_425064;
   reg _425065_425065 ; 
   reg __425065_425065;
   reg _425066_425066 ; 
   reg __425066_425066;
   reg _425067_425067 ; 
   reg __425067_425067;
   reg _425068_425068 ; 
   reg __425068_425068;
   reg _425069_425069 ; 
   reg __425069_425069;
   reg _425070_425070 ; 
   reg __425070_425070;
   reg _425071_425071 ; 
   reg __425071_425071;
   reg _425072_425072 ; 
   reg __425072_425072;
   reg _425073_425073 ; 
   reg __425073_425073;
   reg _425074_425074 ; 
   reg __425074_425074;
   reg _425075_425075 ; 
   reg __425075_425075;
   reg _425076_425076 ; 
   reg __425076_425076;
   reg _425077_425077 ; 
   reg __425077_425077;
   reg _425078_425078 ; 
   reg __425078_425078;
   reg _425079_425079 ; 
   reg __425079_425079;
   reg _425080_425080 ; 
   reg __425080_425080;
   reg _425081_425081 ; 
   reg __425081_425081;
   reg _425082_425082 ; 
   reg __425082_425082;
   reg _425083_425083 ; 
   reg __425083_425083;
   reg _425084_425084 ; 
   reg __425084_425084;
   reg _425085_425085 ; 
   reg __425085_425085;
   reg _425086_425086 ; 
   reg __425086_425086;
   reg _425087_425087 ; 
   reg __425087_425087;
   reg _425088_425088 ; 
   reg __425088_425088;
   reg _425089_425089 ; 
   reg __425089_425089;
   reg _425090_425090 ; 
   reg __425090_425090;
   reg _425091_425091 ; 
   reg __425091_425091;
   reg _425092_425092 ; 
   reg __425092_425092;
   reg _425093_425093 ; 
   reg __425093_425093;
   reg _425094_425094 ; 
   reg __425094_425094;
   reg _425095_425095 ; 
   reg __425095_425095;
   reg _425096_425096 ; 
   reg __425096_425096;
   reg _425097_425097 ; 
   reg __425097_425097;
   reg _425098_425098 ; 
   reg __425098_425098;
   reg _425099_425099 ; 
   reg __425099_425099;
   reg _425100_425100 ; 
   reg __425100_425100;
   reg _425101_425101 ; 
   reg __425101_425101;
   reg _425102_425102 ; 
   reg __425102_425102;
   reg _425103_425103 ; 
   reg __425103_425103;
   reg _425104_425104 ; 
   reg __425104_425104;
   reg _425105_425105 ; 
   reg __425105_425105;
   reg _425106_425106 ; 
   reg __425106_425106;
   reg _425107_425107 ; 
   reg __425107_425107;
   reg _425108_425108 ; 
   reg __425108_425108;
   reg _425109_425109 ; 
   reg __425109_425109;
   reg _425110_425110 ; 
   reg __425110_425110;
   reg _425111_425111 ; 
   reg __425111_425111;
   reg _425112_425112 ; 
   reg __425112_425112;
   reg _425113_425113 ; 
   reg __425113_425113;
   reg _425114_425114 ; 
   reg __425114_425114;
   reg _425115_425115 ; 
   reg __425115_425115;
   reg _425116_425116 ; 
   reg __425116_425116;
   reg _425117_425117 ; 
   reg __425117_425117;
   reg _425118_425118 ; 
   reg __425118_425118;
   reg _425119_425119 ; 
   reg __425119_425119;
   reg _425120_425120 ; 
   reg __425120_425120;
   reg _425121_425121 ; 
   reg __425121_425121;
   reg _425122_425122 ; 
   reg __425122_425122;
   reg _425123_425123 ; 
   reg __425123_425123;
   reg _425124_425124 ; 
   reg __425124_425124;
   reg _425125_425125 ; 
   reg __425125_425125;
   reg _425126_425126 ; 
   reg __425126_425126;
   reg _425127_425127 ; 
   reg __425127_425127;
   reg _425128_425128 ; 
   reg __425128_425128;
   reg _425129_425129 ; 
   reg __425129_425129;
   reg _425130_425130 ; 
   reg __425130_425130;
   reg _425131_425131 ; 
   reg __425131_425131;
   reg _425132_425132 ; 
   reg __425132_425132;
   reg _425133_425133 ; 
   reg __425133_425133;
   reg _425134_425134 ; 
   reg __425134_425134;
   reg _425135_425135 ; 
   reg __425135_425135;
   reg _425136_425136 ; 
   reg __425136_425136;
   reg _425137_425137 ; 
   reg __425137_425137;
   reg _425138_425138 ; 
   reg __425138_425138;
   reg _425139_425139 ; 
   reg __425139_425139;
   reg _425140_425140 ; 
   reg __425140_425140;
   reg _425141_425141 ; 
   reg __425141_425141;
   reg _425142_425142 ; 
   reg __425142_425142;
   reg _425143_425143 ; 
   reg __425143_425143;
   reg _425144_425144 ; 
   reg __425144_425144;
   reg _425145_425145 ; 
   reg __425145_425145;
   reg _425146_425146 ; 
   reg __425146_425146;
   reg _425147_425147 ; 
   reg __425147_425147;
   reg _425148_425148 ; 
   reg __425148_425148;
   reg _425149_425149 ; 
   reg __425149_425149;
   reg _425150_425150 ; 
   reg __425150_425150;
   reg _425151_425151 ; 
   reg __425151_425151;
   reg _425152_425152 ; 
   reg __425152_425152;
   reg _425153_425153 ; 
   reg __425153_425153;
   reg _425154_425154 ; 
   reg __425154_425154;
   reg _425155_425155 ; 
   reg __425155_425155;
   reg _425156_425156 ; 
   reg __425156_425156;
   reg _425157_425157 ; 
   reg __425157_425157;
   reg _425158_425158 ; 
   reg __425158_425158;
   reg _425159_425159 ; 
   reg __425159_425159;
   reg _425160_425160 ; 
   reg __425160_425160;
   reg _425161_425161 ; 
   reg __425161_425161;
   reg _425162_425162 ; 
   reg __425162_425162;
   reg _425163_425163 ; 
   reg __425163_425163;
   reg _425164_425164 ; 
   reg __425164_425164;
   reg _425165_425165 ; 
   reg __425165_425165;
   reg _425166_425166 ; 
   reg __425166_425166;
   reg _425167_425167 ; 
   reg __425167_425167;
   reg _425168_425168 ; 
   reg __425168_425168;
   reg _425169_425169 ; 
   reg __425169_425169;
   reg _425170_425170 ; 
   reg __425170_425170;
   reg _425171_425171 ; 
   reg __425171_425171;
   reg _425172_425172 ; 
   reg __425172_425172;
   reg _425173_425173 ; 
   reg __425173_425173;
   reg _425174_425174 ; 
   reg __425174_425174;
   reg _425175_425175 ; 
   reg __425175_425175;
   reg _425176_425176 ; 
   reg __425176_425176;
   reg _425177_425177 ; 
   reg __425177_425177;
   reg _425178_425178 ; 
   reg __425178_425178;
   reg _425179_425179 ; 
   reg __425179_425179;
   reg _425180_425180 ; 
   reg __425180_425180;
   reg _425181_425181 ; 
   reg __425181_425181;
   reg _425182_425182 ; 
   reg __425182_425182;
   reg _425183_425183 ; 
   reg __425183_425183;
   reg _425184_425184 ; 
   reg __425184_425184;
   reg _425185_425185 ; 
   reg __425185_425185;
   reg _425186_425186 ; 
   reg __425186_425186;
   reg _425187_425187 ; 
   reg __425187_425187;
   reg _425188_425188 ; 
   reg __425188_425188;
   reg _425189_425189 ; 
   reg __425189_425189;
   reg _425190_425190 ; 
   reg __425190_425190;
   reg _425191_425191 ; 
   reg __425191_425191;
   reg _425192_425192 ; 
   reg __425192_425192;
   reg _425193_425193 ; 
   reg __425193_425193;
   reg _425194_425194 ; 
   reg __425194_425194;
   reg _425195_425195 ; 
   reg __425195_425195;
   reg _425196_425196 ; 
   reg __425196_425196;
   reg _425197_425197 ; 
   reg __425197_425197;
   reg _425198_425198 ; 
   reg __425198_425198;
   reg _425199_425199 ; 
   reg __425199_425199;
   reg _425200_425200 ; 
   reg __425200_425200;
   reg _425201_425201 ; 
   reg __425201_425201;
   reg _425202_425202 ; 
   reg __425202_425202;
   reg _425203_425203 ; 
   reg __425203_425203;
   reg _425204_425204 ; 
   reg __425204_425204;
   reg _425205_425205 ; 
   reg __425205_425205;
   reg _425206_425206 ; 
   reg __425206_425206;
   reg _425207_425207 ; 
   reg __425207_425207;
   reg _425208_425208 ; 
   reg __425208_425208;
   reg _425209_425209 ; 
   reg __425209_425209;
   reg _425210_425210 ; 
   reg __425210_425210;
   reg _425211_425211 ; 
   reg __425211_425211;
   reg _425212_425212 ; 
   reg __425212_425212;
   reg _425213_425213 ; 
   reg __425213_425213;
   reg _425214_425214 ; 
   reg __425214_425214;
   reg _425215_425215 ; 
   reg __425215_425215;
   reg _425216_425216 ; 
   reg __425216_425216;
   reg _425217_425217 ; 
   reg __425217_425217;
   reg _425218_425218 ; 
   reg __425218_425218;
   reg _425219_425219 ; 
   reg __425219_425219;
   reg _425220_425220 ; 
   reg __425220_425220;
   reg _425221_425221 ; 
   reg __425221_425221;
   reg _425222_425222 ; 
   reg __425222_425222;
   reg _425223_425223 ; 
   reg __425223_425223;
   reg _425224_425224 ; 
   reg __425224_425224;
   reg _425225_425225 ; 
   reg __425225_425225;
   reg _425226_425226 ; 
   reg __425226_425226;
   reg _425227_425227 ; 
   reg __425227_425227;
   reg _425228_425228 ; 
   reg __425228_425228;
   reg _425229_425229 ; 
   reg __425229_425229;
   reg _425230_425230 ; 
   reg __425230_425230;
   reg _425231_425231 ; 
   reg __425231_425231;
   reg _425232_425232 ; 
   reg __425232_425232;
   reg _425233_425233 ; 
   reg __425233_425233;
   reg _425234_425234 ; 
   reg __425234_425234;
   reg _425235_425235 ; 
   reg __425235_425235;
   reg _425236_425236 ; 
   reg __425236_425236;
   reg _425237_425237 ; 
   reg __425237_425237;
   reg _425238_425238 ; 
   reg __425238_425238;
   reg _425239_425239 ; 
   reg __425239_425239;
   reg _425240_425240 ; 
   reg __425240_425240;
   reg _425241_425241 ; 
   reg __425241_425241;
   reg _425242_425242 ; 
   reg __425242_425242;
   reg _425243_425243 ; 
   reg __425243_425243;
   reg _425244_425244 ; 
   reg __425244_425244;
   reg _425245_425245 ; 
   reg __425245_425245;
   reg _425246_425246 ; 
   reg __425246_425246;
   reg _425247_425247 ; 
   reg __425247_425247;
   reg _425248_425248 ; 
   reg __425248_425248;
   reg _425249_425249 ; 
   reg __425249_425249;
   reg _425250_425250 ; 
   reg __425250_425250;
   reg _425251_425251 ; 
   reg __425251_425251;
   reg _425252_425252 ; 
   reg __425252_425252;
   reg _425253_425253 ; 
   reg __425253_425253;
   reg _425254_425254 ; 
   reg __425254_425254;
   reg _425255_425255 ; 
   reg __425255_425255;
   reg _425256_425256 ; 
   reg __425256_425256;
   reg _425257_425257 ; 
   reg __425257_425257;
   reg _425258_425258 ; 
   reg __425258_425258;
   reg _425259_425259 ; 
   reg __425259_425259;
   reg _425260_425260 ; 
   reg __425260_425260;
   reg _425261_425261 ; 
   reg __425261_425261;
   reg _425262_425262 ; 
   reg __425262_425262;
   reg _425263_425263 ; 
   reg __425263_425263;
   reg _425264_425264 ; 
   reg __425264_425264;
   reg _425265_425265 ; 
   reg __425265_425265;
   reg _425266_425266 ; 
   reg __425266_425266;
   reg _425267_425267 ; 
   reg __425267_425267;
   reg _425268_425268 ; 
   reg __425268_425268;
   reg _425269_425269 ; 
   reg __425269_425269;
   reg _425270_425270 ; 
   reg __425270_425270;
   reg _425271_425271 ; 
   reg __425271_425271;
   reg _425272_425272 ; 
   reg __425272_425272;
   reg _425273_425273 ; 
   reg __425273_425273;
   reg _425274_425274 ; 
   reg __425274_425274;
   reg _425275_425275 ; 
   reg __425275_425275;
   reg _425276_425276 ; 
   reg __425276_425276;
   reg _425277_425277 ; 
   reg __425277_425277;
   reg _425278_425278 ; 
   reg __425278_425278;
   reg _425279_425279 ; 
   reg __425279_425279;
   reg _425280_425280 ; 
   reg __425280_425280;
   reg _425281_425281 ; 
   reg __425281_425281;
   reg _425282_425282 ; 
   reg __425282_425282;
   reg _425283_425283 ; 
   reg __425283_425283;
   reg _425284_425284 ; 
   reg __425284_425284;
   reg _425285_425285 ; 
   reg __425285_425285;
   reg _425286_425286 ; 
   reg __425286_425286;
   reg _425287_425287 ; 
   reg __425287_425287;
   reg _425288_425288 ; 
   reg __425288_425288;
   reg _425289_425289 ; 
   reg __425289_425289;
   reg _425290_425290 ; 
   reg __425290_425290;
   reg _425291_425291 ; 
   reg __425291_425291;
   reg _425292_425292 ; 
   reg __425292_425292;
   reg _425293_425293 ; 
   reg __425293_425293;
   reg _425294_425294 ; 
   reg __425294_425294;
   reg _425295_425295 ; 
   reg __425295_425295;
   reg _425296_425296 ; 
   reg __425296_425296;
   reg _425297_425297 ; 
   reg __425297_425297;
   reg _425298_425298 ; 
   reg __425298_425298;
   reg _425299_425299 ; 
   reg __425299_425299;
   reg _425300_425300 ; 
   reg __425300_425300;
   reg _425301_425301 ; 
   reg __425301_425301;
   reg _425302_425302 ; 
   reg __425302_425302;
   reg _425303_425303 ; 
   reg __425303_425303;
   reg _425304_425304 ; 
   reg __425304_425304;
   reg _425305_425305 ; 
   reg __425305_425305;
   reg _425306_425306 ; 
   reg __425306_425306;
   reg _425307_425307 ; 
   reg __425307_425307;
   reg _425308_425308 ; 
   reg __425308_425308;
   reg _425309_425309 ; 
   reg __425309_425309;
   reg _425310_425310 ; 
   reg __425310_425310;
   reg _425311_425311 ; 
   reg __425311_425311;
   reg _425312_425312 ; 
   reg __425312_425312;
   reg _425313_425313 ; 
   reg __425313_425313;
   reg _425314_425314 ; 
   reg __425314_425314;
   reg _425315_425315 ; 
   reg __425315_425315;
   reg _425316_425316 ; 
   reg __425316_425316;
   reg _425317_425317 ; 
   reg __425317_425317;
   reg _425318_425318 ; 
   reg __425318_425318;
   reg _425319_425319 ; 
   reg __425319_425319;
   reg _425320_425320 ; 
   reg __425320_425320;
   reg _425321_425321 ; 
   reg __425321_425321;
   reg _425322_425322 ; 
   reg __425322_425322;
   reg _425323_425323 ; 
   reg __425323_425323;
   reg _425324_425324 ; 
   reg __425324_425324;
   reg _425325_425325 ; 
   reg __425325_425325;
   reg _425326_425326 ; 
   reg __425326_425326;
   reg _425327_425327 ; 
   reg __425327_425327;
   reg _425328_425328 ; 
   reg __425328_425328;
   reg _425329_425329 ; 
   reg __425329_425329;
   reg _425330_425330 ; 
   reg __425330_425330;
   reg _425331_425331 ; 
   reg __425331_425331;
   reg _425332_425332 ; 
   reg __425332_425332;
   reg _425333_425333 ; 
   reg __425333_425333;
   reg _425334_425334 ; 
   reg __425334_425334;
   reg _425335_425335 ; 
   reg __425335_425335;
   reg _425336_425336 ; 
   reg __425336_425336;
   reg _425337_425337 ; 
   reg __425337_425337;
   reg _425338_425338 ; 
   reg __425338_425338;
   reg _425339_425339 ; 
   reg __425339_425339;
   reg _425340_425340 ; 
   reg __425340_425340;
   reg _425341_425341 ; 
   reg __425341_425341;
   reg _425342_425342 ; 
   reg __425342_425342;
   reg _425343_425343 ; 
   reg __425343_425343;
   reg _425344_425344 ; 
   reg __425344_425344;
   reg _425345_425345 ; 
   reg __425345_425345;
   reg _425346_425346 ; 
   reg __425346_425346;
   reg _425347_425347 ; 
   reg __425347_425347;
   reg _425348_425348 ; 
   reg __425348_425348;
   reg _425349_425349 ; 
   reg __425349_425349;
   reg _425350_425350 ; 
   reg __425350_425350;
   reg _425351_425351 ; 
   reg __425351_425351;
   reg _425352_425352 ; 
   reg __425352_425352;
   reg _425353_425353 ; 
   reg __425353_425353;
   reg _425354_425354 ; 
   reg __425354_425354;
   reg _425355_425355 ; 
   reg __425355_425355;
   reg _425356_425356 ; 
   reg __425356_425356;
   reg _425357_425357 ; 
   reg __425357_425357;
   reg _425358_425358 ; 
   reg __425358_425358;
   reg _425359_425359 ; 
   reg __425359_425359;
   reg _425360_425360 ; 
   reg __425360_425360;
   reg _425361_425361 ; 
   reg __425361_425361;
   reg _425362_425362 ; 
   reg __425362_425362;
   reg _425363_425363 ; 
   reg __425363_425363;
   reg _425364_425364 ; 
   reg __425364_425364;
   reg _425365_425365 ; 
   reg __425365_425365;
   reg _425366_425366 ; 
   reg __425366_425366;
   reg _425367_425367 ; 
   reg __425367_425367;
   reg _425368_425368 ; 
   reg __425368_425368;
   reg _425369_425369 ; 
   reg __425369_425369;
   reg _425370_425370 ; 
   reg __425370_425370;
   reg _425371_425371 ; 
   reg __425371_425371;
   reg _425372_425372 ; 
   reg __425372_425372;
   reg _425373_425373 ; 
   reg __425373_425373;
   reg _425374_425374 ; 
   reg __425374_425374;
   reg _425375_425375 ; 
   reg __425375_425375;
   reg _425376_425376 ; 
   reg __425376_425376;
   reg _425377_425377 ; 
   reg __425377_425377;
   reg _425378_425378 ; 
   reg __425378_425378;
   reg _425379_425379 ; 
   reg __425379_425379;
   reg _425380_425380 ; 
   reg __425380_425380;
   reg _425381_425381 ; 
   reg __425381_425381;
   reg _425382_425382 ; 
   reg __425382_425382;
   reg _425383_425383 ; 
   reg __425383_425383;
   reg _425384_425384 ; 
   reg __425384_425384;
   reg _425385_425385 ; 
   reg __425385_425385;
   reg _425386_425386 ; 
   reg __425386_425386;
   reg _425387_425387 ; 
   reg __425387_425387;
   reg _425388_425388 ; 
   reg __425388_425388;
   reg _425389_425389 ; 
   reg __425389_425389;
   reg _425390_425390 ; 
   reg __425390_425390;
   reg _425391_425391 ; 
   reg __425391_425391;
   reg _425392_425392 ; 
   reg __425392_425392;
   reg _425393_425393 ; 
   reg __425393_425393;
   reg _425394_425394 ; 
   reg __425394_425394;
   reg _425395_425395 ; 
   reg __425395_425395;
   reg _425396_425396 ; 
   reg __425396_425396;
   reg _425397_425397 ; 
   reg __425397_425397;
   reg _425398_425398 ; 
   reg __425398_425398;
   reg _425399_425399 ; 
   reg __425399_425399;
   reg _425400_425400 ; 
   reg __425400_425400;
   reg _425401_425401 ; 
   reg __425401_425401;
   reg _425402_425402 ; 
   reg __425402_425402;
   reg _425403_425403 ; 
   reg __425403_425403;
   reg _425404_425404 ; 
   reg __425404_425404;
   reg _425405_425405 ; 
   reg __425405_425405;
   reg _425406_425406 ; 
   reg __425406_425406;
   reg _425407_425407 ; 
   reg __425407_425407;
   reg _425408_425408 ; 
   reg __425408_425408;
   reg _425409_425409 ; 
   reg __425409_425409;
   reg _425410_425410 ; 
   reg __425410_425410;
   reg _425411_425411 ; 
   reg __425411_425411;
   reg _425412_425412 ; 
   reg __425412_425412;
   reg _425413_425413 ; 
   reg __425413_425413;
   reg _425414_425414 ; 
   reg __425414_425414;
   reg _425415_425415 ; 
   reg __425415_425415;
   reg _425416_425416 ; 
   reg __425416_425416;
   reg _425417_425417 ; 
   reg __425417_425417;
   reg _425418_425418 ; 
   reg __425418_425418;
   reg _425419_425419 ; 
   reg __425419_425419;
   reg _425420_425420 ; 
   reg __425420_425420;
   reg _425421_425421 ; 
   reg __425421_425421;
   reg _425422_425422 ; 
   reg __425422_425422;
   reg _425423_425423 ; 
   reg __425423_425423;
   reg _425424_425424 ; 
   reg __425424_425424;
   reg _425425_425425 ; 
   reg __425425_425425;
   reg _425426_425426 ; 
   reg __425426_425426;
   reg _425427_425427 ; 
   reg __425427_425427;
   reg _425428_425428 ; 
   reg __425428_425428;
   reg _425429_425429 ; 
   reg __425429_425429;
   reg _425430_425430 ; 
   reg __425430_425430;
   reg _425431_425431 ; 
   reg __425431_425431;
   reg _425432_425432 ; 
   reg __425432_425432;
   reg _425433_425433 ; 
   reg __425433_425433;
   reg _425434_425434 ; 
   reg __425434_425434;
   reg _425435_425435 ; 
   reg __425435_425435;
   reg _425436_425436 ; 
   reg __425436_425436;
   reg _425437_425437 ; 
   reg __425437_425437;
   reg _425438_425438 ; 
   reg __425438_425438;
   reg _425439_425439 ; 
   reg __425439_425439;
   reg _425440_425440 ; 
   reg __425440_425440;
   reg _425441_425441 ; 
   reg __425441_425441;
   reg _425442_425442 ; 
   reg __425442_425442;
   reg _425443_425443 ; 
   reg __425443_425443;
   reg _425444_425444 ; 
   reg __425444_425444;
   reg _425445_425445 ; 
   reg __425445_425445;
   reg _425446_425446 ; 
   reg __425446_425446;
   reg _425447_425447 ; 
   reg __425447_425447;
   reg _425448_425448 ; 
   reg __425448_425448;
   reg _425449_425449 ; 
   reg __425449_425449;
   reg _425450_425450 ; 
   reg __425450_425450;
   reg _425451_425451 ; 
   reg __425451_425451;
   reg _425452_425452 ; 
   reg __425452_425452;
   reg _425453_425453 ; 
   reg __425453_425453;
   reg _425454_425454 ; 
   reg __425454_425454;
   reg _425455_425455 ; 
   reg __425455_425455;
   reg _425456_425456 ; 
   reg __425456_425456;
   reg _425457_425457 ; 
   reg __425457_425457;
   reg _425458_425458 ; 
   reg __425458_425458;
   reg _425459_425459 ; 
   reg __425459_425459;
   reg _425460_425460 ; 
   reg __425460_425460;
   reg _425461_425461 ; 
   reg __425461_425461;
   reg _425462_425462 ; 
   reg __425462_425462;
   reg _425463_425463 ; 
   reg __425463_425463;
   reg _425464_425464 ; 
   reg __425464_425464;
   reg _425465_425465 ; 
   reg __425465_425465;
   reg _425466_425466 ; 
   reg __425466_425466;
   reg _425467_425467 ; 
   reg __425467_425467;
   reg _425468_425468 ; 
   reg __425468_425468;
   reg _425469_425469 ; 
   reg __425469_425469;
   reg _425470_425470 ; 
   reg __425470_425470;
   reg _425471_425471 ; 
   reg __425471_425471;
   reg _425472_425472 ; 
   reg __425472_425472;
   reg _425473_425473 ; 
   reg __425473_425473;
   reg _425474_425474 ; 
   reg __425474_425474;
   reg _425475_425475 ; 
   reg __425475_425475;
   reg _425476_425476 ; 
   reg __425476_425476;
   reg _425477_425477 ; 
   reg __425477_425477;
   reg _425478_425478 ; 
   reg __425478_425478;
   reg _425479_425479 ; 
   reg __425479_425479;
   reg _425480_425480 ; 
   reg __425480_425480;
   reg _425481_425481 ; 
   reg __425481_425481;
   reg _425482_425482 ; 
   reg __425482_425482;
   reg _425483_425483 ; 
   reg __425483_425483;
   reg _425484_425484 ; 
   reg __425484_425484;
   reg _425485_425485 ; 
   reg __425485_425485;
   reg _425486_425486 ; 
   reg __425486_425486;
   reg _425487_425487 ; 
   reg __425487_425487;
   reg _425488_425488 ; 
   reg __425488_425488;
   reg _425489_425489 ; 
   reg __425489_425489;
   reg _425490_425490 ; 
   reg __425490_425490;
   reg _425491_425491 ; 
   reg __425491_425491;
   reg _425492_425492 ; 
   reg __425492_425492;
   reg _425493_425493 ; 
   reg __425493_425493;
   reg _425494_425494 ; 
   reg __425494_425494;
   reg _425495_425495 ; 
   reg __425495_425495;
   reg _425496_425496 ; 
   reg __425496_425496;
   reg _425497_425497 ; 
   reg __425497_425497;
   reg _425498_425498 ; 
   reg __425498_425498;
   reg _425499_425499 ; 
   reg __425499_425499;
   reg _425500_425500 ; 
   reg __425500_425500;
   reg _425501_425501 ; 
   reg __425501_425501;
   reg _425502_425502 ; 
   reg __425502_425502;
   reg _425503_425503 ; 
   reg __425503_425503;
   reg _425504_425504 ; 
   reg __425504_425504;
   reg _425505_425505 ; 
   reg __425505_425505;
   reg _425506_425506 ; 
   reg __425506_425506;
   reg _425507_425507 ; 
   reg __425507_425507;
   reg _425508_425508 ; 
   reg __425508_425508;
   reg _425509_425509 ; 
   reg __425509_425509;
   reg _425510_425510 ; 
   reg __425510_425510;
   reg _425511_425511 ; 
   reg __425511_425511;
   reg _425512_425512 ; 
   reg __425512_425512;
   reg _425513_425513 ; 
   reg __425513_425513;
   reg _425514_425514 ; 
   reg __425514_425514;
   reg _425515_425515 ; 
   reg __425515_425515;
   reg _425516_425516 ; 
   reg __425516_425516;
   reg _425517_425517 ; 
   reg __425517_425517;
   reg _425518_425518 ; 
   reg __425518_425518;
   reg _425519_425519 ; 
   reg __425519_425519;
   reg _425520_425520 ; 
   reg __425520_425520;
   reg _425521_425521 ; 
   reg __425521_425521;
   reg _425522_425522 ; 
   reg __425522_425522;
   reg _425523_425523 ; 
   reg __425523_425523;
   reg _425524_425524 ; 
   reg __425524_425524;
   reg _425525_425525 ; 
   reg __425525_425525;
   reg _425526_425526 ; 
   reg __425526_425526;
   reg _425527_425527 ; 
   reg __425527_425527;
   reg _425528_425528 ; 
   reg __425528_425528;
   reg _425529_425529 ; 
   reg __425529_425529;
   reg _425530_425530 ; 
   reg __425530_425530;
   reg _425531_425531 ; 
   reg __425531_425531;
   reg _425532_425532 ; 
   reg __425532_425532;
   reg _425533_425533 ; 
   reg __425533_425533;
   reg _425534_425534 ; 
   reg __425534_425534;
   reg _425535_425535 ; 
   reg __425535_425535;
   reg _425536_425536 ; 
   reg __425536_425536;
   reg _425537_425537 ; 
   reg __425537_425537;
   reg _425538_425538 ; 
   reg __425538_425538;
   reg _425539_425539 ; 
   reg __425539_425539;
   reg _425540_425540 ; 
   reg __425540_425540;
   reg _425541_425541 ; 
   reg __425541_425541;
   reg _425542_425542 ; 
   reg __425542_425542;
   reg _425543_425543 ; 
   reg __425543_425543;
   reg _425544_425544 ; 
   reg __425544_425544;
   reg _425545_425545 ; 
   reg __425545_425545;
   reg _425546_425546 ; 
   reg __425546_425546;
   reg _425547_425547 ; 
   reg __425547_425547;
   reg _425548_425548 ; 
   reg __425548_425548;
   reg _425549_425549 ; 
   reg __425549_425549;
   reg _425550_425550 ; 
   reg __425550_425550;
   reg _425551_425551 ; 
   reg __425551_425551;
   reg _425552_425552 ; 
   reg __425552_425552;
   reg _425553_425553 ; 
   reg __425553_425553;
   reg _425554_425554 ; 
   reg __425554_425554;
   reg _425555_425555 ; 
   reg __425555_425555;
   reg _425556_425556 ; 
   reg __425556_425556;
   reg _425557_425557 ; 
   reg __425557_425557;
   reg _425558_425558 ; 
   reg __425558_425558;
   reg _425559_425559 ; 
   reg __425559_425559;
   reg _425560_425560 ; 
   reg __425560_425560;
   reg _425561_425561 ; 
   reg __425561_425561;
   reg _425562_425562 ; 
   reg __425562_425562;
   reg _425563_425563 ; 
   reg __425563_425563;
   reg _425564_425564 ; 
   reg __425564_425564;
   reg _425565_425565 ; 
   reg __425565_425565;
   reg _425566_425566 ; 
   reg __425566_425566;
   reg _425567_425567 ; 
   reg __425567_425567;
   reg _425568_425568 ; 
   reg __425568_425568;
   reg _425569_425569 ; 
   reg __425569_425569;
   reg _425570_425570 ; 
   reg __425570_425570;
   reg _425571_425571 ; 
   reg __425571_425571;
   reg _425572_425572 ; 
   reg __425572_425572;
   reg _425573_425573 ; 
   reg __425573_425573;
   reg _425574_425574 ; 
   reg __425574_425574;
   reg _425575_425575 ; 
   reg __425575_425575;
   reg _425576_425576 ; 
   reg __425576_425576;
   reg _425577_425577 ; 
   reg __425577_425577;
   reg _425578_425578 ; 
   reg __425578_425578;
   reg _425579_425579 ; 
   reg __425579_425579;
   reg _425580_425580 ; 
   reg __425580_425580;
   reg _425581_425581 ; 
   reg __425581_425581;
   reg _425582_425582 ; 
   reg __425582_425582;
   reg _425583_425583 ; 
   reg __425583_425583;
   reg _425584_425584 ; 
   reg __425584_425584;
   reg _425585_425585 ; 
   reg __425585_425585;
   reg _425586_425586 ; 
   reg __425586_425586;
   reg _425587_425587 ; 
   reg __425587_425587;
   reg _425588_425588 ; 
   reg __425588_425588;
   reg _425589_425589 ; 
   reg __425589_425589;
   reg _425590_425590 ; 
   reg __425590_425590;
   reg _425591_425591 ; 
   reg __425591_425591;
   reg _425592_425592 ; 
   reg __425592_425592;
   reg _425593_425593 ; 
   reg __425593_425593;
   reg _425594_425594 ; 
   reg __425594_425594;
   reg _425595_425595 ; 
   reg __425595_425595;
   reg _425596_425596 ; 
   reg __425596_425596;
   reg _425597_425597 ; 
   reg __425597_425597;
   reg _425598_425598 ; 
   reg __425598_425598;
   reg _425599_425599 ; 
   reg __425599_425599;
   reg _425600_425600 ; 
   reg __425600_425600;
   reg _425601_425601 ; 
   reg __425601_425601;
   reg _425602_425602 ; 
   reg __425602_425602;
   reg _425603_425603 ; 
   reg __425603_425603;
   reg _425604_425604 ; 
   reg __425604_425604;
   reg _425605_425605 ; 
   reg __425605_425605;
   reg _425606_425606 ; 
   reg __425606_425606;
   reg _425607_425607 ; 
   reg __425607_425607;
   reg _425608_425608 ; 
   reg __425608_425608;
   reg _425609_425609 ; 
   reg __425609_425609;
   reg _425610_425610 ; 
   reg __425610_425610;
   reg _425611_425611 ; 
   reg __425611_425611;
   reg _425612_425612 ; 
   reg __425612_425612;
   reg _425613_425613 ; 
   reg __425613_425613;
   reg _425614_425614 ; 
   reg __425614_425614;
   reg _425615_425615 ; 
   reg __425615_425615;
   reg _425616_425616 ; 
   reg __425616_425616;
   reg _425617_425617 ; 
   reg __425617_425617;
   reg _425618_425618 ; 
   reg __425618_425618;
   reg _425619_425619 ; 
   reg __425619_425619;
   reg _425620_425620 ; 
   reg __425620_425620;
   reg _425621_425621 ; 
   reg __425621_425621;
   reg _425622_425622 ; 
   reg __425622_425622;
   reg _425623_425623 ; 
   reg __425623_425623;
   reg _425624_425624 ; 
   reg __425624_425624;
   reg _425625_425625 ; 
   reg __425625_425625;
   reg _425626_425626 ; 
   reg __425626_425626;
   reg _425627_425627 ; 
   reg __425627_425627;
   reg _425628_425628 ; 
   reg __425628_425628;
   reg _425629_425629 ; 
   reg __425629_425629;
   reg _425630_425630 ; 
   reg __425630_425630;
   reg _425631_425631 ; 
   reg __425631_425631;
   reg _425632_425632 ; 
   reg __425632_425632;
   reg _425633_425633 ; 
   reg __425633_425633;
   reg _425634_425634 ; 
   reg __425634_425634;
   reg _425635_425635 ; 
   reg __425635_425635;
   reg _425636_425636 ; 
   reg __425636_425636;
   reg _425637_425637 ; 
   reg __425637_425637;
   reg _425638_425638 ; 
   reg __425638_425638;
   reg _425639_425639 ; 
   reg __425639_425639;
   reg _425640_425640 ; 
   reg __425640_425640;
   reg _425641_425641 ; 
   reg __425641_425641;
   reg _425642_425642 ; 
   reg __425642_425642;
   reg _425643_425643 ; 
   reg __425643_425643;
   reg _425644_425644 ; 
   reg __425644_425644;
   reg _425645_425645 ; 
   reg __425645_425645;
   reg _425646_425646 ; 
   reg __425646_425646;
   reg _425647_425647 ; 
   reg __425647_425647;
   reg _425648_425648 ; 
   reg __425648_425648;
   reg _425649_425649 ; 
   reg __425649_425649;
   reg _425650_425650 ; 
   reg __425650_425650;
   reg _425651_425651 ; 
   reg __425651_425651;
   reg _425652_425652 ; 
   reg __425652_425652;
   reg _425653_425653 ; 
   reg __425653_425653;
   reg _425654_425654 ; 
   reg __425654_425654;
   reg _425655_425655 ; 
   reg __425655_425655;
   reg _425656_425656 ; 
   reg __425656_425656;
   reg _425657_425657 ; 
   reg __425657_425657;
   reg _425658_425658 ; 
   reg __425658_425658;
   reg _425659_425659 ; 
   reg __425659_425659;
   reg _425660_425660 ; 
   reg __425660_425660;
   reg _425661_425661 ; 
   reg __425661_425661;
   reg _425662_425662 ; 
   reg __425662_425662;
   reg _425663_425663 ; 
   reg __425663_425663;
   reg _425664_425664 ; 
   reg __425664_425664;
   reg _425665_425665 ; 
   reg __425665_425665;
   reg _425666_425666 ; 
   reg __425666_425666;
   reg _425667_425667 ; 
   reg __425667_425667;
   reg _425668_425668 ; 
   reg __425668_425668;
   reg _425669_425669 ; 
   reg __425669_425669;
   reg _425670_425670 ; 
   reg __425670_425670;
   reg _425671_425671 ; 
   reg __425671_425671;
   reg _425672_425672 ; 
   reg __425672_425672;
   reg _425673_425673 ; 
   reg __425673_425673;
   reg _425674_425674 ; 
   reg __425674_425674;
   reg _425675_425675 ; 
   reg __425675_425675;
   reg _425676_425676 ; 
   reg __425676_425676;
   reg _425677_425677 ; 
   reg __425677_425677;
   reg _425678_425678 ; 
   reg __425678_425678;
   reg _425679_425679 ; 
   reg __425679_425679;
   reg _425680_425680 ; 
   reg __425680_425680;
   reg _425681_425681 ; 
   reg __425681_425681;
   reg _425682_425682 ; 
   reg __425682_425682;
   reg _425683_425683 ; 
   reg __425683_425683;
   reg _425684_425684 ; 
   reg __425684_425684;
   reg _425685_425685 ; 
   reg __425685_425685;
   reg _425686_425686 ; 
   reg __425686_425686;
   reg _425687_425687 ; 
   reg __425687_425687;
   reg _425688_425688 ; 
   reg __425688_425688;
   reg _425689_425689 ; 
   reg __425689_425689;
   reg _425690_425690 ; 
   reg __425690_425690;
   reg _425691_425691 ; 
   reg __425691_425691;
   reg _425692_425692 ; 
   reg __425692_425692;
   reg _425693_425693 ; 
   reg __425693_425693;
   reg _425694_425694 ; 
   reg __425694_425694;
   reg _425695_425695 ; 
   reg __425695_425695;
   reg _425696_425696 ; 
   reg __425696_425696;
   reg _425697_425697 ; 
   reg __425697_425697;
   reg _425698_425698 ; 
   reg __425698_425698;
   reg _425699_425699 ; 
   reg __425699_425699;
   reg _425700_425700 ; 
   reg __425700_425700;
   reg _425701_425701 ; 
   reg __425701_425701;
   reg _425702_425702 ; 
   reg __425702_425702;
   reg _425703_425703 ; 
   reg __425703_425703;
   reg _425704_425704 ; 
   reg __425704_425704;
   reg _425705_425705 ; 
   reg __425705_425705;
   reg _425706_425706 ; 
   reg __425706_425706;
   reg _425707_425707 ; 
   reg __425707_425707;
   reg _425708_425708 ; 
   reg __425708_425708;
   reg _425709_425709 ; 
   reg __425709_425709;
   reg _425710_425710 ; 
   reg __425710_425710;
   reg _425711_425711 ; 
   reg __425711_425711;
   reg _425712_425712 ; 
   reg __425712_425712;
   reg _425713_425713 ; 
   reg __425713_425713;
   reg _425714_425714 ; 
   reg __425714_425714;
   reg _425715_425715 ; 
   reg __425715_425715;
   reg _425716_425716 ; 
   reg __425716_425716;
   reg _425717_425717 ; 
   reg __425717_425717;
   reg _425718_425718 ; 
   reg __425718_425718;
   reg _425719_425719 ; 
   reg __425719_425719;
   reg _425720_425720 ; 
   reg __425720_425720;
   reg _425721_425721 ; 
   reg __425721_425721;
   reg _425722_425722 ; 
   reg __425722_425722;
   reg _425723_425723 ; 
   reg __425723_425723;
   reg _425724_425724 ; 
   reg __425724_425724;
   reg _425725_425725 ; 
   reg __425725_425725;
   reg _425726_425726 ; 
   reg __425726_425726;
   reg _425727_425727 ; 
   reg __425727_425727;
   reg _425728_425728 ; 
   reg __425728_425728;
   reg _425729_425729 ; 
   reg __425729_425729;
   reg _425730_425730 ; 
   reg __425730_425730;
   reg _425731_425731 ; 
   reg __425731_425731;
   reg _425732_425732 ; 
   reg __425732_425732;
   reg _425733_425733 ; 
   reg __425733_425733;
   reg _425734_425734 ; 
   reg __425734_425734;
   reg _425735_425735 ; 
   reg __425735_425735;
   reg _425736_425736 ; 
   reg __425736_425736;
   reg _425737_425737 ; 
   reg __425737_425737;
   reg _425738_425738 ; 
   reg __425738_425738;
   reg _425739_425739 ; 
   reg __425739_425739;
   reg _425740_425740 ; 
   reg __425740_425740;
   reg _425741_425741 ; 
   reg __425741_425741;
   reg _425742_425742 ; 
   reg __425742_425742;
   reg _425743_425743 ; 
   reg __425743_425743;
   reg _425744_425744 ; 
   reg __425744_425744;
   reg _425745_425745 ; 
   reg __425745_425745;
   reg _425746_425746 ; 
   reg __425746_425746;
   reg _425747_425747 ; 
   reg __425747_425747;
   reg _425748_425748 ; 
   reg __425748_425748;
   reg _425749_425749 ; 
   reg __425749_425749;
   reg _425750_425750 ; 
   reg __425750_425750;
   reg _425751_425751 ; 
   reg __425751_425751;
   reg _425752_425752 ; 
   reg __425752_425752;
   reg _425753_425753 ; 
   reg __425753_425753;
   reg _425754_425754 ; 
   reg __425754_425754;
   reg _425755_425755 ; 
   reg __425755_425755;
   reg _425756_425756 ; 
   reg __425756_425756;
   reg _425757_425757 ; 
   reg __425757_425757;
   reg _425758_425758 ; 
   reg __425758_425758;
   reg _425759_425759 ; 
   reg __425759_425759;
   reg _425760_425760 ; 
   reg __425760_425760;
   reg _425761_425761 ; 
   reg __425761_425761;
   reg _425762_425762 ; 
   reg __425762_425762;
   reg _425763_425763 ; 
   reg __425763_425763;
   reg _425764_425764 ; 
   reg __425764_425764;
   reg _425765_425765 ; 
   reg __425765_425765;
   reg _425766_425766 ; 
   reg __425766_425766;
   reg _425767_425767 ; 
   reg __425767_425767;
   reg _425768_425768 ; 
   reg __425768_425768;
   reg _425769_425769 ; 
   reg __425769_425769;
   reg _425770_425770 ; 
   reg __425770_425770;
   reg _425771_425771 ; 
   reg __425771_425771;
   reg _425772_425772 ; 
   reg __425772_425772;
   reg _425773_425773 ; 
   reg __425773_425773;
   reg _425774_425774 ; 
   reg __425774_425774;
   reg _425775_425775 ; 
   reg __425775_425775;
   reg _425776_425776 ; 
   reg __425776_425776;
   reg _425777_425777 ; 
   reg __425777_425777;
   reg _425778_425778 ; 
   reg __425778_425778;
   reg _425779_425779 ; 
   reg __425779_425779;
   reg _425780_425780 ; 
   reg __425780_425780;
   reg _425781_425781 ; 
   reg __425781_425781;
   reg _425782_425782 ; 
   reg __425782_425782;
   reg _425783_425783 ; 
   reg __425783_425783;
   reg _425784_425784 ; 
   reg __425784_425784;
   reg _425785_425785 ; 
   reg __425785_425785;
   reg _425786_425786 ; 
   reg __425786_425786;
   reg _425787_425787 ; 
   reg __425787_425787;
   reg _425788_425788 ; 
   reg __425788_425788;
   reg _425789_425789 ; 
   reg __425789_425789;
   reg _425790_425790 ; 
   reg __425790_425790;
   reg _425791_425791 ; 
   reg __425791_425791;
   reg _425792_425792 ; 
   reg __425792_425792;
   reg _425793_425793 ; 
   reg __425793_425793;
   reg _425794_425794 ; 
   reg __425794_425794;
   reg _425795_425795 ; 
   reg __425795_425795;
   reg _425796_425796 ; 
   reg __425796_425796;
   reg _425797_425797 ; 
   reg __425797_425797;
   reg _425798_425798 ; 
   reg __425798_425798;
   reg _425799_425799 ; 
   reg __425799_425799;
   reg _425800_425800 ; 
   reg __425800_425800;
   reg _425801_425801 ; 
   reg __425801_425801;
   reg _425802_425802 ; 
   reg __425802_425802;
   reg _425803_425803 ; 
   reg __425803_425803;
   reg _425804_425804 ; 
   reg __425804_425804;
   reg _425805_425805 ; 
   reg __425805_425805;
   reg _425806_425806 ; 
   reg __425806_425806;
   reg _425807_425807 ; 
   reg __425807_425807;
   reg _425808_425808 ; 
   reg __425808_425808;
   reg _425809_425809 ; 
   reg __425809_425809;
   reg _425810_425810 ; 
   reg __425810_425810;
   reg _425811_425811 ; 
   reg __425811_425811;
   reg _425812_425812 ; 
   reg __425812_425812;
   reg _425813_425813 ; 
   reg __425813_425813;
   reg _425814_425814 ; 
   reg __425814_425814;
   reg _425815_425815 ; 
   reg __425815_425815;
   reg _425816_425816 ; 
   reg __425816_425816;
   reg _425817_425817 ; 
   reg __425817_425817;
   reg _425818_425818 ; 
   reg __425818_425818;
   reg _425819_425819 ; 
   reg __425819_425819;
   reg _425820_425820 ; 
   reg __425820_425820;
   reg _425821_425821 ; 
   reg __425821_425821;
   reg _425822_425822 ; 
   reg __425822_425822;
   reg _425823_425823 ; 
   reg __425823_425823;
   reg _425824_425824 ; 
   reg __425824_425824;
   reg _425825_425825 ; 
   reg __425825_425825;
   reg _425826_425826 ; 
   reg __425826_425826;
   reg _425827_425827 ; 
   reg __425827_425827;
   reg _425828_425828 ; 
   reg __425828_425828;
   reg _425829_425829 ; 
   reg __425829_425829;
   reg _425830_425830 ; 
   reg __425830_425830;
   reg _425831_425831 ; 
   reg __425831_425831;
   reg _425832_425832 ; 
   reg __425832_425832;
   reg _425833_425833 ; 
   reg __425833_425833;
   reg _425834_425834 ; 
   reg __425834_425834;
   reg _425835_425835 ; 
   reg __425835_425835;
   reg _425836_425836 ; 
   reg __425836_425836;
   reg _425837_425837 ; 
   reg __425837_425837;
   reg _425838_425838 ; 
   reg __425838_425838;
   reg _425839_425839 ; 
   reg __425839_425839;
   reg _425840_425840 ; 
   reg __425840_425840;
   reg _425841_425841 ; 
   reg __425841_425841;
   reg _425842_425842 ; 
   reg __425842_425842;
   reg _425843_425843 ; 
   reg __425843_425843;
   reg _425844_425844 ; 
   reg __425844_425844;
   reg _425845_425845 ; 
   reg __425845_425845;
   reg _425846_425846 ; 
   reg __425846_425846;
   reg _425847_425847 ; 
   reg __425847_425847;
   reg _425848_425848 ; 
   reg __425848_425848;
   reg _425849_425849 ; 
   reg __425849_425849;
   reg _425850_425850 ; 
   reg __425850_425850;
   reg _425851_425851 ; 
   reg __425851_425851;
   reg _425852_425852 ; 
   reg __425852_425852;
   reg _425853_425853 ; 
   reg __425853_425853;
   reg _425854_425854 ; 
   reg __425854_425854;
   reg _425855_425855 ; 
   reg __425855_425855;
   reg _425856_425856 ; 
   reg __425856_425856;
   reg _425857_425857 ; 
   reg __425857_425857;
   reg _425858_425858 ; 
   reg __425858_425858;
   reg _425859_425859 ; 
   reg __425859_425859;
   reg _425860_425860 ; 
   reg __425860_425860;
   reg _425861_425861 ; 
   reg __425861_425861;
   reg _425862_425862 ; 
   reg __425862_425862;
   reg _425863_425863 ; 
   reg __425863_425863;
   reg _425864_425864 ; 
   reg __425864_425864;
   reg _425865_425865 ; 
   reg __425865_425865;
   reg _425866_425866 ; 
   reg __425866_425866;
   reg _425867_425867 ; 
   reg __425867_425867;
   reg _425868_425868 ; 
   reg __425868_425868;
   reg _425869_425869 ; 
   reg __425869_425869;
   reg _425870_425870 ; 
   reg __425870_425870;
   reg _425871_425871 ; 
   reg __425871_425871;
   reg _425872_425872 ; 
   reg __425872_425872;
   reg _425873_425873 ; 
   reg __425873_425873;
   reg _425874_425874 ; 
   reg __425874_425874;
   reg _425875_425875 ; 
   reg __425875_425875;
   reg _425876_425876 ; 
   reg __425876_425876;
   reg _425877_425877 ; 
   reg __425877_425877;
   reg _425878_425878 ; 
   reg __425878_425878;
   reg _425879_425879 ; 
   reg __425879_425879;
   reg _425880_425880 ; 
   reg __425880_425880;
   reg _425881_425881 ; 
   reg __425881_425881;
   reg _425882_425882 ; 
   reg __425882_425882;
   reg _425883_425883 ; 
   reg __425883_425883;
   reg _425884_425884 ; 
   reg __425884_425884;
   reg _425885_425885 ; 
   reg __425885_425885;
   reg _425886_425886 ; 
   reg __425886_425886;
   reg _425887_425887 ; 
   reg __425887_425887;
   reg _425888_425888 ; 
   reg __425888_425888;
   reg _425889_425889 ; 
   reg __425889_425889;
   reg _425890_425890 ; 
   reg __425890_425890;
   reg _425891_425891 ; 
   reg __425891_425891;
   reg _425892_425892 ; 
   reg __425892_425892;
   reg _425893_425893 ; 
   reg __425893_425893;
   reg _425894_425894 ; 
   reg __425894_425894;
   reg _425895_425895 ; 
   reg __425895_425895;
   reg _425896_425896 ; 
   reg __425896_425896;
   reg _425897_425897 ; 
   reg __425897_425897;
   reg _425898_425898 ; 
   reg __425898_425898;
   reg _425899_425899 ; 
   reg __425899_425899;
   reg _425900_425900 ; 
   reg __425900_425900;
   reg _425901_425901 ; 
   reg __425901_425901;
   reg _425902_425902 ; 
   reg __425902_425902;
   reg _425903_425903 ; 
   reg __425903_425903;
   reg _425904_425904 ; 
   reg __425904_425904;
   reg _425905_425905 ; 
   reg __425905_425905;
   reg _425906_425906 ; 
   reg __425906_425906;
   reg _425907_425907 ; 
   reg __425907_425907;
   reg _425908_425908 ; 
   reg __425908_425908;
   reg _425909_425909 ; 
   reg __425909_425909;
   reg _425910_425910 ; 
   reg __425910_425910;
   reg _425911_425911 ; 
   reg __425911_425911;
   reg _425912_425912 ; 
   reg __425912_425912;
   reg _425913_425913 ; 
   reg __425913_425913;
   reg _425914_425914 ; 
   reg __425914_425914;
   reg _425915_425915 ; 
   reg __425915_425915;
   reg _425916_425916 ; 
   reg __425916_425916;
   reg _425917_425917 ; 
   reg __425917_425917;
   reg _425918_425918 ; 
   reg __425918_425918;
   reg _425919_425919 ; 
   reg __425919_425919;
   reg _425920_425920 ; 
   reg __425920_425920;
   reg _425921_425921 ; 
   reg __425921_425921;
   reg _425922_425922 ; 
   reg __425922_425922;
   reg _425923_425923 ; 
   reg __425923_425923;
   reg _425924_425924 ; 
   reg __425924_425924;
   reg _425925_425925 ; 
   reg __425925_425925;
   reg _425926_425926 ; 
   reg __425926_425926;
   reg _425927_425927 ; 
   reg __425927_425927;
   reg _425928_425928 ; 
   reg __425928_425928;
   reg _425929_425929 ; 
   reg __425929_425929;
   reg _425930_425930 ; 
   reg __425930_425930;
   reg _425931_425931 ; 
   reg __425931_425931;
   reg _425932_425932 ; 
   reg __425932_425932;
   reg _425933_425933 ; 
   reg __425933_425933;
   reg _425934_425934 ; 
   reg __425934_425934;
   reg _425935_425935 ; 
   reg __425935_425935;
   reg _425936_425936 ; 
   reg __425936_425936;
   reg _425937_425937 ; 
   reg __425937_425937;
   reg _425938_425938 ; 
   reg __425938_425938;
   reg _425939_425939 ; 
   reg __425939_425939;
   reg _425940_425940 ; 
   reg __425940_425940;
   reg _425941_425941 ; 
   reg __425941_425941;
   reg _425942_425942 ; 
   reg __425942_425942;
   reg _425943_425943 ; 
   reg __425943_425943;
   reg _425944_425944 ; 
   reg __425944_425944;
   reg _425945_425945 ; 
   reg __425945_425945;
   reg _425946_425946 ; 
   reg __425946_425946;
   reg _425947_425947 ; 
   reg __425947_425947;
   reg _425948_425948 ; 
   reg __425948_425948;
   reg _425949_425949 ; 
   reg __425949_425949;
   reg _425950_425950 ; 
   reg __425950_425950;
   reg _425951_425951 ; 
   reg __425951_425951;
   reg _425952_425952 ; 
   reg __425952_425952;
   reg _425953_425953 ; 
   reg __425953_425953;
   reg _425954_425954 ; 
   reg __425954_425954;
   reg _425955_425955 ; 
   reg __425955_425955;
   reg _425956_425956 ; 
   reg __425956_425956;
   reg _425957_425957 ; 
   reg __425957_425957;
   reg _425958_425958 ; 
   reg __425958_425958;
   reg _425959_425959 ; 
   reg __425959_425959;
   reg _425960_425960 ; 
   reg __425960_425960;
   reg _425961_425961 ; 
   reg __425961_425961;
   reg _425962_425962 ; 
   reg __425962_425962;
   reg _425963_425963 ; 
   reg __425963_425963;
   reg _425964_425964 ; 
   reg __425964_425964;
   reg _425965_425965 ; 
   reg __425965_425965;
   reg _425966_425966 ; 
   reg __425966_425966;
   reg _425967_425967 ; 
   reg __425967_425967;
   reg _425968_425968 ; 
   reg __425968_425968;
   reg _425969_425969 ; 
   reg __425969_425969;
   reg _425970_425970 ; 
   reg __425970_425970;
   reg _425971_425971 ; 
   reg __425971_425971;
   reg _425972_425972 ; 
   reg __425972_425972;
   reg _425973_425973 ; 
   reg __425973_425973;
   reg _425974_425974 ; 
   reg __425974_425974;
   reg _425975_425975 ; 
   reg __425975_425975;
   reg _425976_425976 ; 
   reg __425976_425976;
   reg _425977_425977 ; 
   reg __425977_425977;
   reg _425978_425978 ; 
   reg __425978_425978;
   reg _425979_425979 ; 
   reg __425979_425979;
   reg _425980_425980 ; 
   reg __425980_425980;
   reg _425981_425981 ; 
   reg __425981_425981;
   reg _425982_425982 ; 
   reg __425982_425982;
   reg _425983_425983 ; 
   reg __425983_425983;
   reg _425984_425984 ; 
   reg __425984_425984;
   reg _425985_425985 ; 
   reg __425985_425985;
   reg _425986_425986 ; 
   reg __425986_425986;
   reg _425987_425987 ; 
   reg __425987_425987;
   reg _425988_425988 ; 
   reg __425988_425988;
   reg _425989_425989 ; 
   reg __425989_425989;
   reg _425990_425990 ; 
   reg __425990_425990;
   reg _425991_425991 ; 
   reg __425991_425991;
   reg _425992_425992 ; 
   reg __425992_425992;
   reg _425993_425993 ; 
   reg __425993_425993;
   reg _425994_425994 ; 
   reg __425994_425994;
   reg _425995_425995 ; 
   reg __425995_425995;
   reg _425996_425996 ; 
   reg __425996_425996;
   reg _425997_425997 ; 
   reg __425997_425997;
   reg _425998_425998 ; 
   reg __425998_425998;
   reg _425999_425999 ; 
   reg __425999_425999;
   reg _426000_426000 ; 
   reg __426000_426000;
   reg _426001_426001 ; 
   reg __426001_426001;
   reg _426002_426002 ; 
   reg __426002_426002;
   reg _426003_426003 ; 
   reg __426003_426003;
   reg _426004_426004 ; 
   reg __426004_426004;
   reg _426005_426005 ; 
   reg __426005_426005;
   reg _426006_426006 ; 
   reg __426006_426006;
   reg _426007_426007 ; 
   reg __426007_426007;
   reg _426008_426008 ; 
   reg __426008_426008;
   reg _426009_426009 ; 
   reg __426009_426009;
   reg _426010_426010 ; 
   reg __426010_426010;
   reg _426011_426011 ; 
   reg __426011_426011;
   reg _426012_426012 ; 
   reg __426012_426012;
   reg _426013_426013 ; 
   reg __426013_426013;
   reg _426014_426014 ; 
   reg __426014_426014;
   reg _426015_426015 ; 
   reg __426015_426015;
   reg _426016_426016 ; 
   reg __426016_426016;
   reg _426017_426017 ; 
   reg __426017_426017;
   reg _426018_426018 ; 
   reg __426018_426018;
   reg _426019_426019 ; 
   reg __426019_426019;
   reg _426020_426020 ; 
   reg __426020_426020;
   reg _426021_426021 ; 
   reg __426021_426021;
   reg _426022_426022 ; 
   reg __426022_426022;
   reg _426023_426023 ; 
   reg __426023_426023;
   reg _426024_426024 ; 
   reg __426024_426024;
   reg _426025_426025 ; 
   reg __426025_426025;
   reg _426026_426026 ; 
   reg __426026_426026;
   reg _426027_426027 ; 
   reg __426027_426027;
   reg _426028_426028 ; 
   reg __426028_426028;
   reg _426029_426029 ; 
   reg __426029_426029;
   reg _426030_426030 ; 
   reg __426030_426030;
   reg _426031_426031 ; 
   reg __426031_426031;
   reg _426032_426032 ; 
   reg __426032_426032;
   reg _426033_426033 ; 
   reg __426033_426033;
   reg _426034_426034 ; 
   reg __426034_426034;
   reg _426035_426035 ; 
   reg __426035_426035;
   reg _426036_426036 ; 
   reg __426036_426036;
   reg _426037_426037 ; 
   reg __426037_426037;
   reg _426038_426038 ; 
   reg __426038_426038;
   reg _426039_426039 ; 
   reg __426039_426039;
   reg _426040_426040 ; 
   reg __426040_426040;
   reg _426041_426041 ; 
   reg __426041_426041;
   reg _426042_426042 ; 
   reg __426042_426042;
   reg _426043_426043 ; 
   reg __426043_426043;
   reg _426044_426044 ; 
   reg __426044_426044;
   reg _426045_426045 ; 
   reg __426045_426045;
   reg _426046_426046 ; 
   reg __426046_426046;
   reg _426047_426047 ; 
   reg __426047_426047;
   reg _426048_426048 ; 
   reg __426048_426048;
   reg _426049_426049 ; 
   reg __426049_426049;
   reg _426050_426050 ; 
   reg __426050_426050;
   reg _426051_426051 ; 
   reg __426051_426051;
   reg _426052_426052 ; 
   reg __426052_426052;
   reg _426053_426053 ; 
   reg __426053_426053;
   reg _426054_426054 ; 
   reg __426054_426054;
   reg _426055_426055 ; 
   reg __426055_426055;
   reg _426056_426056 ; 
   reg __426056_426056;
   reg _426057_426057 ; 
   reg __426057_426057;
   reg _426058_426058 ; 
   reg __426058_426058;
   reg _426059_426059 ; 
   reg __426059_426059;
   reg _426060_426060 ; 
   reg __426060_426060;
   reg _426061_426061 ; 
   reg __426061_426061;
   reg _426062_426062 ; 
   reg __426062_426062;
   reg _426063_426063 ; 
   reg __426063_426063;
   reg _426064_426064 ; 
   reg __426064_426064;
   reg _426065_426065 ; 
   reg __426065_426065;
   reg _426066_426066 ; 
   reg __426066_426066;
   reg _426067_426067 ; 
   reg __426067_426067;
   reg _426068_426068 ; 
   reg __426068_426068;
   reg _426069_426069 ; 
   reg __426069_426069;
   reg _426070_426070 ; 
   reg __426070_426070;
   reg _426071_426071 ; 
   reg __426071_426071;
   reg _426072_426072 ; 
   reg __426072_426072;
   reg _426073_426073 ; 
   reg __426073_426073;
   reg _426074_426074 ; 
   reg __426074_426074;
   reg _426075_426075 ; 
   reg __426075_426075;
   reg _426076_426076 ; 
   reg __426076_426076;
   reg _426077_426077 ; 
   reg __426077_426077;
   reg _426078_426078 ; 
   reg __426078_426078;
   reg _426079_426079 ; 
   reg __426079_426079;
   reg _426080_426080 ; 
   reg __426080_426080;
   reg _426081_426081 ; 
   reg __426081_426081;
   reg _426082_426082 ; 
   reg __426082_426082;
   reg _426083_426083 ; 
   reg __426083_426083;
   reg _426084_426084 ; 
   reg __426084_426084;
   reg _426085_426085 ; 
   reg __426085_426085;
   reg _426086_426086 ; 
   reg __426086_426086;
   reg _426087_426087 ; 
   reg __426087_426087;
   reg _426088_426088 ; 
   reg __426088_426088;
   reg _426089_426089 ; 
   reg __426089_426089;
   reg _426090_426090 ; 
   reg __426090_426090;
   reg _426091_426091 ; 
   reg __426091_426091;
   reg _426092_426092 ; 
   reg __426092_426092;
   reg _426093_426093 ; 
   reg __426093_426093;
   reg _426094_426094 ; 
   reg __426094_426094;
   reg _426095_426095 ; 
   reg __426095_426095;
   reg _426096_426096 ; 
   reg __426096_426096;
   reg _426097_426097 ; 
   reg __426097_426097;
   reg _426098_426098 ; 
   reg __426098_426098;
   reg _426099_426099 ; 
   reg __426099_426099;
   reg _426100_426100 ; 
   reg __426100_426100;
   reg _426101_426101 ; 
   reg __426101_426101;
   reg _426102_426102 ; 
   reg __426102_426102;
   reg _426103_426103 ; 
   reg __426103_426103;
   reg _426104_426104 ; 
   reg __426104_426104;
   reg _426105_426105 ; 
   reg __426105_426105;
   reg _426106_426106 ; 
   reg __426106_426106;
   reg _426107_426107 ; 
   reg __426107_426107;
   reg _426108_426108 ; 
   reg __426108_426108;
   reg _426109_426109 ; 
   reg __426109_426109;
   reg _426110_426110 ; 
   reg __426110_426110;
   reg _426111_426111 ; 
   reg __426111_426111;
   reg _426112_426112 ; 
   reg __426112_426112;
   reg _426113_426113 ; 
   reg __426113_426113;
   reg _426114_426114 ; 
   reg __426114_426114;
   reg _426115_426115 ; 
   reg __426115_426115;
   reg _426116_426116 ; 
   reg __426116_426116;
   reg _426117_426117 ; 
   reg __426117_426117;
   reg _426118_426118 ; 
   reg __426118_426118;
   reg _426119_426119 ; 
   reg __426119_426119;
   reg _426120_426120 ; 
   reg __426120_426120;
   reg _426121_426121 ; 
   reg __426121_426121;
   reg _426122_426122 ; 
   reg __426122_426122;
   reg _426123_426123 ; 
   reg __426123_426123;
   reg _426124_426124 ; 
   reg __426124_426124;
   reg _426125_426125 ; 
   reg __426125_426125;
   reg _426126_426126 ; 
   reg __426126_426126;
   reg _426127_426127 ; 
   reg __426127_426127;
   reg _426128_426128 ; 
   reg __426128_426128;
   reg _426129_426129 ; 
   reg __426129_426129;
   reg _426130_426130 ; 
   reg __426130_426130;
   reg _426131_426131 ; 
   reg __426131_426131;
   reg _426132_426132 ; 
   reg __426132_426132;
   reg _426133_426133 ; 
   reg __426133_426133;
   reg _426134_426134 ; 
   reg __426134_426134;
   reg _426135_426135 ; 
   reg __426135_426135;
   reg _426136_426136 ; 
   reg __426136_426136;
   reg _426137_426137 ; 
   reg __426137_426137;
   reg _426138_426138 ; 
   reg __426138_426138;
   reg _426139_426139 ; 
   reg __426139_426139;
   reg _426140_426140 ; 
   reg __426140_426140;
   reg _426141_426141 ; 
   reg __426141_426141;
   reg _426142_426142 ; 
   reg __426142_426142;
   reg _426143_426143 ; 
   reg __426143_426143;
   reg _426144_426144 ; 
   reg __426144_426144;
   reg _426145_426145 ; 
   reg __426145_426145;
   reg _426146_426146 ; 
   reg __426146_426146;
   reg _426147_426147 ; 
   reg __426147_426147;
   reg _426148_426148 ; 
   reg __426148_426148;
   reg _426149_426149 ; 
   reg __426149_426149;
   reg _426150_426150 ; 
   reg __426150_426150;
   reg _426151_426151 ; 
   reg __426151_426151;
   reg _426152_426152 ; 
   reg __426152_426152;
   reg _426153_426153 ; 
   reg __426153_426153;
   reg _426154_426154 ; 
   reg __426154_426154;
   reg _426155_426155 ; 
   reg __426155_426155;
   reg _426156_426156 ; 
   reg __426156_426156;
   reg _426157_426157 ; 
   reg __426157_426157;
   reg _426158_426158 ; 
   reg __426158_426158;
   reg _426159_426159 ; 
   reg __426159_426159;
   reg _426160_426160 ; 
   reg __426160_426160;
   reg _426161_426161 ; 
   reg __426161_426161;
   reg _426162_426162 ; 
   reg __426162_426162;
   reg _426163_426163 ; 
   reg __426163_426163;
   reg _426164_426164 ; 
   reg __426164_426164;
   reg _426165_426165 ; 
   reg __426165_426165;
   reg _426166_426166 ; 
   reg __426166_426166;
   reg _426167_426167 ; 
   reg __426167_426167;
   reg _426168_426168 ; 
   reg __426168_426168;
   reg _426169_426169 ; 
   reg __426169_426169;
   reg _426170_426170 ; 
   reg __426170_426170;
   reg _426171_426171 ; 
   reg __426171_426171;
   reg _426172_426172 ; 
   reg __426172_426172;
   reg _426173_426173 ; 
   reg __426173_426173;
   reg _426174_426174 ; 
   reg __426174_426174;
   reg _426175_426175 ; 
   reg __426175_426175;
   reg _426176_426176 ; 
   reg __426176_426176;
   reg _426177_426177 ; 
   reg __426177_426177;
   reg _426178_426178 ; 
   reg __426178_426178;
   reg _426179_426179 ; 
   reg __426179_426179;
   reg _426180_426180 ; 
   reg __426180_426180;
   reg _426181_426181 ; 
   reg __426181_426181;
   reg _426182_426182 ; 
   reg __426182_426182;
   reg _426183_426183 ; 
   reg __426183_426183;
   reg _426184_426184 ; 
   reg __426184_426184;
   reg _426185_426185 ; 
   reg __426185_426185;
   reg _426186_426186 ; 
   reg __426186_426186;
   reg _426187_426187 ; 
   reg __426187_426187;
   reg _426188_426188 ; 
   reg __426188_426188;
   reg _426189_426189 ; 
   reg __426189_426189;
   reg _426190_426190 ; 
   reg __426190_426190;
   reg _426191_426191 ; 
   reg __426191_426191;
   reg _426192_426192 ; 
   reg __426192_426192;
   reg _426193_426193 ; 
   reg __426193_426193;
   reg _426194_426194 ; 
   reg __426194_426194;
   reg _426195_426195 ; 
   reg __426195_426195;
   reg _426196_426196 ; 
   reg __426196_426196;
   reg _426197_426197 ; 
   reg __426197_426197;
   reg _426198_426198 ; 
   reg __426198_426198;
   reg _426199_426199 ; 
   reg __426199_426199;
   reg _426200_426200 ; 
   reg __426200_426200;
   reg _426201_426201 ; 
   reg __426201_426201;
   reg _426202_426202 ; 
   reg __426202_426202;
   reg _426203_426203 ; 
   reg __426203_426203;
   reg _426204_426204 ; 
   reg __426204_426204;
   reg _426205_426205 ; 
   reg __426205_426205;
   reg _426206_426206 ; 
   reg __426206_426206;
   reg _426207_426207 ; 
   reg __426207_426207;
   reg _426208_426208 ; 
   reg __426208_426208;
   reg _426209_426209 ; 
   reg __426209_426209;
   reg _426210_426210 ; 
   reg __426210_426210;
   reg _426211_426211 ; 
   reg __426211_426211;
   reg _426212_426212 ; 
   reg __426212_426212;
   reg _426213_426213 ; 
   reg __426213_426213;
   reg _426214_426214 ; 
   reg __426214_426214;
   reg _426215_426215 ; 
   reg __426215_426215;
   reg _426216_426216 ; 
   reg __426216_426216;
   reg _426217_426217 ; 
   reg __426217_426217;
   reg _426218_426218 ; 
   reg __426218_426218;
   reg _426219_426219 ; 
   reg __426219_426219;
   reg _426220_426220 ; 
   reg __426220_426220;
   reg _426221_426221 ; 
   reg __426221_426221;
   reg _426222_426222 ; 
   reg __426222_426222;
   reg _426223_426223 ; 
   reg __426223_426223;
   reg _426224_426224 ; 
   reg __426224_426224;
   reg _426225_426225 ; 
   reg __426225_426225;
   reg _426226_426226 ; 
   reg __426226_426226;
   reg _426227_426227 ; 
   reg __426227_426227;
   reg _426228_426228 ; 
   reg __426228_426228;
   reg _426229_426229 ; 
   reg __426229_426229;
   reg _426230_426230 ; 
   reg __426230_426230;
   reg _426231_426231 ; 
   reg __426231_426231;
   reg _426232_426232 ; 
   reg __426232_426232;
   reg _426233_426233 ; 
   reg __426233_426233;
   reg _426234_426234 ; 
   reg __426234_426234;
   reg _426235_426235 ; 
   reg __426235_426235;
   reg _426236_426236 ; 
   reg __426236_426236;
   reg _426237_426237 ; 
   reg __426237_426237;
   reg _426238_426238 ; 
   reg __426238_426238;
   reg _426239_426239 ; 
   reg __426239_426239;
   reg _426240_426240 ; 
   reg __426240_426240;
   reg _426241_426241 ; 
   reg __426241_426241;
   reg _426242_426242 ; 
   reg __426242_426242;
   reg _426243_426243 ; 
   reg __426243_426243;
   reg _426244_426244 ; 
   reg __426244_426244;
   reg _426245_426245 ; 
   reg __426245_426245;
   reg _426246_426246 ; 
   reg __426246_426246;
   reg _426247_426247 ; 
   reg __426247_426247;
   reg _426248_426248 ; 
   reg __426248_426248;
   reg _426249_426249 ; 
   reg __426249_426249;
   reg _426250_426250 ; 
   reg __426250_426250;
   reg _426251_426251 ; 
   reg __426251_426251;
   reg _426252_426252 ; 
   reg __426252_426252;
   reg _426253_426253 ; 
   reg __426253_426253;
   reg _426254_426254 ; 
   reg __426254_426254;
   reg _426255_426255 ; 
   reg __426255_426255;
   reg _426256_426256 ; 
   reg __426256_426256;
   reg _426257_426257 ; 
   reg __426257_426257;
   reg _426258_426258 ; 
   reg __426258_426258;
   reg _426259_426259 ; 
   reg __426259_426259;
   reg _426260_426260 ; 
   reg __426260_426260;
   reg _426261_426261 ; 
   reg __426261_426261;
   reg _426262_426262 ; 
   reg __426262_426262;
   reg _426263_426263 ; 
   reg __426263_426263;
   reg _426264_426264 ; 
   reg __426264_426264;
   reg _426265_426265 ; 
   reg __426265_426265;
   reg _426266_426266 ; 
   reg __426266_426266;
   reg _426267_426267 ; 
   reg __426267_426267;
   reg _426268_426268 ; 
   reg __426268_426268;
   reg _426269_426269 ; 
   reg __426269_426269;
   reg _426270_426270 ; 
   reg __426270_426270;
   reg _426271_426271 ; 
   reg __426271_426271;
   reg _426272_426272 ; 
   reg __426272_426272;
   reg _426273_426273 ; 
   reg __426273_426273;
   reg _426274_426274 ; 
   reg __426274_426274;
   reg _426275_426275 ; 
   reg __426275_426275;
   reg _426276_426276 ; 
   reg __426276_426276;
   reg _426277_426277 ; 
   reg __426277_426277;
   reg _426278_426278 ; 
   reg __426278_426278;
   reg _426279_426279 ; 
   reg __426279_426279;
   reg _426280_426280 ; 
   reg __426280_426280;
   reg _426281_426281 ; 
   reg __426281_426281;
   reg _426282_426282 ; 
   reg __426282_426282;
   reg _426283_426283 ; 
   reg __426283_426283;
   reg _426284_426284 ; 
   reg __426284_426284;
   reg _426285_426285 ; 
   reg __426285_426285;
   reg _426286_426286 ; 
   reg __426286_426286;
   reg _426287_426287 ; 
   reg __426287_426287;
   reg _426288_426288 ; 
   reg __426288_426288;
   reg _426289_426289 ; 
   reg __426289_426289;
   reg _426290_426290 ; 
   reg __426290_426290;
   reg _426291_426291 ; 
   reg __426291_426291;
   reg _426292_426292 ; 
   reg __426292_426292;
   reg _426293_426293 ; 
   reg __426293_426293;
   reg _426294_426294 ; 
   reg __426294_426294;
   reg _426295_426295 ; 
   reg __426295_426295;
   reg _426296_426296 ; 
   reg __426296_426296;
   reg _426297_426297 ; 
   reg __426297_426297;
   reg _426298_426298 ; 
   reg __426298_426298;
   reg _426299_426299 ; 
   reg __426299_426299;
   reg _426300_426300 ; 
   reg __426300_426300;
   reg _426301_426301 ; 
   reg __426301_426301;
   reg _426302_426302 ; 
   reg __426302_426302;
   reg _426303_426303 ; 
   reg __426303_426303;
   reg _426304_426304 ; 
   reg __426304_426304;
   reg _426305_426305 ; 
   reg __426305_426305;
   reg _426306_426306 ; 
   reg __426306_426306;
   reg _426307_426307 ; 
   reg __426307_426307;
   reg _426308_426308 ; 
   reg __426308_426308;
   reg _426309_426309 ; 
   reg __426309_426309;
   reg _426310_426310 ; 
   reg __426310_426310;
   reg _426311_426311 ; 
   reg __426311_426311;
   reg _426312_426312 ; 
   reg __426312_426312;
   reg _426313_426313 ; 
   reg __426313_426313;
   reg _426314_426314 ; 
   reg __426314_426314;
   reg _426315_426315 ; 
   reg __426315_426315;
   reg _426316_426316 ; 
   reg __426316_426316;
   reg _426317_426317 ; 
   reg __426317_426317;
   reg _426318_426318 ; 
   reg __426318_426318;
   reg _426319_426319 ; 
   reg __426319_426319;
   reg _426320_426320 ; 
   reg __426320_426320;
   reg _426321_426321 ; 
   reg __426321_426321;
   reg _426322_426322 ; 
   reg __426322_426322;
   reg _426323_426323 ; 
   reg __426323_426323;
   reg _426324_426324 ; 
   reg __426324_426324;
   reg _426325_426325 ; 
   reg __426325_426325;
   reg _426326_426326 ; 
   reg __426326_426326;
   reg _426327_426327 ; 
   reg __426327_426327;
   reg _426328_426328 ; 
   reg __426328_426328;
   reg _426329_426329 ; 
   reg __426329_426329;
   reg _426330_426330 ; 
   reg __426330_426330;
   reg _426331_426331 ; 
   reg __426331_426331;
   reg _426332_426332 ; 
   reg __426332_426332;
   reg _426333_426333 ; 
   reg __426333_426333;
   reg _426334_426334 ; 
   reg __426334_426334;
   reg _426335_426335 ; 
   reg __426335_426335;
   reg _426336_426336 ; 
   reg __426336_426336;
   reg _426337_426337 ; 
   reg __426337_426337;
   reg _426338_426338 ; 
   reg __426338_426338;
   reg _426339_426339 ; 
   reg __426339_426339;
   reg _426340_426340 ; 
   reg __426340_426340;
   reg _426341_426341 ; 
   reg __426341_426341;
   reg _426342_426342 ; 
   reg __426342_426342;
   reg _426343_426343 ; 
   reg __426343_426343;
   reg _426344_426344 ; 
   reg __426344_426344;
   reg _426345_426345 ; 
   reg __426345_426345;
   reg _426346_426346 ; 
   reg __426346_426346;
   reg _426347_426347 ; 
   reg __426347_426347;
   reg _426348_426348 ; 
   reg __426348_426348;
   reg _426349_426349 ; 
   reg __426349_426349;
   reg _426350_426350 ; 
   reg __426350_426350;
   reg _426351_426351 ; 
   reg __426351_426351;
   reg _426352_426352 ; 
   reg __426352_426352;
   reg _426353_426353 ; 
   reg __426353_426353;
   reg _426354_426354 ; 
   reg __426354_426354;
   reg _426355_426355 ; 
   reg __426355_426355;
   reg _426356_426356 ; 
   reg __426356_426356;
   reg _426357_426357 ; 
   reg __426357_426357;
   reg _426358_426358 ; 
   reg __426358_426358;
   reg _426359_426359 ; 
   reg __426359_426359;
   reg _426360_426360 ; 
   reg __426360_426360;
   reg _426361_426361 ; 
   reg __426361_426361;
   reg _426362_426362 ; 
   reg __426362_426362;
   reg _426363_426363 ; 
   reg __426363_426363;
   reg _426364_426364 ; 
   reg __426364_426364;
   reg _426365_426365 ; 
   reg __426365_426365;
   reg _426366_426366 ; 
   reg __426366_426366;
   reg _426367_426367 ; 
   reg __426367_426367;
   reg _426368_426368 ; 
   reg __426368_426368;
   reg _426369_426369 ; 
   reg __426369_426369;
   reg _426370_426370 ; 
   reg __426370_426370;
   reg _426371_426371 ; 
   reg __426371_426371;
   reg _426372_426372 ; 
   reg __426372_426372;
   reg _426373_426373 ; 
   reg __426373_426373;
   reg _426374_426374 ; 
   reg __426374_426374;
   reg _426375_426375 ; 
   reg __426375_426375;
   reg _426376_426376 ; 
   reg __426376_426376;
   reg _426377_426377 ; 
   reg __426377_426377;
   reg _426378_426378 ; 
   reg __426378_426378;
   reg _426379_426379 ; 
   reg __426379_426379;
   reg _426380_426380 ; 
   reg __426380_426380;
   reg _426381_426381 ; 
   reg __426381_426381;
   reg _426382_426382 ; 
   reg __426382_426382;
   reg _426383_426383 ; 
   reg __426383_426383;
   reg _426384_426384 ; 
   reg __426384_426384;
   reg _426385_426385 ; 
   reg __426385_426385;
   reg _426386_426386 ; 
   reg __426386_426386;
   reg _426387_426387 ; 
   reg __426387_426387;
   reg _426388_426388 ; 
   reg __426388_426388;
   reg _426389_426389 ; 
   reg __426389_426389;
   reg _426390_426390 ; 
   reg __426390_426390;
   reg _426391_426391 ; 
   reg __426391_426391;
   reg _426392_426392 ; 
   reg __426392_426392;
   reg _426393_426393 ; 
   reg __426393_426393;
   reg _426394_426394 ; 
   reg __426394_426394;
   reg _426395_426395 ; 
   reg __426395_426395;
   reg _426396_426396 ; 
   reg __426396_426396;
   reg _426397_426397 ; 
   reg __426397_426397;
   reg _426398_426398 ; 
   reg __426398_426398;
   reg _426399_426399 ; 
   reg __426399_426399;
   reg _426400_426400 ; 
   reg __426400_426400;
   reg _426401_426401 ; 
   reg __426401_426401;
   reg _426402_426402 ; 
   reg __426402_426402;
   reg _426403_426403 ; 
   reg __426403_426403;
   reg _426404_426404 ; 
   reg __426404_426404;
   reg _426405_426405 ; 
   reg __426405_426405;
   reg _426406_426406 ; 
   reg __426406_426406;
   reg _426407_426407 ; 
   reg __426407_426407;
   reg _426408_426408 ; 
   reg __426408_426408;
   reg _426409_426409 ; 
   reg __426409_426409;
   reg _426410_426410 ; 
   reg __426410_426410;
   reg _426411_426411 ; 
   reg __426411_426411;
   reg _426412_426412 ; 
   reg __426412_426412;
   reg _426413_426413 ; 
   reg __426413_426413;
   reg _426414_426414 ; 
   reg __426414_426414;
   reg _426415_426415 ; 
   reg __426415_426415;
   reg _426416_426416 ; 
   reg __426416_426416;
   reg _426417_426417 ; 
   reg __426417_426417;
   reg _426418_426418 ; 
   reg __426418_426418;
   reg _426419_426419 ; 
   reg __426419_426419;
   reg _426420_426420 ; 
   reg __426420_426420;
   reg _426421_426421 ; 
   reg __426421_426421;
   reg _426422_426422 ; 
   reg __426422_426422;
   reg _426423_426423 ; 
   reg __426423_426423;
   reg _426424_426424 ; 
   reg __426424_426424;
   reg _426425_426425 ; 
   reg __426425_426425;
   reg _426426_426426 ; 
   reg __426426_426426;
   reg _426427_426427 ; 
   reg __426427_426427;
   reg _426428_426428 ; 
   reg __426428_426428;
   reg _426429_426429 ; 
   reg __426429_426429;
   reg _426430_426430 ; 
   reg __426430_426430;
   reg _426431_426431 ; 
   reg __426431_426431;
   reg _426432_426432 ; 
   reg __426432_426432;
   reg _426433_426433 ; 
   reg __426433_426433;
   reg _426434_426434 ; 
   reg __426434_426434;
   reg _426435_426435 ; 
   reg __426435_426435;
   reg _426436_426436 ; 
   reg __426436_426436;
   reg _426437_426437 ; 
   reg __426437_426437;
   reg _426438_426438 ; 
   reg __426438_426438;
   reg _426439_426439 ; 
   reg __426439_426439;
   reg _426440_426440 ; 
   reg __426440_426440;
   reg _426441_426441 ; 
   reg __426441_426441;
   reg _426442_426442 ; 
   reg __426442_426442;
   reg _426443_426443 ; 
   reg __426443_426443;
   reg _426444_426444 ; 
   reg __426444_426444;
   reg _426445_426445 ; 
   reg __426445_426445;
   reg _426446_426446 ; 
   reg __426446_426446;
   reg _426447_426447 ; 
   reg __426447_426447;
   reg _426448_426448 ; 
   reg __426448_426448;
   reg _426449_426449 ; 
   reg __426449_426449;
   reg _426450_426450 ; 
   reg __426450_426450;
   reg _426451_426451 ; 
   reg __426451_426451;
   reg _426452_426452 ; 
   reg __426452_426452;
   reg _426453_426453 ; 
   reg __426453_426453;
   reg _426454_426454 ; 
   reg __426454_426454;
   reg _426455_426455 ; 
   reg __426455_426455;
   reg _426456_426456 ; 
   reg __426456_426456;
   reg _426457_426457 ; 
   reg __426457_426457;
   reg _426458_426458 ; 
   reg __426458_426458;
   reg _426459_426459 ; 
   reg __426459_426459;
   reg _426460_426460 ; 
   reg __426460_426460;
   reg _426461_426461 ; 
   reg __426461_426461;
   reg _426462_426462 ; 
   reg __426462_426462;
   reg _426463_426463 ; 
   reg __426463_426463;
   reg _426464_426464 ; 
   reg __426464_426464;
   reg _426465_426465 ; 
   reg __426465_426465;
   reg _426466_426466 ; 
   reg __426466_426466;
   reg _426467_426467 ; 
   reg __426467_426467;
   reg _426468_426468 ; 
   reg __426468_426468;
   reg _426469_426469 ; 
   reg __426469_426469;
   reg _426470_426470 ; 
   reg __426470_426470;
   reg _426471_426471 ; 
   reg __426471_426471;
   reg _426472_426472 ; 
   reg __426472_426472;
   reg _426473_426473 ; 
   reg __426473_426473;
   reg _426474_426474 ; 
   reg __426474_426474;
   reg _426475_426475 ; 
   reg __426475_426475;
   reg _426476_426476 ; 
   reg __426476_426476;
   reg _426477_426477 ; 
   reg __426477_426477;
   reg _426478_426478 ; 
   reg __426478_426478;
   reg _426479_426479 ; 
   reg __426479_426479;
   reg _426480_426480 ; 
   reg __426480_426480;
   reg _426481_426481 ; 
   reg __426481_426481;
   reg _426482_426482 ; 
   reg __426482_426482;
   reg _426483_426483 ; 
   reg __426483_426483;
   reg _426484_426484 ; 
   reg __426484_426484;
   reg _426485_426485 ; 
   reg __426485_426485;
   reg _426486_426486 ; 
   reg __426486_426486;
   reg _426487_426487 ; 
   reg __426487_426487;
   reg _426488_426488 ; 
   reg __426488_426488;
   reg _426489_426489 ; 
   reg __426489_426489;
   reg _426490_426490 ; 
   reg __426490_426490;
   reg _426491_426491 ; 
   reg __426491_426491;
   reg _426492_426492 ; 
   reg __426492_426492;
   reg _426493_426493 ; 
   reg __426493_426493;
   reg _426494_426494 ; 
   reg __426494_426494;
   reg _426495_426495 ; 
   reg __426495_426495;
   reg _426496_426496 ; 
   reg __426496_426496;
   reg _426497_426497 ; 
   reg __426497_426497;
   reg _426498_426498 ; 
   reg __426498_426498;
   reg _426499_426499 ; 
   reg __426499_426499;
   reg _426500_426500 ; 
   reg __426500_426500;
   reg _426501_426501 ; 
   reg __426501_426501;
   reg _426502_426502 ; 
   reg __426502_426502;
   reg _426503_426503 ; 
   reg __426503_426503;
   reg _426504_426504 ; 
   reg __426504_426504;
   reg _426505_426505 ; 
   reg __426505_426505;
   reg _426506_426506 ; 
   reg __426506_426506;
   reg _426507_426507 ; 
   reg __426507_426507;
   reg _426508_426508 ; 
   reg __426508_426508;
   reg _426509_426509 ; 
   reg __426509_426509;
   reg _426510_426510 ; 
   reg __426510_426510;
   reg _426511_426511 ; 
   reg __426511_426511;
   reg _426512_426512 ; 
   reg __426512_426512;
   reg _426513_426513 ; 
   reg __426513_426513;
   reg _426514_426514 ; 
   reg __426514_426514;
   reg _426515_426515 ; 
   reg __426515_426515;
   reg _426516_426516 ; 
   reg __426516_426516;
   reg _426517_426517 ; 
   reg __426517_426517;
   reg _426518_426518 ; 
   reg __426518_426518;
   reg _426519_426519 ; 
   reg __426519_426519;
   reg _426520_426520 ; 
   reg __426520_426520;
   reg _426521_426521 ; 
   reg __426521_426521;
   reg _426522_426522 ; 
   reg __426522_426522;
   reg _426523_426523 ; 
   reg __426523_426523;
   reg _426524_426524 ; 
   reg __426524_426524;
   reg _426525_426525 ; 
   reg __426525_426525;
   reg _426526_426526 ; 
   reg __426526_426526;
   reg _426527_426527 ; 
   reg __426527_426527;
   reg _426528_426528 ; 
   reg __426528_426528;
   reg _426529_426529 ; 
   reg __426529_426529;
   reg _426530_426530 ; 
   reg __426530_426530;
   reg _426531_426531 ; 
   reg __426531_426531;
   reg _426532_426532 ; 
   reg __426532_426532;
   reg _426533_426533 ; 
   reg __426533_426533;
   reg _426534_426534 ; 
   reg __426534_426534;
   reg _426535_426535 ; 
   reg __426535_426535;
   reg _426536_426536 ; 
   reg __426536_426536;
   reg _426537_426537 ; 
   reg __426537_426537;
   reg _426538_426538 ; 
   reg __426538_426538;
   reg _426539_426539 ; 
   reg __426539_426539;
   reg _426540_426540 ; 
   reg __426540_426540;
   reg _426541_426541 ; 
   reg __426541_426541;
   reg _426542_426542 ; 
   reg __426542_426542;
   reg _426543_426543 ; 
   reg __426543_426543;
   reg _426544_426544 ; 
   reg __426544_426544;
   reg _426545_426545 ; 
   reg __426545_426545;
   reg _426546_426546 ; 
   reg __426546_426546;
   reg _426547_426547 ; 
   reg __426547_426547;
   reg _426548_426548 ; 
   reg __426548_426548;
   reg _426549_426549 ; 
   reg __426549_426549;
   reg _426550_426550 ; 
   reg __426550_426550;
   reg _426551_426551 ; 
   reg __426551_426551;
   reg _426552_426552 ; 
   reg __426552_426552;
   reg _426553_426553 ; 
   reg __426553_426553;
   reg _426554_426554 ; 
   reg __426554_426554;
   reg _426555_426555 ; 
   reg __426555_426555;
   reg _426556_426556 ; 
   reg __426556_426556;
   reg _426557_426557 ; 
   reg __426557_426557;
   reg _426558_426558 ; 
   reg __426558_426558;
   reg _426559_426559 ; 
   reg __426559_426559;
   reg _426560_426560 ; 
   reg __426560_426560;
   reg _426561_426561 ; 
   reg __426561_426561;
   reg _426562_426562 ; 
   reg __426562_426562;
   reg _426563_426563 ; 
   reg __426563_426563;
   reg _426564_426564 ; 
   reg __426564_426564;
   reg _426565_426565 ; 
   reg __426565_426565;
   reg _426566_426566 ; 
   reg __426566_426566;
   reg _426567_426567 ; 
   reg __426567_426567;
   reg _426568_426568 ; 
   reg __426568_426568;
   reg _426569_426569 ; 
   reg __426569_426569;
   reg _426570_426570 ; 
   reg __426570_426570;
   reg _426571_426571 ; 
   reg __426571_426571;
   reg _426572_426572 ; 
   reg __426572_426572;
   reg _426573_426573 ; 
   reg __426573_426573;
   reg _426574_426574 ; 
   reg __426574_426574;
   reg _426575_426575 ; 
   reg __426575_426575;
   reg _426576_426576 ; 
   reg __426576_426576;
   reg _426577_426577 ; 
   reg __426577_426577;
   reg _426578_426578 ; 
   reg __426578_426578;
   reg _426579_426579 ; 
   reg __426579_426579;
   reg _426580_426580 ; 
   reg __426580_426580;
   reg _426581_426581 ; 
   reg __426581_426581;
   reg _426582_426582 ; 
   reg __426582_426582;
   reg _426583_426583 ; 
   reg __426583_426583;
   reg _426584_426584 ; 
   reg __426584_426584;
   reg _426585_426585 ; 
   reg __426585_426585;
   reg _426586_426586 ; 
   reg __426586_426586;
   reg _426587_426587 ; 
   reg __426587_426587;
   reg _426588_426588 ; 
   reg __426588_426588;
   reg _426589_426589 ; 
   reg __426589_426589;
   reg _426590_426590 ; 
   reg __426590_426590;
   reg _426591_426591 ; 
   reg __426591_426591;
   reg _426592_426592 ; 
   reg __426592_426592;
   reg _426593_426593 ; 
   reg __426593_426593;
   reg _426594_426594 ; 
   reg __426594_426594;
   reg _426595_426595 ; 
   reg __426595_426595;
   reg _426596_426596 ; 
   reg __426596_426596;
   reg _426597_426597 ; 
   reg __426597_426597;
   reg _426598_426598 ; 
   reg __426598_426598;
   reg _426599_426599 ; 
   reg __426599_426599;
   reg _426600_426600 ; 
   reg __426600_426600;
   reg _426601_426601 ; 
   reg __426601_426601;
   reg _426602_426602 ; 
   reg __426602_426602;
   reg _426603_426603 ; 
   reg __426603_426603;
   reg _426604_426604 ; 
   reg __426604_426604;
   reg _426605_426605 ; 
   reg __426605_426605;
   reg _426606_426606 ; 
   reg __426606_426606;
   reg _426607_426607 ; 
   reg __426607_426607;
   reg _426608_426608 ; 
   reg __426608_426608;
   reg _426609_426609 ; 
   reg __426609_426609;
   reg _426610_426610 ; 
   reg __426610_426610;
   reg _426611_426611 ; 
   reg __426611_426611;
   reg _426612_426612 ; 
   reg __426612_426612;
   reg _426613_426613 ; 
   reg __426613_426613;
   reg _426614_426614 ; 
   reg __426614_426614;
   reg _426615_426615 ; 
   reg __426615_426615;
   reg _426616_426616 ; 
   reg __426616_426616;
   reg _426617_426617 ; 
   reg __426617_426617;
   reg _426618_426618 ; 
   reg __426618_426618;
   reg _426619_426619 ; 
   reg __426619_426619;
   reg _426620_426620 ; 
   reg __426620_426620;
   reg _426621_426621 ; 
   reg __426621_426621;
   reg _426622_426622 ; 
   reg __426622_426622;
   reg _426623_426623 ; 
   reg __426623_426623;
   reg _426624_426624 ; 
   reg __426624_426624;
   reg _426625_426625 ; 
   reg __426625_426625;
   reg _426626_426626 ; 
   reg __426626_426626;
   reg _426627_426627 ; 
   reg __426627_426627;
   reg _426628_426628 ; 
   reg __426628_426628;
   reg _426629_426629 ; 
   reg __426629_426629;
   reg _426630_426630 ; 
   reg __426630_426630;
   reg _426631_426631 ; 
   reg __426631_426631;
   reg _426632_426632 ; 
   reg __426632_426632;
   reg _426633_426633 ; 
   reg __426633_426633;
   reg _426634_426634 ; 
   reg __426634_426634;
   reg _426635_426635 ; 
   reg __426635_426635;
   reg _426636_426636 ; 
   reg __426636_426636;
   reg _426637_426637 ; 
   reg __426637_426637;
   reg _426638_426638 ; 
   reg __426638_426638;
   reg _426639_426639 ; 
   reg __426639_426639;
   reg _426640_426640 ; 
   reg __426640_426640;
   reg _426641_426641 ; 
   reg __426641_426641;
   reg _426642_426642 ; 
   reg __426642_426642;
   reg _426643_426643 ; 
   reg __426643_426643;
   reg _426644_426644 ; 
   reg __426644_426644;
   reg _426645_426645 ; 
   reg __426645_426645;
   reg _426646_426646 ; 
   reg __426646_426646;
   reg _426647_426647 ; 
   reg __426647_426647;
   reg _426648_426648 ; 
   reg __426648_426648;
   reg _426649_426649 ; 
   reg __426649_426649;
   reg _426650_426650 ; 
   reg __426650_426650;
   reg _426651_426651 ; 
   reg __426651_426651;
   reg _426652_426652 ; 
   reg __426652_426652;
   reg _426653_426653 ; 
   reg __426653_426653;
   reg _426654_426654 ; 
   reg __426654_426654;
   reg _426655_426655 ; 
   reg __426655_426655;
   reg _426656_426656 ; 
   reg __426656_426656;
   reg _426657_426657 ; 
   reg __426657_426657;
   reg _426658_426658 ; 
   reg __426658_426658;
   reg _426659_426659 ; 
   reg __426659_426659;
   reg _426660_426660 ; 
   reg __426660_426660;
   reg _426661_426661 ; 
   reg __426661_426661;
   reg _426662_426662 ; 
   reg __426662_426662;
   reg _426663_426663 ; 
   reg __426663_426663;
   reg _426664_426664 ; 
   reg __426664_426664;
   reg _426665_426665 ; 
   reg __426665_426665;
   reg _426666_426666 ; 
   reg __426666_426666;
   reg _426667_426667 ; 
   reg __426667_426667;
   reg _426668_426668 ; 
   reg __426668_426668;
   reg _426669_426669 ; 
   reg __426669_426669;
   reg _426670_426670 ; 
   reg __426670_426670;
   reg _426671_426671 ; 
   reg __426671_426671;
   reg _426672_426672 ; 
   reg __426672_426672;
   reg _426673_426673 ; 
   reg __426673_426673;
   reg _426674_426674 ; 
   reg __426674_426674;
   reg _426675_426675 ; 
   reg __426675_426675;
   reg _426676_426676 ; 
   reg __426676_426676;
   reg _426677_426677 ; 
   reg __426677_426677;
   reg _426678_426678 ; 
   reg __426678_426678;
   reg _426679_426679 ; 
   reg __426679_426679;
   reg _426680_426680 ; 
   reg __426680_426680;
   reg _426681_426681 ; 
   reg __426681_426681;
   reg _426682_426682 ; 
   reg __426682_426682;
   reg _426683_426683 ; 
   reg __426683_426683;
   reg _426684_426684 ; 
   reg __426684_426684;
   reg _426685_426685 ; 
   reg __426685_426685;
   reg _426686_426686 ; 
   reg __426686_426686;
   reg _426687_426687 ; 
   reg __426687_426687;
   reg _426688_426688 ; 
   reg __426688_426688;
   reg _426689_426689 ; 
   reg __426689_426689;
   reg _426690_426690 ; 
   reg __426690_426690;
   reg _426691_426691 ; 
   reg __426691_426691;
   reg _426692_426692 ; 
   reg __426692_426692;
   reg _426693_426693 ; 
   reg __426693_426693;
   reg _426694_426694 ; 
   reg __426694_426694;
   reg _426695_426695 ; 
   reg __426695_426695;
   reg _426696_426696 ; 
   reg __426696_426696;
   reg _426697_426697 ; 
   reg __426697_426697;
   reg _426698_426698 ; 
   reg __426698_426698;
   reg _426699_426699 ; 
   reg __426699_426699;
   reg _426700_426700 ; 
   reg __426700_426700;
   reg _426701_426701 ; 
   reg __426701_426701;
   reg _426702_426702 ; 
   reg __426702_426702;
   reg _426703_426703 ; 
   reg __426703_426703;
   reg _426704_426704 ; 
   reg __426704_426704;
   reg _426705_426705 ; 
   reg __426705_426705;
   reg _426706_426706 ; 
   reg __426706_426706;
   reg _426707_426707 ; 
   reg __426707_426707;
   reg _426708_426708 ; 
   reg __426708_426708;
   reg _426709_426709 ; 
   reg __426709_426709;
   reg _426710_426710 ; 
   reg __426710_426710;
   reg _426711_426711 ; 
   reg __426711_426711;
   reg _426712_426712 ; 
   reg __426712_426712;
   reg _426713_426713 ; 
   reg __426713_426713;
   reg _426714_426714 ; 
   reg __426714_426714;
   reg _426715_426715 ; 
   reg __426715_426715;
   reg _426716_426716 ; 
   reg __426716_426716;
   reg _426717_426717 ; 
   reg __426717_426717;
   reg _426718_426718 ; 
   reg __426718_426718;
   reg _426719_426719 ; 
   reg __426719_426719;
   reg _426720_426720 ; 
   reg __426720_426720;
   reg _426721_426721 ; 
   reg __426721_426721;
   reg _426722_426722 ; 
   reg __426722_426722;
   reg _426723_426723 ; 
   reg __426723_426723;
   reg _426724_426724 ; 
   reg __426724_426724;
   reg _426725_426725 ; 
   reg __426725_426725;
   reg _426726_426726 ; 
   reg __426726_426726;
   reg _426727_426727 ; 
   reg __426727_426727;
   reg _426728_426728 ; 
   reg __426728_426728;
   reg _426729_426729 ; 
   reg __426729_426729;
   reg _426730_426730 ; 
   reg __426730_426730;
   reg _426731_426731 ; 
   reg __426731_426731;
   reg _426732_426732 ; 
   reg __426732_426732;
   reg _426733_426733 ; 
   reg __426733_426733;
   reg _426734_426734 ; 
   reg __426734_426734;
   reg _426735_426735 ; 
   reg __426735_426735;
   reg _426736_426736 ; 
   reg __426736_426736;
   reg _426737_426737 ; 
   reg __426737_426737;
   reg _426738_426738 ; 
   reg __426738_426738;
   reg _426739_426739 ; 
   reg __426739_426739;
   reg _426740_426740 ; 
   reg __426740_426740;
   reg _426741_426741 ; 
   reg __426741_426741;
   reg _426742_426742 ; 
   reg __426742_426742;
   reg _426743_426743 ; 
   reg __426743_426743;
   reg _426744_426744 ; 
   reg __426744_426744;
   reg _426745_426745 ; 
   reg __426745_426745;
   reg _426746_426746 ; 
   reg __426746_426746;
   reg _426747_426747 ; 
   reg __426747_426747;
   reg _426748_426748 ; 
   reg __426748_426748;
   reg _426749_426749 ; 
   reg __426749_426749;
   reg _426750_426750 ; 
   reg __426750_426750;
   reg _426751_426751 ; 
   reg __426751_426751;
   reg _426752_426752 ; 
   reg __426752_426752;
   reg _426753_426753 ; 
   reg __426753_426753;
   reg _426754_426754 ; 
   reg __426754_426754;
   reg _426755_426755 ; 
   reg __426755_426755;
   reg _426756_426756 ; 
   reg __426756_426756;
   reg _426757_426757 ; 
   reg __426757_426757;
   reg _426758_426758 ; 
   reg __426758_426758;
   reg _426759_426759 ; 
   reg __426759_426759;
   reg _426760_426760 ; 
   reg __426760_426760;
   reg _426761_426761 ; 
   reg __426761_426761;
   reg _426762_426762 ; 
   reg __426762_426762;
   reg _426763_426763 ; 
   reg __426763_426763;
   reg _426764_426764 ; 
   reg __426764_426764;
   reg _426765_426765 ; 
   reg __426765_426765;
   reg _426766_426766 ; 
   reg __426766_426766;
   reg _426767_426767 ; 
   reg __426767_426767;
   reg _426768_426768 ; 
   reg __426768_426768;
   reg _426769_426769 ; 
   reg __426769_426769;
   reg _426770_426770 ; 
   reg __426770_426770;
   reg _426771_426771 ; 
   reg __426771_426771;
   reg _426772_426772 ; 
   reg __426772_426772;
   reg _426773_426773 ; 
   reg __426773_426773;
   reg _426774_426774 ; 
   reg __426774_426774;
   reg _426775_426775 ; 
   reg __426775_426775;
   reg _426776_426776 ; 
   reg __426776_426776;
   reg _426777_426777 ; 
   reg __426777_426777;
   reg _426778_426778 ; 
   reg __426778_426778;
   reg _426779_426779 ; 
   reg __426779_426779;
   reg _426780_426780 ; 
   reg __426780_426780;
   reg _426781_426781 ; 
   reg __426781_426781;
   reg _426782_426782 ; 
   reg __426782_426782;
   reg _426783_426783 ; 
   reg __426783_426783;
   reg _426784_426784 ; 
   reg __426784_426784;
   reg _426785_426785 ; 
   reg __426785_426785;
   reg _426786_426786 ; 
   reg __426786_426786;
   reg _426787_426787 ; 
   reg __426787_426787;
   reg _426788_426788 ; 
   reg __426788_426788;
   reg _426789_426789 ; 
   reg __426789_426789;
   reg _426790_426790 ; 
   reg __426790_426790;
   reg _426791_426791 ; 
   reg __426791_426791;
   reg _426792_426792 ; 
   reg __426792_426792;
   reg _426793_426793 ; 
   reg __426793_426793;
   reg _426794_426794 ; 
   reg __426794_426794;
   reg _426795_426795 ; 
   reg __426795_426795;
   reg _426796_426796 ; 
   reg __426796_426796;
   reg _426797_426797 ; 
   reg __426797_426797;
   reg _426798_426798 ; 
   reg __426798_426798;
   reg _426799_426799 ; 
   reg __426799_426799;
   reg _426800_426800 ; 
   reg __426800_426800;
   reg _426801_426801 ; 
   reg __426801_426801;
   reg _426802_426802 ; 
   reg __426802_426802;
   reg _426803_426803 ; 
   reg __426803_426803;
   reg _426804_426804 ; 
   reg __426804_426804;
   reg _426805_426805 ; 
   reg __426805_426805;
   reg _426806_426806 ; 
   reg __426806_426806;
   reg _426807_426807 ; 
   reg __426807_426807;
   reg _426808_426808 ; 
   reg __426808_426808;
   reg _426809_426809 ; 
   reg __426809_426809;
   reg _426810_426810 ; 
   reg __426810_426810;
   reg _426811_426811 ; 
   reg __426811_426811;
   reg _426812_426812 ; 
   reg __426812_426812;
   reg _426813_426813 ; 
   reg __426813_426813;
   reg _426814_426814 ; 
   reg __426814_426814;
   reg _426815_426815 ; 
   reg __426815_426815;
   reg _426816_426816 ; 
   reg __426816_426816;
   reg _426817_426817 ; 
   reg __426817_426817;
   reg _426818_426818 ; 
   reg __426818_426818;
   reg _426819_426819 ; 
   reg __426819_426819;
   reg _426820_426820 ; 
   reg __426820_426820;
   reg _426821_426821 ; 
   reg __426821_426821;
   reg _426822_426822 ; 
   reg __426822_426822;
   reg _426823_426823 ; 
   reg __426823_426823;
   reg _426824_426824 ; 
   reg __426824_426824;
   reg _426825_426825 ; 
   reg __426825_426825;
   reg _426826_426826 ; 
   reg __426826_426826;
   reg _426827_426827 ; 
   reg __426827_426827;
   reg _426828_426828 ; 
   reg __426828_426828;
   reg _426829_426829 ; 
   reg __426829_426829;
   reg _426830_426830 ; 
   reg __426830_426830;
   reg _426831_426831 ; 
   reg __426831_426831;
   reg _426832_426832 ; 
   reg __426832_426832;
   reg _426833_426833 ; 
   reg __426833_426833;
   reg _426834_426834 ; 
   reg __426834_426834;
   reg _426835_426835 ; 
   reg __426835_426835;
   reg _426836_426836 ; 
   reg __426836_426836;
   reg _426837_426837 ; 
   reg __426837_426837;
   reg _426838_426838 ; 
   reg __426838_426838;
   reg _426839_426839 ; 
   reg __426839_426839;
   reg _426840_426840 ; 
   reg __426840_426840;
   reg _426841_426841 ; 
   reg __426841_426841;
   reg _426842_426842 ; 
   reg __426842_426842;
   reg _426843_426843 ; 
   reg __426843_426843;
   reg _426844_426844 ; 
   reg __426844_426844;
   reg _426845_426845 ; 
   reg __426845_426845;
   reg _426846_426846 ; 
   reg __426846_426846;
   reg _426847_426847 ; 
   reg __426847_426847;
   reg _426848_426848 ; 
   reg __426848_426848;
   reg _426849_426849 ; 
   reg __426849_426849;
   reg _426850_426850 ; 
   reg __426850_426850;
   reg _426851_426851 ; 
   reg __426851_426851;
   reg _426852_426852 ; 
   reg __426852_426852;
   reg _426853_426853 ; 
   reg __426853_426853;
   reg _426854_426854 ; 
   reg __426854_426854;
   reg _426855_426855 ; 
   reg __426855_426855;
   reg _426856_426856 ; 
   reg __426856_426856;
   reg _426857_426857 ; 
   reg __426857_426857;
   reg _426858_426858 ; 
   reg __426858_426858;
   reg _426859_426859 ; 
   reg __426859_426859;
   reg _426860_426860 ; 
   reg __426860_426860;
   reg _426861_426861 ; 
   reg __426861_426861;
   reg _426862_426862 ; 
   reg __426862_426862;
   reg _426863_426863 ; 
   reg __426863_426863;
   reg _426864_426864 ; 
   reg __426864_426864;
   reg _426865_426865 ; 
   reg __426865_426865;
   reg _426866_426866 ; 
   reg __426866_426866;
   reg _426867_426867 ; 
   reg __426867_426867;
   reg _426868_426868 ; 
   reg __426868_426868;
   reg _426869_426869 ; 
   reg __426869_426869;
   reg _426870_426870 ; 
   reg __426870_426870;
   reg _426871_426871 ; 
   reg __426871_426871;
   reg _426872_426872 ; 
   reg __426872_426872;
   reg _426873_426873 ; 
   reg __426873_426873;
   reg _426874_426874 ; 
   reg __426874_426874;
   reg _426875_426875 ; 
   reg __426875_426875;
   reg _426876_426876 ; 
   reg __426876_426876;
   reg _426877_426877 ; 
   reg __426877_426877;
   reg _426878_426878 ; 
   reg __426878_426878;
   reg _426879_426879 ; 
   reg __426879_426879;
   reg _426880_426880 ; 
   reg __426880_426880;
   reg _426881_426881 ; 
   reg __426881_426881;
   reg _426882_426882 ; 
   reg __426882_426882;
   reg _426883_426883 ; 
   reg __426883_426883;
   reg _426884_426884 ; 
   reg __426884_426884;
   reg _426885_426885 ; 
   reg __426885_426885;
   reg _426886_426886 ; 
   reg __426886_426886;
   reg _426887_426887 ; 
   reg __426887_426887;
   reg _426888_426888 ; 
   reg __426888_426888;
   reg _426889_426889 ; 
   reg __426889_426889;
   reg _426890_426890 ; 
   reg __426890_426890;
   reg _426891_426891 ; 
   reg __426891_426891;
   reg _426892_426892 ; 
   reg __426892_426892;
   reg _426893_426893 ; 
   reg __426893_426893;
   reg _426894_426894 ; 
   reg __426894_426894;
   reg _426895_426895 ; 
   reg __426895_426895;
   reg _426896_426896 ; 
   reg __426896_426896;
   reg _426897_426897 ; 
   reg __426897_426897;
   reg _426898_426898 ; 
   reg __426898_426898;
   reg _426899_426899 ; 
   reg __426899_426899;
   reg _426900_426900 ; 
   reg __426900_426900;
   reg _426901_426901 ; 
   reg __426901_426901;
   reg _426902_426902 ; 
   reg __426902_426902;
   reg _426903_426903 ; 
   reg __426903_426903;
   reg _426904_426904 ; 
   reg __426904_426904;
   reg _426905_426905 ; 
   reg __426905_426905;
   reg _426906_426906 ; 
   reg __426906_426906;
   reg _426907_426907 ; 
   reg __426907_426907;
   reg _426908_426908 ; 
   reg __426908_426908;
   reg _426909_426909 ; 
   reg __426909_426909;
   reg _426910_426910 ; 
   reg __426910_426910;
   reg _426911_426911 ; 
   reg __426911_426911;
   reg _426912_426912 ; 
   reg __426912_426912;
   reg _426913_426913 ; 
   reg __426913_426913;
   reg _426914_426914 ; 
   reg __426914_426914;
   reg _426915_426915 ; 
   reg __426915_426915;
   reg _426916_426916 ; 
   reg __426916_426916;
   reg _426917_426917 ; 
   reg __426917_426917;
   reg _426918_426918 ; 
   reg __426918_426918;
   reg _426919_426919 ; 
   reg __426919_426919;
   reg _426920_426920 ; 
   reg __426920_426920;
   reg _426921_426921 ; 
   reg __426921_426921;
   reg _426922_426922 ; 
   reg __426922_426922;
   reg _426923_426923 ; 
   reg __426923_426923;
   reg _426924_426924 ; 
   reg __426924_426924;
   reg _426925_426925 ; 
   reg __426925_426925;
   reg _426926_426926 ; 
   reg __426926_426926;
   reg _426927_426927 ; 
   reg __426927_426927;
   reg _426928_426928 ; 
   reg __426928_426928;
   reg _426929_426929 ; 
   reg __426929_426929;
   reg _426930_426930 ; 
   reg __426930_426930;
   reg _426931_426931 ; 
   reg __426931_426931;
   reg _426932_426932 ; 
   reg __426932_426932;
   reg _426933_426933 ; 
   reg __426933_426933;
   reg _426934_426934 ; 
   reg __426934_426934;
   reg _426935_426935 ; 
   reg __426935_426935;
   reg _426936_426936 ; 
   reg __426936_426936;
   reg _426937_426937 ; 
   reg __426937_426937;
   reg _426938_426938 ; 
   reg __426938_426938;
   reg _426939_426939 ; 
   reg __426939_426939;
   reg _426940_426940 ; 
   reg __426940_426940;
   reg _426941_426941 ; 
   reg __426941_426941;
   reg _426942_426942 ; 
   reg __426942_426942;
   reg _426943_426943 ; 
   reg __426943_426943;
   reg _426944_426944 ; 
   reg __426944_426944;
   reg _426945_426945 ; 
   reg __426945_426945;
   reg _426946_426946 ; 
   reg __426946_426946;
   reg _426947_426947 ; 
   reg __426947_426947;
   reg _426948_426948 ; 
   reg __426948_426948;
   reg _426949_426949 ; 
   reg __426949_426949;
   reg _426950_426950 ; 
   reg __426950_426950;
   reg _426951_426951 ; 
   reg __426951_426951;
   reg _426952_426952 ; 
   reg __426952_426952;
   reg _426953_426953 ; 
   reg __426953_426953;
   reg _426954_426954 ; 
   reg __426954_426954;
   reg _426955_426955 ; 
   reg __426955_426955;
   reg _426956_426956 ; 
   reg __426956_426956;
   reg _426957_426957 ; 
   reg __426957_426957;
   reg _426958_426958 ; 
   reg __426958_426958;
   reg _426959_426959 ; 
   reg __426959_426959;
   reg _426960_426960 ; 
   reg __426960_426960;
   reg _426961_426961 ; 
   reg __426961_426961;
   reg _426962_426962 ; 
   reg __426962_426962;
   reg _426963_426963 ; 
   reg __426963_426963;
   reg _426964_426964 ; 
   reg __426964_426964;
   reg _426965_426965 ; 
   reg __426965_426965;
   reg _426966_426966 ; 
   reg __426966_426966;
   reg _426967_426967 ; 
   reg __426967_426967;
   reg _426968_426968 ; 
   reg __426968_426968;
   reg _426969_426969 ; 
   reg __426969_426969;
   reg _426970_426970 ; 
   reg __426970_426970;
   reg _426971_426971 ; 
   reg __426971_426971;
   reg _426972_426972 ; 
   reg __426972_426972;
   reg _426973_426973 ; 
   reg __426973_426973;
   reg _426974_426974 ; 
   reg __426974_426974;
   reg _426975_426975 ; 
   reg __426975_426975;
   reg _426976_426976 ; 
   reg __426976_426976;
   reg _426977_426977 ; 
   reg __426977_426977;
   reg _426978_426978 ; 
   reg __426978_426978;
   reg _426979_426979 ; 
   reg __426979_426979;
   reg _426980_426980 ; 
   reg __426980_426980;
   reg _426981_426981 ; 
   reg __426981_426981;
   reg _426982_426982 ; 
   reg __426982_426982;
   reg _426983_426983 ; 
   reg __426983_426983;
   reg _426984_426984 ; 
   reg __426984_426984;
   reg _426985_426985 ; 
   reg __426985_426985;
   reg _426986_426986 ; 
   reg __426986_426986;
   reg _426987_426987 ; 
   reg __426987_426987;
   reg _426988_426988 ; 
   reg __426988_426988;
   reg _426989_426989 ; 
   reg __426989_426989;
   reg _426990_426990 ; 
   reg __426990_426990;
   reg _426991_426991 ; 
   reg __426991_426991;
   reg _426992_426992 ; 
   reg __426992_426992;
   reg _426993_426993 ; 
   reg __426993_426993;
   reg _426994_426994 ; 
   reg __426994_426994;
   reg _426995_426995 ; 
   reg __426995_426995;
   reg _426996_426996 ; 
   reg __426996_426996;
   reg _426997_426997 ; 
   reg __426997_426997;
   reg _426998_426998 ; 
   reg __426998_426998;
   reg _426999_426999 ; 
   reg __426999_426999;
   reg _427000_427000 ; 
   reg __427000_427000;
   reg _427001_427001 ; 
   reg __427001_427001;
   reg _427002_427002 ; 
   reg __427002_427002;
   reg _427003_427003 ; 
   reg __427003_427003;
   reg _427004_427004 ; 
   reg __427004_427004;
   reg _427005_427005 ; 
   reg __427005_427005;
   reg _427006_427006 ; 
   reg __427006_427006;
   reg _427007_427007 ; 
   reg __427007_427007;
   reg _427008_427008 ; 
   reg __427008_427008;
   reg _427009_427009 ; 
   reg __427009_427009;
   reg _427010_427010 ; 
   reg __427010_427010;
   reg _427011_427011 ; 
   reg __427011_427011;
   reg _427012_427012 ; 
   reg __427012_427012;
   reg _427013_427013 ; 
   reg __427013_427013;
   reg _427014_427014 ; 
   reg __427014_427014;
   reg _427015_427015 ; 
   reg __427015_427015;
   reg _427016_427016 ; 
   reg __427016_427016;
   reg _427017_427017 ; 
   reg __427017_427017;
   reg _427018_427018 ; 
   reg __427018_427018;
   reg _427019_427019 ; 
   reg __427019_427019;
   reg _427020_427020 ; 
   reg __427020_427020;
   reg _427021_427021 ; 
   reg __427021_427021;
   reg _427022_427022 ; 
   reg __427022_427022;
   reg _427023_427023 ; 
   reg __427023_427023;
   reg _427024_427024 ; 
   reg __427024_427024;
   reg _427025_427025 ; 
   reg __427025_427025;
   reg _427026_427026 ; 
   reg __427026_427026;
   reg _427027_427027 ; 
   reg __427027_427027;
   reg _427028_427028 ; 
   reg __427028_427028;
   reg _427029_427029 ; 
   reg __427029_427029;
   reg _427030_427030 ; 
   reg __427030_427030;
   reg _427031_427031 ; 
   reg __427031_427031;
   reg _427032_427032 ; 
   reg __427032_427032;
   reg _427033_427033 ; 
   reg __427033_427033;
   reg _427034_427034 ; 
   reg __427034_427034;
   reg _427035_427035 ; 
   reg __427035_427035;
   reg _427036_427036 ; 
   reg __427036_427036;
   reg _427037_427037 ; 
   reg __427037_427037;
   reg _427038_427038 ; 
   reg __427038_427038;
   reg _427039_427039 ; 
   reg __427039_427039;
   reg _427040_427040 ; 
   reg __427040_427040;
   reg _427041_427041 ; 
   reg __427041_427041;
   reg _427042_427042 ; 
   reg __427042_427042;
   reg _427043_427043 ; 
   reg __427043_427043;
   reg _427044_427044 ; 
   reg __427044_427044;
   reg _427045_427045 ; 
   reg __427045_427045;
   reg _427046_427046 ; 
   reg __427046_427046;
   reg _427047_427047 ; 
   reg __427047_427047;
   reg _427048_427048 ; 
   reg __427048_427048;
   reg _427049_427049 ; 
   reg __427049_427049;
   reg _427050_427050 ; 
   reg __427050_427050;
   reg _427051_427051 ; 
   reg __427051_427051;
   reg _427052_427052 ; 
   reg __427052_427052;
   reg _427053_427053 ; 
   reg __427053_427053;
   reg _427054_427054 ; 
   reg __427054_427054;
   reg _427055_427055 ; 
   reg __427055_427055;
   reg _427056_427056 ; 
   reg __427056_427056;
   reg _427057_427057 ; 
   reg __427057_427057;
   reg _427058_427058 ; 
   reg __427058_427058;
   reg _427059_427059 ; 
   reg __427059_427059;
   reg _427060_427060 ; 
   reg __427060_427060;
   reg _427061_427061 ; 
   reg __427061_427061;
   reg _427062_427062 ; 
   reg __427062_427062;
   reg _427063_427063 ; 
   reg __427063_427063;
   reg _427064_427064 ; 
   reg __427064_427064;
   reg _427065_427065 ; 
   reg __427065_427065;
   reg _427066_427066 ; 
   reg __427066_427066;
   reg _427067_427067 ; 
   reg __427067_427067;
   reg _427068_427068 ; 
   reg __427068_427068;
   reg _427069_427069 ; 
   reg __427069_427069;
   reg _427070_427070 ; 
   reg __427070_427070;
   reg _427071_427071 ; 
   reg __427071_427071;
   reg _427072_427072 ; 
   reg __427072_427072;
   reg _427073_427073 ; 
   reg __427073_427073;
   reg _427074_427074 ; 
   reg __427074_427074;
   reg _427075_427075 ; 
   reg __427075_427075;
   reg _427076_427076 ; 
   reg __427076_427076;
   reg _427077_427077 ; 
   reg __427077_427077;
   reg _427078_427078 ; 
   reg __427078_427078;
   reg _427079_427079 ; 
   reg __427079_427079;
   reg _427080_427080 ; 
   reg __427080_427080;
   reg _427081_427081 ; 
   reg __427081_427081;
   reg _427082_427082 ; 
   reg __427082_427082;
   reg _427083_427083 ; 
   reg __427083_427083;
   reg _427084_427084 ; 
   reg __427084_427084;
   reg _427085_427085 ; 
   reg __427085_427085;
   reg _427086_427086 ; 
   reg __427086_427086;
   reg _427087_427087 ; 
   reg __427087_427087;
   reg _427088_427088 ; 
   reg __427088_427088;
   reg _427089_427089 ; 
   reg __427089_427089;
   reg _427090_427090 ; 
   reg __427090_427090;
   reg _427091_427091 ; 
   reg __427091_427091;
   reg _427092_427092 ; 
   reg __427092_427092;
   reg _427093_427093 ; 
   reg __427093_427093;
   reg _427094_427094 ; 
   reg __427094_427094;
   reg _427095_427095 ; 
   reg __427095_427095;
   reg _427096_427096 ; 
   reg __427096_427096;
   reg _427097_427097 ; 
   reg __427097_427097;
   reg _427098_427098 ; 
   reg __427098_427098;
   reg _427099_427099 ; 
   reg __427099_427099;
   reg _427100_427100 ; 
   reg __427100_427100;
   reg _427101_427101 ; 
   reg __427101_427101;
   reg _427102_427102 ; 
   reg __427102_427102;
   reg _427103_427103 ; 
   reg __427103_427103;
   reg _427104_427104 ; 
   reg __427104_427104;
   reg _427105_427105 ; 
   reg __427105_427105;
   reg _427106_427106 ; 
   reg __427106_427106;
   reg _427107_427107 ; 
   reg __427107_427107;
   reg _427108_427108 ; 
   reg __427108_427108;
   reg _427109_427109 ; 
   reg __427109_427109;
   reg _427110_427110 ; 
   reg __427110_427110;
   reg _427111_427111 ; 
   reg __427111_427111;
   reg _427112_427112 ; 
   reg __427112_427112;
   reg _427113_427113 ; 
   reg __427113_427113;
   reg _427114_427114 ; 
   reg __427114_427114;
   reg _427115_427115 ; 
   reg __427115_427115;
   reg _427116_427116 ; 
   reg __427116_427116;
   reg _427117_427117 ; 
   reg __427117_427117;
   reg _427118_427118 ; 
   reg __427118_427118;
   reg _427119_427119 ; 
   reg __427119_427119;
   reg _427120_427120 ; 
   reg __427120_427120;
   reg _427121_427121 ; 
   reg __427121_427121;
   reg _427122_427122 ; 
   reg __427122_427122;
   reg _427123_427123 ; 
   reg __427123_427123;
   reg _427124_427124 ; 
   reg __427124_427124;
   reg _427125_427125 ; 
   reg __427125_427125;
   reg _427126_427126 ; 
   reg __427126_427126;
   reg _427127_427127 ; 
   reg __427127_427127;
   reg _427128_427128 ; 
   reg __427128_427128;
   reg _427129_427129 ; 
   reg __427129_427129;
   reg _427130_427130 ; 
   reg __427130_427130;
   reg _427131_427131 ; 
   reg __427131_427131;
   reg _427132_427132 ; 
   reg __427132_427132;
   reg _427133_427133 ; 
   reg __427133_427133;
   reg _427134_427134 ; 
   reg __427134_427134;
   reg _427135_427135 ; 
   reg __427135_427135;
   reg _427136_427136 ; 
   reg __427136_427136;
   reg _427137_427137 ; 
   reg __427137_427137;
   reg _427138_427138 ; 
   reg __427138_427138;
   reg _427139_427139 ; 
   reg __427139_427139;
   reg _427140_427140 ; 
   reg __427140_427140;
   reg _427141_427141 ; 
   reg __427141_427141;
   reg _427142_427142 ; 
   reg __427142_427142;
   reg _427143_427143 ; 
   reg __427143_427143;
   reg _427144_427144 ; 
   reg __427144_427144;
   reg _427145_427145 ; 
   reg __427145_427145;
   reg _427146_427146 ; 
   reg __427146_427146;
   reg _427147_427147 ; 
   reg __427147_427147;
   reg _427148_427148 ; 
   reg __427148_427148;
   reg _427149_427149 ; 
   reg __427149_427149;
   reg _427150_427150 ; 
   reg __427150_427150;
   reg _427151_427151 ; 
   reg __427151_427151;
   reg _427152_427152 ; 
   reg __427152_427152;
   reg _427153_427153 ; 
   reg __427153_427153;
   reg _427154_427154 ; 
   reg __427154_427154;
   reg _427155_427155 ; 
   reg __427155_427155;
   reg _427156_427156 ; 
   reg __427156_427156;
   reg _427157_427157 ; 
   reg __427157_427157;
   reg _427158_427158 ; 
   reg __427158_427158;
   reg _427159_427159 ; 
   reg __427159_427159;
   reg _427160_427160 ; 
   reg __427160_427160;
   reg _427161_427161 ; 
   reg __427161_427161;
   reg _427162_427162 ; 
   reg __427162_427162;
   reg _427163_427163 ; 
   reg __427163_427163;
   reg _427164_427164 ; 
   reg __427164_427164;
   reg _427165_427165 ; 
   reg __427165_427165;
   reg _427166_427166 ; 
   reg __427166_427166;
   reg _427167_427167 ; 
   reg __427167_427167;
   reg _427168_427168 ; 
   reg __427168_427168;
   reg _427169_427169 ; 
   reg __427169_427169;
   reg _427170_427170 ; 
   reg __427170_427170;
   reg _427171_427171 ; 
   reg __427171_427171;
   reg _427172_427172 ; 
   reg __427172_427172;
   reg _427173_427173 ; 
   reg __427173_427173;
   reg _427174_427174 ; 
   reg __427174_427174;
   reg _427175_427175 ; 
   reg __427175_427175;
   reg _427176_427176 ; 
   reg __427176_427176;
   reg _427177_427177 ; 
   reg __427177_427177;
   reg _427178_427178 ; 
   reg __427178_427178;
   reg _427179_427179 ; 
   reg __427179_427179;
   reg _427180_427180 ; 
   reg __427180_427180;
   reg _427181_427181 ; 
   reg __427181_427181;
   reg _427182_427182 ; 
   reg __427182_427182;
   reg _427183_427183 ; 
   reg __427183_427183;
   reg _427184_427184 ; 
   reg __427184_427184;
   reg _427185_427185 ; 
   reg __427185_427185;
   reg _427186_427186 ; 
   reg __427186_427186;
   reg _427187_427187 ; 
   reg __427187_427187;
   reg _427188_427188 ; 
   reg __427188_427188;
   reg _427189_427189 ; 
   reg __427189_427189;
   reg _427190_427190 ; 
   reg __427190_427190;
   reg _427191_427191 ; 
   reg __427191_427191;
   reg _427192_427192 ; 
   reg __427192_427192;
   reg _427193_427193 ; 
   reg __427193_427193;
   reg _427194_427194 ; 
   reg __427194_427194;
   reg _427195_427195 ; 
   reg __427195_427195;
   reg _427196_427196 ; 
   reg __427196_427196;
   reg _427197_427197 ; 
   reg __427197_427197;
   reg _427198_427198 ; 
   reg __427198_427198;
   reg _427199_427199 ; 
   reg __427199_427199;
   reg _427200_427200 ; 
   reg __427200_427200;
   reg _427201_427201 ; 
   reg __427201_427201;
   reg _427202_427202 ; 
   reg __427202_427202;
   reg _427203_427203 ; 
   reg __427203_427203;
   reg _427204_427204 ; 
   reg __427204_427204;
   reg _427205_427205 ; 
   reg __427205_427205;
   reg _427206_427206 ; 
   reg __427206_427206;
   reg _427207_427207 ; 
   reg __427207_427207;
   reg _427208_427208 ; 
   reg __427208_427208;
   reg _427209_427209 ; 
   reg __427209_427209;
   reg _427210_427210 ; 
   reg __427210_427210;
   reg _427211_427211 ; 
   reg __427211_427211;
   reg _427212_427212 ; 
   reg __427212_427212;
   reg _427213_427213 ; 
   reg __427213_427213;
   reg _427214_427214 ; 
   reg __427214_427214;
   reg _427215_427215 ; 
   reg __427215_427215;
   reg _427216_427216 ; 
   reg __427216_427216;
   reg _427217_427217 ; 
   reg __427217_427217;
   reg _427218_427218 ; 
   reg __427218_427218;
   reg _427219_427219 ; 
   reg __427219_427219;
   reg _427220_427220 ; 
   reg __427220_427220;
   reg _427221_427221 ; 
   reg __427221_427221;
   reg _427222_427222 ; 
   reg __427222_427222;
   reg _427223_427223 ; 
   reg __427223_427223;
   reg _427224_427224 ; 
   reg __427224_427224;
   reg _427225_427225 ; 
   reg __427225_427225;
   reg _427226_427226 ; 
   reg __427226_427226;
   reg _427227_427227 ; 
   reg __427227_427227;
   reg _427228_427228 ; 
   reg __427228_427228;
   reg _427229_427229 ; 
   reg __427229_427229;
   reg _427230_427230 ; 
   reg __427230_427230;
   reg _427231_427231 ; 
   reg __427231_427231;
   reg _427232_427232 ; 
   reg __427232_427232;
   reg _427233_427233 ; 
   reg __427233_427233;
   reg _427234_427234 ; 
   reg __427234_427234;
   reg _427235_427235 ; 
   reg __427235_427235;
   reg _427236_427236 ; 
   reg __427236_427236;
   reg _427237_427237 ; 
   reg __427237_427237;
   reg _427238_427238 ; 
   reg __427238_427238;
   reg _427239_427239 ; 
   reg __427239_427239;
   reg _427240_427240 ; 
   reg __427240_427240;
   reg _427241_427241 ; 
   reg __427241_427241;
   reg _427242_427242 ; 
   reg __427242_427242;
   reg _427243_427243 ; 
   reg __427243_427243;
   reg _427244_427244 ; 
   reg __427244_427244;
   reg _427245_427245 ; 
   reg __427245_427245;
   reg _427246_427246 ; 
   reg __427246_427246;
   reg _427247_427247 ; 
   reg __427247_427247;
   reg _427248_427248 ; 
   reg __427248_427248;
   reg _427249_427249 ; 
   reg __427249_427249;
   reg _427250_427250 ; 
   reg __427250_427250;
   reg _427251_427251 ; 
   reg __427251_427251;
   reg _427252_427252 ; 
   reg __427252_427252;
   reg _427253_427253 ; 
   reg __427253_427253;
   reg _427254_427254 ; 
   reg __427254_427254;
   reg _427255_427255 ; 
   reg __427255_427255;
   reg _427256_427256 ; 
   reg __427256_427256;
   reg _427257_427257 ; 
   reg __427257_427257;
   reg _427258_427258 ; 
   reg __427258_427258;
   reg _427259_427259 ; 
   reg __427259_427259;
   reg _427260_427260 ; 
   reg __427260_427260;
   reg _427261_427261 ; 
   reg __427261_427261;
   reg _427262_427262 ; 
   reg __427262_427262;
   reg _427263_427263 ; 
   reg __427263_427263;
   reg _427264_427264 ; 
   reg __427264_427264;
   reg _427265_427265 ; 
   reg __427265_427265;
   reg _427266_427266 ; 
   reg __427266_427266;
   reg _427267_427267 ; 
   reg __427267_427267;
   reg _427268_427268 ; 
   reg __427268_427268;
   reg _427269_427269 ; 
   reg __427269_427269;
   reg _427270_427270 ; 
   reg __427270_427270;
   reg _427271_427271 ; 
   reg __427271_427271;
   reg _427272_427272 ; 
   reg __427272_427272;
   reg _427273_427273 ; 
   reg __427273_427273;
   reg _427274_427274 ; 
   reg __427274_427274;
   reg _427275_427275 ; 
   reg __427275_427275;
   reg _427276_427276 ; 
   reg __427276_427276;
   reg _427277_427277 ; 
   reg __427277_427277;
   reg _427278_427278 ; 
   reg __427278_427278;
   reg _427279_427279 ; 
   reg __427279_427279;
   reg _427280_427280 ; 
   reg __427280_427280;
   reg _427281_427281 ; 
   reg __427281_427281;
   reg _427282_427282 ; 
   reg __427282_427282;
   reg _427283_427283 ; 
   reg __427283_427283;
   reg _427284_427284 ; 
   reg __427284_427284;
   reg _427285_427285 ; 
   reg __427285_427285;
   reg _427286_427286 ; 
   reg __427286_427286;
   reg _427287_427287 ; 
   reg __427287_427287;
   reg _427288_427288 ; 
   reg __427288_427288;
   reg _427289_427289 ; 
   reg __427289_427289;
   reg _427290_427290 ; 
   reg __427290_427290;
   reg _427291_427291 ; 
   reg __427291_427291;
   reg _427292_427292 ; 
   reg __427292_427292;
   reg _427293_427293 ; 
   reg __427293_427293;
   reg _427294_427294 ; 
   reg __427294_427294;
   reg _427295_427295 ; 
   reg __427295_427295;
   reg _427296_427296 ; 
   reg __427296_427296;
   reg _427297_427297 ; 
   reg __427297_427297;
   reg _427298_427298 ; 
   reg __427298_427298;
   reg _427299_427299 ; 
   reg __427299_427299;
   reg _427300_427300 ; 
   reg __427300_427300;
   reg _427301_427301 ; 
   reg __427301_427301;
   reg _427302_427302 ; 
   reg __427302_427302;
   reg _427303_427303 ; 
   reg __427303_427303;
   reg _427304_427304 ; 
   reg __427304_427304;
   reg _427305_427305 ; 
   reg __427305_427305;
   reg _427306_427306 ; 
   reg __427306_427306;
   reg _427307_427307 ; 
   reg __427307_427307;
   reg _427308_427308 ; 
   reg __427308_427308;
   reg _427309_427309 ; 
   reg __427309_427309;
   reg _427310_427310 ; 
   reg __427310_427310;
   reg _427311_427311 ; 
   reg __427311_427311;
   reg _427312_427312 ; 
   reg __427312_427312;
   reg _427313_427313 ; 
   reg __427313_427313;
   reg _427314_427314 ; 
   reg __427314_427314;
   reg _427315_427315 ; 
   reg __427315_427315;
   reg _427316_427316 ; 
   reg __427316_427316;
   reg _427317_427317 ; 
   reg __427317_427317;
   reg _427318_427318 ; 
   reg __427318_427318;
   reg _427319_427319 ; 
   reg __427319_427319;
   reg _427320_427320 ; 
   reg __427320_427320;
   reg _427321_427321 ; 
   reg __427321_427321;
   reg _427322_427322 ; 
   reg __427322_427322;
   reg _427323_427323 ; 
   reg __427323_427323;
   reg _427324_427324 ; 
   reg __427324_427324;
   reg _427325_427325 ; 
   reg __427325_427325;
   reg _427326_427326 ; 
   reg __427326_427326;
   reg _427327_427327 ; 
   reg __427327_427327;
   reg _427328_427328 ; 
   reg __427328_427328;
   reg _427329_427329 ; 
   reg __427329_427329;
   reg _427330_427330 ; 
   reg __427330_427330;
   reg _427331_427331 ; 
   reg __427331_427331;
   reg _427332_427332 ; 
   reg __427332_427332;
   reg _427333_427333 ; 
   reg __427333_427333;
   reg _427334_427334 ; 
   reg __427334_427334;
   reg _427335_427335 ; 
   reg __427335_427335;
   reg _427336_427336 ; 
   reg __427336_427336;
   reg _427337_427337 ; 
   reg __427337_427337;
   reg _427338_427338 ; 
   reg __427338_427338;
   reg _427339_427339 ; 
   reg __427339_427339;
   reg _427340_427340 ; 
   reg __427340_427340;
   reg _427341_427341 ; 
   reg __427341_427341;
   reg _427342_427342 ; 
   reg __427342_427342;
   reg _427343_427343 ; 
   reg __427343_427343;
   reg _427344_427344 ; 
   reg __427344_427344;
   reg _427345_427345 ; 
   reg __427345_427345;
   reg _427346_427346 ; 
   reg __427346_427346;
   reg _427347_427347 ; 
   reg __427347_427347;
   reg _427348_427348 ; 
   reg __427348_427348;
   reg _427349_427349 ; 
   reg __427349_427349;
   reg _427350_427350 ; 
   reg __427350_427350;
   reg _427351_427351 ; 
   reg __427351_427351;
   reg _427352_427352 ; 
   reg __427352_427352;
   reg _427353_427353 ; 
   reg __427353_427353;
   reg _427354_427354 ; 
   reg __427354_427354;
   reg _427355_427355 ; 
   reg __427355_427355;
   reg _427356_427356 ; 
   reg __427356_427356;
   reg _427357_427357 ; 
   reg __427357_427357;
   reg _427358_427358 ; 
   reg __427358_427358;
   reg _427359_427359 ; 
   reg __427359_427359;
   reg _427360_427360 ; 
   reg __427360_427360;
   reg _427361_427361 ; 
   reg __427361_427361;
   reg _427362_427362 ; 
   reg __427362_427362;
   reg _427363_427363 ; 
   reg __427363_427363;
   reg _427364_427364 ; 
   reg __427364_427364;
   reg _427365_427365 ; 
   reg __427365_427365;
   reg _427366_427366 ; 
   reg __427366_427366;
   reg _427367_427367 ; 
   reg __427367_427367;
   reg _427368_427368 ; 
   reg __427368_427368;
   reg _427369_427369 ; 
   reg __427369_427369;
   reg _427370_427370 ; 
   reg __427370_427370;
   reg _427371_427371 ; 
   reg __427371_427371;
   reg _427372_427372 ; 
   reg __427372_427372;
   reg _427373_427373 ; 
   reg __427373_427373;
   reg _427374_427374 ; 
   reg __427374_427374;
   reg _427375_427375 ; 
   reg __427375_427375;
   reg _427376_427376 ; 
   reg __427376_427376;
   reg _427377_427377 ; 
   reg __427377_427377;
   reg _427378_427378 ; 
   reg __427378_427378;
   reg _427379_427379 ; 
   reg __427379_427379;
   reg _427380_427380 ; 
   reg __427380_427380;
   reg _427381_427381 ; 
   reg __427381_427381;
   reg _427382_427382 ; 
   reg __427382_427382;
   reg _427383_427383 ; 
   reg __427383_427383;
   reg _427384_427384 ; 
   reg __427384_427384;
   reg _427385_427385 ; 
   reg __427385_427385;
   reg _427386_427386 ; 
   reg __427386_427386;
   reg _427387_427387 ; 
   reg __427387_427387;
   reg _427388_427388 ; 
   reg __427388_427388;
   reg _427389_427389 ; 
   reg __427389_427389;
   reg _427390_427390 ; 
   reg __427390_427390;
   reg _427391_427391 ; 
   reg __427391_427391;
   reg _427392_427392 ; 
   reg __427392_427392;
   reg _427393_427393 ; 
   reg __427393_427393;
   reg _427394_427394 ; 
   reg __427394_427394;
   reg _427395_427395 ; 
   reg __427395_427395;
   reg _427396_427396 ; 
   reg __427396_427396;
   reg _427397_427397 ; 
   reg __427397_427397;
   reg _427398_427398 ; 
   reg __427398_427398;
   reg _427399_427399 ; 
   reg __427399_427399;
   reg _427400_427400 ; 
   reg __427400_427400;
   reg _427401_427401 ; 
   reg __427401_427401;
   reg _427402_427402 ; 
   reg __427402_427402;
   reg _427403_427403 ; 
   reg __427403_427403;
   reg _427404_427404 ; 
   reg __427404_427404;
   reg _427405_427405 ; 
   reg __427405_427405;
   reg _427406_427406 ; 
   reg __427406_427406;
   reg _427407_427407 ; 
   reg __427407_427407;
   reg _427408_427408 ; 
   reg __427408_427408;
   reg _427409_427409 ; 
   reg __427409_427409;
   reg _427410_427410 ; 
   reg __427410_427410;
   reg _427411_427411 ; 
   reg __427411_427411;
   reg _427412_427412 ; 
   reg __427412_427412;
   reg _427413_427413 ; 
   reg __427413_427413;
   reg _427414_427414 ; 
   reg __427414_427414;
   reg _427415_427415 ; 
   reg __427415_427415;
   reg _427416_427416 ; 
   reg __427416_427416;
   reg _427417_427417 ; 
   reg __427417_427417;
   reg _427418_427418 ; 
   reg __427418_427418;
   reg _427419_427419 ; 
   reg __427419_427419;
   reg _427420_427420 ; 
   reg __427420_427420;
   reg _427421_427421 ; 
   reg __427421_427421;
   reg _427422_427422 ; 
   reg __427422_427422;
   reg _427423_427423 ; 
   reg __427423_427423;
   reg _427424_427424 ; 
   reg __427424_427424;
   reg _427425_427425 ; 
   reg __427425_427425;
   reg _427426_427426 ; 
   reg __427426_427426;
   reg _427427_427427 ; 
   reg __427427_427427;
   reg _427428_427428 ; 
   reg __427428_427428;
   reg _427429_427429 ; 
   reg __427429_427429;
   reg _427430_427430 ; 
   reg __427430_427430;
   reg _427431_427431 ; 
   reg __427431_427431;
   reg _427432_427432 ; 
   reg __427432_427432;
   reg _427433_427433 ; 
   reg __427433_427433;
   reg _427434_427434 ; 
   reg __427434_427434;
   reg _427435_427435 ; 
   reg __427435_427435;
   reg _427436_427436 ; 
   reg __427436_427436;
   reg _427437_427437 ; 
   reg __427437_427437;
   reg _427438_427438 ; 
   reg __427438_427438;
   reg _427439_427439 ; 
   reg __427439_427439;
   reg _427440_427440 ; 
   reg __427440_427440;
   reg _427441_427441 ; 
   reg __427441_427441;
   reg _427442_427442 ; 
   reg __427442_427442;
   reg _427443_427443 ; 
   reg __427443_427443;
   reg _427444_427444 ; 
   reg __427444_427444;
   reg _427445_427445 ; 
   reg __427445_427445;
   reg _427446_427446 ; 
   reg __427446_427446;
   reg _427447_427447 ; 
   reg __427447_427447;
   reg _427448_427448 ; 
   reg __427448_427448;
   reg _427449_427449 ; 
   reg __427449_427449;
   reg _427450_427450 ; 
   reg __427450_427450;
   reg _427451_427451 ; 
   reg __427451_427451;
   reg _427452_427452 ; 
   reg __427452_427452;
   reg _427453_427453 ; 
   reg __427453_427453;
   reg _427454_427454 ; 
   reg __427454_427454;
   reg _427455_427455 ; 
   reg __427455_427455;
   reg _427456_427456 ; 
   reg __427456_427456;
   reg _427457_427457 ; 
   reg __427457_427457;
   reg _427458_427458 ; 
   reg __427458_427458;
   reg _427459_427459 ; 
   reg __427459_427459;
   reg _427460_427460 ; 
   reg __427460_427460;
   reg _427461_427461 ; 
   reg __427461_427461;
   reg _427462_427462 ; 
   reg __427462_427462;
   reg _427463_427463 ; 
   reg __427463_427463;
   reg _427464_427464 ; 
   reg __427464_427464;
   reg _427465_427465 ; 
   reg __427465_427465;
   reg _427466_427466 ; 
   reg __427466_427466;
   reg _427467_427467 ; 
   reg __427467_427467;
   reg _427468_427468 ; 
   reg __427468_427468;
   reg _427469_427469 ; 
   reg __427469_427469;
   reg _427470_427470 ; 
   reg __427470_427470;
   reg _427471_427471 ; 
   reg __427471_427471;
   reg _427472_427472 ; 
   reg __427472_427472;
   reg _427473_427473 ; 
   reg __427473_427473;
   reg _427474_427474 ; 
   reg __427474_427474;
   reg _427475_427475 ; 
   reg __427475_427475;
   reg _427476_427476 ; 
   reg __427476_427476;
   reg _427477_427477 ; 
   reg __427477_427477;
   reg _427478_427478 ; 
   reg __427478_427478;
   reg _427479_427479 ; 
   reg __427479_427479;
   reg _427480_427480 ; 
   reg __427480_427480;
   reg _427481_427481 ; 
   reg __427481_427481;
   reg _427482_427482 ; 
   reg __427482_427482;
   reg _427483_427483 ; 
   reg __427483_427483;
   reg _427484_427484 ; 
   reg __427484_427484;
   reg _427485_427485 ; 
   reg __427485_427485;
   reg _427486_427486 ; 
   reg __427486_427486;
   reg _427487_427487 ; 
   reg __427487_427487;
   reg _427488_427488 ; 
   reg __427488_427488;
   reg _427489_427489 ; 
   reg __427489_427489;
   reg _427490_427490 ; 
   reg __427490_427490;
   reg _427491_427491 ; 
   reg __427491_427491;
   reg _427492_427492 ; 
   reg __427492_427492;
   reg _427493_427493 ; 
   reg __427493_427493;
   reg _427494_427494 ; 
   reg __427494_427494;
   reg _427495_427495 ; 
   reg __427495_427495;
   reg _427496_427496 ; 
   reg __427496_427496;
   reg _427497_427497 ; 
   reg __427497_427497;
   reg _427498_427498 ; 
   reg __427498_427498;
   reg _427499_427499 ; 
   reg __427499_427499;
   reg _427500_427500 ; 
   reg __427500_427500;
   reg _427501_427501 ; 
   reg __427501_427501;
   reg _427502_427502 ; 
   reg __427502_427502;
   reg _427503_427503 ; 
   reg __427503_427503;
   reg _427504_427504 ; 
   reg __427504_427504;
   reg _427505_427505 ; 
   reg __427505_427505;
   reg _427506_427506 ; 
   reg __427506_427506;
   reg _427507_427507 ; 
   reg __427507_427507;
   reg _427508_427508 ; 
   reg __427508_427508;
   reg _427509_427509 ; 
   reg __427509_427509;
   reg _427510_427510 ; 
   reg __427510_427510;
   reg _427511_427511 ; 
   reg __427511_427511;
   reg _427512_427512 ; 
   reg __427512_427512;
   reg _427513_427513 ; 
   reg __427513_427513;
   reg _427514_427514 ; 
   reg __427514_427514;
   reg _427515_427515 ; 
   reg __427515_427515;
   reg _427516_427516 ; 
   reg __427516_427516;
   reg _427517_427517 ; 
   reg __427517_427517;
   reg _427518_427518 ; 
   reg __427518_427518;
   reg _427519_427519 ; 
   reg __427519_427519;
   reg _427520_427520 ; 
   reg __427520_427520;
   reg _427521_427521 ; 
   reg __427521_427521;
   reg _427522_427522 ; 
   reg __427522_427522;
   reg _427523_427523 ; 
   reg __427523_427523;
   reg _427524_427524 ; 
   reg __427524_427524;
   reg _427525_427525 ; 
   reg __427525_427525;
   reg _427526_427526 ; 
   reg __427526_427526;
   reg _427527_427527 ; 
   reg __427527_427527;
   reg _427528_427528 ; 
   reg __427528_427528;
   reg _427529_427529 ; 
   reg __427529_427529;
   reg _427530_427530 ; 
   reg __427530_427530;
   reg _427531_427531 ; 
   reg __427531_427531;
   reg _427532_427532 ; 
   reg __427532_427532;
   reg _427533_427533 ; 
   reg __427533_427533;
   reg _427534_427534 ; 
   reg __427534_427534;
   reg _427535_427535 ; 
   reg __427535_427535;
   reg _427536_427536 ; 
   reg __427536_427536;
   reg _427537_427537 ; 
   reg __427537_427537;
   reg _427538_427538 ; 
   reg __427538_427538;
   reg _427539_427539 ; 
   reg __427539_427539;
   reg _427540_427540 ; 
   reg __427540_427540;
   reg _427541_427541 ; 
   reg __427541_427541;
   reg _427542_427542 ; 
   reg __427542_427542;
   reg _427543_427543 ; 
   reg __427543_427543;
   reg _427544_427544 ; 
   reg __427544_427544;
   reg _427545_427545 ; 
   reg __427545_427545;
   reg _427546_427546 ; 
   reg __427546_427546;
   reg _427547_427547 ; 
   reg __427547_427547;
   reg _427548_427548 ; 
   reg __427548_427548;
   reg _427549_427549 ; 
   reg __427549_427549;
   reg _427550_427550 ; 
   reg __427550_427550;
   reg _427551_427551 ; 
   reg __427551_427551;
   reg _427552_427552 ; 
   reg __427552_427552;
   reg _427553_427553 ; 
   reg __427553_427553;
   reg _427554_427554 ; 
   reg __427554_427554;
   reg _427555_427555 ; 
   reg __427555_427555;
   reg _427556_427556 ; 
   reg __427556_427556;
   reg _427557_427557 ; 
   reg __427557_427557;
   reg _427558_427558 ; 
   reg __427558_427558;
   reg _427559_427559 ; 
   reg __427559_427559;
   reg _427560_427560 ; 
   reg __427560_427560;
   reg _427561_427561 ; 
   reg __427561_427561;
   reg _427562_427562 ; 
   reg __427562_427562;
   reg _427563_427563 ; 
   reg __427563_427563;
   reg _427564_427564 ; 
   reg __427564_427564;
   reg _427565_427565 ; 
   reg __427565_427565;
   reg _427566_427566 ; 
   reg __427566_427566;
   reg _427567_427567 ; 
   reg __427567_427567;
   reg _427568_427568 ; 
   reg __427568_427568;
   reg _427569_427569 ; 
   reg __427569_427569;
   reg _427570_427570 ; 
   reg __427570_427570;
   reg _427571_427571 ; 
   reg __427571_427571;
   reg _427572_427572 ; 
   reg __427572_427572;
   reg _427573_427573 ; 
   reg __427573_427573;
   reg _427574_427574 ; 
   reg __427574_427574;
   reg _427575_427575 ; 
   reg __427575_427575;
   reg _427576_427576 ; 
   reg __427576_427576;
   reg _427577_427577 ; 
   reg __427577_427577;
   reg _427578_427578 ; 
   reg __427578_427578;
   reg _427579_427579 ; 
   reg __427579_427579;
   reg _427580_427580 ; 
   reg __427580_427580;
   reg _427581_427581 ; 
   reg __427581_427581;
   reg _427582_427582 ; 
   reg __427582_427582;
   reg _427583_427583 ; 
   reg __427583_427583;
   reg _427584_427584 ; 
   reg __427584_427584;
   reg _427585_427585 ; 
   reg __427585_427585;
   reg _427586_427586 ; 
   reg __427586_427586;
   reg _427587_427587 ; 
   reg __427587_427587;
   reg _427588_427588 ; 
   reg __427588_427588;
   reg _427589_427589 ; 
   reg __427589_427589;
   reg _427590_427590 ; 
   reg __427590_427590;
   reg _427591_427591 ; 
   reg __427591_427591;
   reg _427592_427592 ; 
   reg __427592_427592;
   reg _427593_427593 ; 
   reg __427593_427593;
   reg _427594_427594 ; 
   reg __427594_427594;
   reg _427595_427595 ; 
   reg __427595_427595;
   reg _427596_427596 ; 
   reg __427596_427596;
   reg _427597_427597 ; 
   reg __427597_427597;
   reg _427598_427598 ; 
   reg __427598_427598;
   reg _427599_427599 ; 
   reg __427599_427599;
   reg _427600_427600 ; 
   reg __427600_427600;
   reg _427601_427601 ; 
   reg __427601_427601;
   reg _427602_427602 ; 
   reg __427602_427602;
   reg _427603_427603 ; 
   reg __427603_427603;
   reg _427604_427604 ; 
   reg __427604_427604;
   reg _427605_427605 ; 
   reg __427605_427605;
   reg _427606_427606 ; 
   reg __427606_427606;
   reg _427607_427607 ; 
   reg __427607_427607;
   reg _427608_427608 ; 
   reg __427608_427608;
   reg _427609_427609 ; 
   reg __427609_427609;
   reg _427610_427610 ; 
   reg __427610_427610;
   reg _427611_427611 ; 
   reg __427611_427611;
   reg _427612_427612 ; 
   reg __427612_427612;
   reg _427613_427613 ; 
   reg __427613_427613;
   reg _427614_427614 ; 
   reg __427614_427614;
   reg _427615_427615 ; 
   reg __427615_427615;
   reg _427616_427616 ; 
   reg __427616_427616;
   reg _427617_427617 ; 
   reg __427617_427617;
   reg _427618_427618 ; 
   reg __427618_427618;
   reg _427619_427619 ; 
   reg __427619_427619;
   reg _427620_427620 ; 
   reg __427620_427620;
   reg _427621_427621 ; 
   reg __427621_427621;
   reg _427622_427622 ; 
   reg __427622_427622;
   reg _427623_427623 ; 
   reg __427623_427623;
   reg _427624_427624 ; 
   reg __427624_427624;
   reg _427625_427625 ; 
   reg __427625_427625;
   reg _427626_427626 ; 
   reg __427626_427626;
   reg _427627_427627 ; 
   reg __427627_427627;
   reg _427628_427628 ; 
   reg __427628_427628;
   reg _427629_427629 ; 
   reg __427629_427629;
   reg _427630_427630 ; 
   reg __427630_427630;
   reg _427631_427631 ; 
   reg __427631_427631;
   reg _427632_427632 ; 
   reg __427632_427632;
   reg _427633_427633 ; 
   reg __427633_427633;
   reg _427634_427634 ; 
   reg __427634_427634;
   reg _427635_427635 ; 
   reg __427635_427635;
   reg _427636_427636 ; 
   reg __427636_427636;
   reg _427637_427637 ; 
   reg __427637_427637;
   reg _427638_427638 ; 
   reg __427638_427638;
   reg _427639_427639 ; 
   reg __427639_427639;
   reg _427640_427640 ; 
   reg __427640_427640;
   reg _427641_427641 ; 
   reg __427641_427641;
   reg _427642_427642 ; 
   reg __427642_427642;
   reg _427643_427643 ; 
   reg __427643_427643;
   reg _427644_427644 ; 
   reg __427644_427644;
   reg _427645_427645 ; 
   reg __427645_427645;
   reg _427646_427646 ; 
   reg __427646_427646;
   reg _427647_427647 ; 
   reg __427647_427647;
   reg _427648_427648 ; 
   reg __427648_427648;
   reg _427649_427649 ; 
   reg __427649_427649;
   reg _427650_427650 ; 
   reg __427650_427650;
   reg _427651_427651 ; 
   reg __427651_427651;
   reg _427652_427652 ; 
   reg __427652_427652;
   reg _427653_427653 ; 
   reg __427653_427653;
   reg _427654_427654 ; 
   reg __427654_427654;
   reg _427655_427655 ; 
   reg __427655_427655;
   reg _427656_427656 ; 
   reg __427656_427656;
   reg _427657_427657 ; 
   reg __427657_427657;
   reg _427658_427658 ; 
   reg __427658_427658;
   reg _427659_427659 ; 
   reg __427659_427659;
   reg _427660_427660 ; 
   reg __427660_427660;
   reg _427661_427661 ; 
   reg __427661_427661;
   reg _427662_427662 ; 
   reg __427662_427662;
   reg _427663_427663 ; 
   reg __427663_427663;
   reg _427664_427664 ; 
   reg __427664_427664;
   reg _427665_427665 ; 
   reg __427665_427665;
   reg _427666_427666 ; 
   reg __427666_427666;
   reg _427667_427667 ; 
   reg __427667_427667;
   reg _427668_427668 ; 
   reg __427668_427668;
   reg _427669_427669 ; 
   reg __427669_427669;
   reg _427670_427670 ; 
   reg __427670_427670;
   reg _427671_427671 ; 
   reg __427671_427671;
   reg _427672_427672 ; 
   reg __427672_427672;
   reg _427673_427673 ; 
   reg __427673_427673;
   reg _427674_427674 ; 
   reg __427674_427674;
   reg _427675_427675 ; 
   reg __427675_427675;
   reg _427676_427676 ; 
   reg __427676_427676;
   reg _427677_427677 ; 
   reg __427677_427677;
   reg _427678_427678 ; 
   reg __427678_427678;
   reg _427679_427679 ; 
   reg __427679_427679;
   reg _427680_427680 ; 
   reg __427680_427680;
   reg _427681_427681 ; 
   reg __427681_427681;
   reg _427682_427682 ; 
   reg __427682_427682;
   reg _427683_427683 ; 
   reg __427683_427683;
   reg _427684_427684 ; 
   reg __427684_427684;
   reg _427685_427685 ; 
   reg __427685_427685;
   reg _427686_427686 ; 
   reg __427686_427686;
   reg _427687_427687 ; 
   reg __427687_427687;
   reg _427688_427688 ; 
   reg __427688_427688;
   reg _427689_427689 ; 
   reg __427689_427689;
   reg _427690_427690 ; 
   reg __427690_427690;
   reg _427691_427691 ; 
   reg __427691_427691;
   reg _427692_427692 ; 
   reg __427692_427692;
   reg _427693_427693 ; 
   reg __427693_427693;
   reg _427694_427694 ; 
   reg __427694_427694;
   reg _427695_427695 ; 
   reg __427695_427695;
   reg _427696_427696 ; 
   reg __427696_427696;
   reg _427697_427697 ; 
   reg __427697_427697;
   reg _427698_427698 ; 
   reg __427698_427698;
   reg _427699_427699 ; 
   reg __427699_427699;
   reg _427700_427700 ; 
   reg __427700_427700;
   reg _427701_427701 ; 
   reg __427701_427701;
   reg _427702_427702 ; 
   reg __427702_427702;
   reg _427703_427703 ; 
   reg __427703_427703;
   reg _427704_427704 ; 
   reg __427704_427704;
   reg _427705_427705 ; 
   reg __427705_427705;
   reg _427706_427706 ; 
   reg __427706_427706;
   reg _427707_427707 ; 
   reg __427707_427707;
   reg _427708_427708 ; 
   reg __427708_427708;
   reg _427709_427709 ; 
   reg __427709_427709;
   reg _427710_427710 ; 
   reg __427710_427710;
   reg _427711_427711 ; 
   reg __427711_427711;
   reg _427712_427712 ; 
   reg __427712_427712;
   reg _427713_427713 ; 
   reg __427713_427713;
   reg _427714_427714 ; 
   reg __427714_427714;
   reg _427715_427715 ; 
   reg __427715_427715;
   reg _427716_427716 ; 
   reg __427716_427716;
   reg _427717_427717 ; 
   reg __427717_427717;
   reg _427718_427718 ; 
   reg __427718_427718;
   reg _427719_427719 ; 
   reg __427719_427719;
   reg _427720_427720 ; 
   reg __427720_427720;
   reg _427721_427721 ; 
   reg __427721_427721;
   reg _427722_427722 ; 
   reg __427722_427722;
   reg _427723_427723 ; 
   reg __427723_427723;
   reg _427724_427724 ; 
   reg __427724_427724;
   reg _427725_427725 ; 
   reg __427725_427725;
   reg _427726_427726 ; 
   reg __427726_427726;
   reg _427727_427727 ; 
   reg __427727_427727;
   reg _427728_427728 ; 
   reg __427728_427728;
   reg _427729_427729 ; 
   reg __427729_427729;
   reg _427730_427730 ; 
   reg __427730_427730;
   reg _427731_427731 ; 
   reg __427731_427731;
   reg _427732_427732 ; 
   reg __427732_427732;
   reg _427733_427733 ; 
   reg __427733_427733;
   reg _427734_427734 ; 
   reg __427734_427734;
   reg _427735_427735 ; 
   reg __427735_427735;
   reg _427736_427736 ; 
   reg __427736_427736;
   reg _427737_427737 ; 
   reg __427737_427737;
   reg _427738_427738 ; 
   reg __427738_427738;
   reg _427739_427739 ; 
   reg __427739_427739;
   reg _427740_427740 ; 
   reg __427740_427740;
   reg _427741_427741 ; 
   reg __427741_427741;
   reg _427742_427742 ; 
   reg __427742_427742;
   reg _427743_427743 ; 
   reg __427743_427743;
   reg _427744_427744 ; 
   reg __427744_427744;
   reg _427745_427745 ; 
   reg __427745_427745;
   reg _427746_427746 ; 
   reg __427746_427746;
   reg _427747_427747 ; 
   reg __427747_427747;
   reg _427748_427748 ; 
   reg __427748_427748;
   reg _427749_427749 ; 
   reg __427749_427749;
   reg _427750_427750 ; 
   reg __427750_427750;
   reg _427751_427751 ; 
   reg __427751_427751;
   reg _427752_427752 ; 
   reg __427752_427752;
   reg _427753_427753 ; 
   reg __427753_427753;
   reg _427754_427754 ; 
   reg __427754_427754;
   reg _427755_427755 ; 
   reg __427755_427755;
   reg _427756_427756 ; 
   reg __427756_427756;
   reg _427757_427757 ; 
   reg __427757_427757;
   reg _427758_427758 ; 
   reg __427758_427758;
   reg _427759_427759 ; 
   reg __427759_427759;
   reg _427760_427760 ; 
   reg __427760_427760;
   reg _427761_427761 ; 
   reg __427761_427761;
   reg _427762_427762 ; 
   reg __427762_427762;
   reg _427763_427763 ; 
   reg __427763_427763;
   reg _427764_427764 ; 
   reg __427764_427764;
   reg _427765_427765 ; 
   reg __427765_427765;
   reg _427766_427766 ; 
   reg __427766_427766;
   reg _427767_427767 ; 
   reg __427767_427767;
   reg _427768_427768 ; 
   reg __427768_427768;
   reg _427769_427769 ; 
   reg __427769_427769;
   reg _427770_427770 ; 
   reg __427770_427770;
   reg _427771_427771 ; 
   reg __427771_427771;
   reg _427772_427772 ; 
   reg __427772_427772;
   reg _427773_427773 ; 
   reg __427773_427773;
   reg _427774_427774 ; 
   reg __427774_427774;
   reg _427775_427775 ; 
   reg __427775_427775;
   reg _427776_427776 ; 
   reg __427776_427776;
   reg _427777_427777 ; 
   reg __427777_427777;
   reg _427778_427778 ; 
   reg __427778_427778;
   reg _427779_427779 ; 
   reg __427779_427779;
   reg _427780_427780 ; 
   reg __427780_427780;
   reg _427781_427781 ; 
   reg __427781_427781;
   reg _427782_427782 ; 
   reg __427782_427782;
   reg _427783_427783 ; 
   reg __427783_427783;
   reg _427784_427784 ; 
   reg __427784_427784;
   reg _427785_427785 ; 
   reg __427785_427785;
   reg _427786_427786 ; 
   reg __427786_427786;
   reg _427787_427787 ; 
   reg __427787_427787;
   reg _427788_427788 ; 
   reg __427788_427788;
   reg _427789_427789 ; 
   reg __427789_427789;
   reg _427790_427790 ; 
   reg __427790_427790;
   reg _427791_427791 ; 
   reg __427791_427791;
   reg _427792_427792 ; 
   reg __427792_427792;
   reg _427793_427793 ; 
   reg __427793_427793;
   reg _427794_427794 ; 
   reg __427794_427794;
   reg _427795_427795 ; 
   reg __427795_427795;
   reg _427796_427796 ; 
   reg __427796_427796;
   reg _427797_427797 ; 
   reg __427797_427797;
   reg _427798_427798 ; 
   reg __427798_427798;
   reg _427799_427799 ; 
   reg __427799_427799;
   reg _427800_427800 ; 
   reg __427800_427800;
   reg _427801_427801 ; 
   reg __427801_427801;
   reg _427802_427802 ; 
   reg __427802_427802;
   reg _427803_427803 ; 
   reg __427803_427803;
   reg _427804_427804 ; 
   reg __427804_427804;
   reg _427805_427805 ; 
   reg __427805_427805;
   reg _427806_427806 ; 
   reg __427806_427806;
   reg _427807_427807 ; 
   reg __427807_427807;
   reg _427808_427808 ; 
   reg __427808_427808;
   reg _427809_427809 ; 
   reg __427809_427809;
   reg _427810_427810 ; 
   reg __427810_427810;
   reg _427811_427811 ; 
   reg __427811_427811;
   reg _427812_427812 ; 
   reg __427812_427812;
   reg _427813_427813 ; 
   reg __427813_427813;
   reg _427814_427814 ; 
   reg __427814_427814;
   reg _427815_427815 ; 
   reg __427815_427815;
   reg _427816_427816 ; 
   reg __427816_427816;
   reg _427817_427817 ; 
   reg __427817_427817;
   reg _427818_427818 ; 
   reg __427818_427818;
   reg _427819_427819 ; 
   reg __427819_427819;
   reg _427820_427820 ; 
   reg __427820_427820;
   reg _427821_427821 ; 
   reg __427821_427821;
   reg _427822_427822 ; 
   reg __427822_427822;
   reg _427823_427823 ; 
   reg __427823_427823;
   reg _427824_427824 ; 
   reg __427824_427824;
   reg _427825_427825 ; 
   reg __427825_427825;
   reg _427826_427826 ; 
   reg __427826_427826;
   reg _427827_427827 ; 
   reg __427827_427827;
   reg _427828_427828 ; 
   reg __427828_427828;
   reg _427829_427829 ; 
   reg __427829_427829;
   reg _427830_427830 ; 
   reg __427830_427830;
   reg _427831_427831 ; 
   reg __427831_427831;
   reg _427832_427832 ; 
   reg __427832_427832;
   reg _427833_427833 ; 
   reg __427833_427833;
   reg _427834_427834 ; 
   reg __427834_427834;
   reg _427835_427835 ; 
   reg __427835_427835;
   reg _427836_427836 ; 
   reg __427836_427836;
   reg _427837_427837 ; 
   reg __427837_427837;
   reg _427838_427838 ; 
   reg __427838_427838;
   reg _427839_427839 ; 
   reg __427839_427839;
   reg _427840_427840 ; 
   reg __427840_427840;
   reg _427841_427841 ; 
   reg __427841_427841;
   reg _427842_427842 ; 
   reg __427842_427842;
   reg _427843_427843 ; 
   reg __427843_427843;
   reg _427844_427844 ; 
   reg __427844_427844;
   reg _427845_427845 ; 
   reg __427845_427845;
   reg _427846_427846 ; 
   reg __427846_427846;
   reg _427847_427847 ; 
   reg __427847_427847;
   reg _427848_427848 ; 
   reg __427848_427848;
   reg _427849_427849 ; 
   reg __427849_427849;
   reg _427850_427850 ; 
   reg __427850_427850;
   reg _427851_427851 ; 
   reg __427851_427851;
   reg _427852_427852 ; 
   reg __427852_427852;
   reg _427853_427853 ; 
   reg __427853_427853;
   reg _427854_427854 ; 
   reg __427854_427854;
   reg _427855_427855 ; 
   reg __427855_427855;
   reg _427856_427856 ; 
   reg __427856_427856;
   reg _427857_427857 ; 
   reg __427857_427857;
   reg _427858_427858 ; 
   reg __427858_427858;
   reg _427859_427859 ; 
   reg __427859_427859;
   reg _427860_427860 ; 
   reg __427860_427860;
   reg _427861_427861 ; 
   reg __427861_427861;
   reg _427862_427862 ; 
   reg __427862_427862;
   reg _427863_427863 ; 
   reg __427863_427863;
   reg _427864_427864 ; 
   reg __427864_427864;
   reg _427865_427865 ; 
   reg __427865_427865;
   reg _427866_427866 ; 
   reg __427866_427866;
   reg _427867_427867 ; 
   reg __427867_427867;
   reg _427868_427868 ; 
   reg __427868_427868;
   reg _427869_427869 ; 
   reg __427869_427869;
   reg _427870_427870 ; 
   reg __427870_427870;
   reg _427871_427871 ; 
   reg __427871_427871;
   reg _427872_427872 ; 
   reg __427872_427872;
   reg _427873_427873 ; 
   reg __427873_427873;
   reg _427874_427874 ; 
   reg __427874_427874;
   reg _427875_427875 ; 
   reg __427875_427875;
   reg _427876_427876 ; 
   reg __427876_427876;
   reg _427877_427877 ; 
   reg __427877_427877;
   reg _427878_427878 ; 
   reg __427878_427878;
   reg _427879_427879 ; 
   reg __427879_427879;
   reg _427880_427880 ; 
   reg __427880_427880;
   reg _427881_427881 ; 
   reg __427881_427881;
   reg _427882_427882 ; 
   reg __427882_427882;
   reg _427883_427883 ; 
   reg __427883_427883;
   reg _427884_427884 ; 
   reg __427884_427884;
   reg _427885_427885 ; 
   reg __427885_427885;
   reg _427886_427886 ; 
   reg __427886_427886;
   reg _427887_427887 ; 
   reg __427887_427887;
   reg _427888_427888 ; 
   reg __427888_427888;
   reg _427889_427889 ; 
   reg __427889_427889;
   reg _427890_427890 ; 
   reg __427890_427890;
   reg _427891_427891 ; 
   reg __427891_427891;
   reg _427892_427892 ; 
   reg __427892_427892;
   reg _427893_427893 ; 
   reg __427893_427893;
   reg _427894_427894 ; 
   reg __427894_427894;
   reg _427895_427895 ; 
   reg __427895_427895;
   reg _427896_427896 ; 
   reg __427896_427896;
   reg _427897_427897 ; 
   reg __427897_427897;
   reg _427898_427898 ; 
   reg __427898_427898;
   reg _427899_427899 ; 
   reg __427899_427899;
   reg _427900_427900 ; 
   reg __427900_427900;
   reg _427901_427901 ; 
   reg __427901_427901;
   reg _427902_427902 ; 
   reg __427902_427902;
   reg _427903_427903 ; 
   reg __427903_427903;
   reg _427904_427904 ; 
   reg __427904_427904;
   reg _427905_427905 ; 
   reg __427905_427905;
   reg _427906_427906 ; 
   reg __427906_427906;
   reg _427907_427907 ; 
   reg __427907_427907;
   reg _427908_427908 ; 
   reg __427908_427908;
   reg _427909_427909 ; 
   reg __427909_427909;
   reg _427910_427910 ; 
   reg __427910_427910;
   reg _427911_427911 ; 
   reg __427911_427911;
   reg _427912_427912 ; 
   reg __427912_427912;
   reg _427913_427913 ; 
   reg __427913_427913;
   reg _427914_427914 ; 
   reg __427914_427914;
   reg _427915_427915 ; 
   reg __427915_427915;
   reg _427916_427916 ; 
   reg __427916_427916;
   reg _427917_427917 ; 
   reg __427917_427917;
   reg _427918_427918 ; 
   reg __427918_427918;
   reg _427919_427919 ; 
   reg __427919_427919;
   reg _427920_427920 ; 
   reg __427920_427920;
   reg _427921_427921 ; 
   reg __427921_427921;
   reg _427922_427922 ; 
   reg __427922_427922;
   reg _427923_427923 ; 
   reg __427923_427923;
   reg _427924_427924 ; 
   reg __427924_427924;
   reg _427925_427925 ; 
   reg __427925_427925;
   reg _427926_427926 ; 
   reg __427926_427926;
   reg _427927_427927 ; 
   reg __427927_427927;
   reg _427928_427928 ; 
   reg __427928_427928;
   reg _427929_427929 ; 
   reg __427929_427929;
   reg _427930_427930 ; 
   reg __427930_427930;
   reg _427931_427931 ; 
   reg __427931_427931;
   reg _427932_427932 ; 
   reg __427932_427932;
   reg _427933_427933 ; 
   reg __427933_427933;
   reg _427934_427934 ; 
   reg __427934_427934;
   reg _427935_427935 ; 
   reg __427935_427935;
   reg _427936_427936 ; 
   reg __427936_427936;
   reg _427937_427937 ; 
   reg __427937_427937;
   reg _427938_427938 ; 
   reg __427938_427938;
   reg _427939_427939 ; 
   reg __427939_427939;
   reg _427940_427940 ; 
   reg __427940_427940;
   reg _427941_427941 ; 
   reg __427941_427941;
   reg _427942_427942 ; 
   reg __427942_427942;
   reg _427943_427943 ; 
   reg __427943_427943;
   reg _427944_427944 ; 
   reg __427944_427944;
   reg _427945_427945 ; 
   reg __427945_427945;
   reg _427946_427946 ; 
   reg __427946_427946;
   reg _427947_427947 ; 
   reg __427947_427947;
   reg _427948_427948 ; 
   reg __427948_427948;
   reg _427949_427949 ; 
   reg __427949_427949;
   reg _427950_427950 ; 
   reg __427950_427950;
   reg _427951_427951 ; 
   reg __427951_427951;
   reg _427952_427952 ; 
   reg __427952_427952;
   reg _427953_427953 ; 
   reg __427953_427953;
   reg _427954_427954 ; 
   reg __427954_427954;
   reg _427955_427955 ; 
   reg __427955_427955;
   reg _427956_427956 ; 
   reg __427956_427956;
   reg _427957_427957 ; 
   reg __427957_427957;
   reg _427958_427958 ; 
   reg __427958_427958;
   reg _427959_427959 ; 
   reg __427959_427959;
   reg _427960_427960 ; 
   reg __427960_427960;
   reg _427961_427961 ; 
   reg __427961_427961;
   reg _427962_427962 ; 
   reg __427962_427962;
   reg _427963_427963 ; 
   reg __427963_427963;
   reg _427964_427964 ; 
   reg __427964_427964;
   reg _427965_427965 ; 
   reg __427965_427965;
   reg _427966_427966 ; 
   reg __427966_427966;
   reg _427967_427967 ; 
   reg __427967_427967;
   reg _427968_427968 ; 
   reg __427968_427968;
   reg _427969_427969 ; 
   reg __427969_427969;
   reg _427970_427970 ; 
   reg __427970_427970;
   reg _427971_427971 ; 
   reg __427971_427971;
   reg _427972_427972 ; 
   reg __427972_427972;
   reg _427973_427973 ; 
   reg __427973_427973;
   reg _427974_427974 ; 
   reg __427974_427974;
   reg _427975_427975 ; 
   reg __427975_427975;
   reg _427976_427976 ; 
   reg __427976_427976;
   reg _427977_427977 ; 
   reg __427977_427977;
   reg _427978_427978 ; 
   reg __427978_427978;
   reg _427979_427979 ; 
   reg __427979_427979;
   reg _427980_427980 ; 
   reg __427980_427980;
   reg _427981_427981 ; 
   reg __427981_427981;
   reg _427982_427982 ; 
   reg __427982_427982;
   reg _427983_427983 ; 
   reg __427983_427983;
   reg _427984_427984 ; 
   reg __427984_427984;
   reg _427985_427985 ; 
   reg __427985_427985;
   reg _427986_427986 ; 
   reg __427986_427986;
   reg _427987_427987 ; 
   reg __427987_427987;
   reg _427988_427988 ; 
   reg __427988_427988;
   reg _427989_427989 ; 
   reg __427989_427989;
   reg _427990_427990 ; 
   reg __427990_427990;
   reg _427991_427991 ; 
   reg __427991_427991;
   reg _427992_427992 ; 
   reg __427992_427992;
   reg _427993_427993 ; 
   reg __427993_427993;
   reg _427994_427994 ; 
   reg __427994_427994;
   reg _427995_427995 ; 
   reg __427995_427995;
   reg _427996_427996 ; 
   reg __427996_427996;
   reg _427997_427997 ; 
   reg __427997_427997;
   reg _427998_427998 ; 
   reg __427998_427998;
   reg _427999_427999 ; 
   reg __427999_427999;
   reg _428000_428000 ; 
   reg __428000_428000;
   reg _428001_428001 ; 
   reg __428001_428001;
   reg _428002_428002 ; 
   reg __428002_428002;
   reg _428003_428003 ; 
   reg __428003_428003;
   reg _428004_428004 ; 
   reg __428004_428004;
   reg _428005_428005 ; 
   reg __428005_428005;
   reg _428006_428006 ; 
   reg __428006_428006;
   reg _428007_428007 ; 
   reg __428007_428007;
   reg _428008_428008 ; 
   reg __428008_428008;
   reg _428009_428009 ; 
   reg __428009_428009;
   reg _428010_428010 ; 
   reg __428010_428010;
   reg _428011_428011 ; 
   reg __428011_428011;
   reg _428012_428012 ; 
   reg __428012_428012;
   reg _428013_428013 ; 
   reg __428013_428013;
   reg _428014_428014 ; 
   reg __428014_428014;
   reg _428015_428015 ; 
   reg __428015_428015;
   reg _428016_428016 ; 
   reg __428016_428016;
   reg _428017_428017 ; 
   reg __428017_428017;
   reg _428018_428018 ; 
   reg __428018_428018;
   reg _428019_428019 ; 
   reg __428019_428019;
   reg _428020_428020 ; 
   reg __428020_428020;
   reg _428021_428021 ; 
   reg __428021_428021;
   reg _428022_428022 ; 
   reg __428022_428022;
   reg _428023_428023 ; 
   reg __428023_428023;
   reg _428024_428024 ; 
   reg __428024_428024;
   reg _428025_428025 ; 
   reg __428025_428025;
   reg _428026_428026 ; 
   reg __428026_428026;
   reg _428027_428027 ; 
   reg __428027_428027;
   reg _428028_428028 ; 
   reg __428028_428028;
   reg _428029_428029 ; 
   reg __428029_428029;
   reg _428030_428030 ; 
   reg __428030_428030;
   reg _428031_428031 ; 
   reg __428031_428031;
   reg _428032_428032 ; 
   reg __428032_428032;
   reg _428033_428033 ; 
   reg __428033_428033;
   reg _428034_428034 ; 
   reg __428034_428034;
   reg _428035_428035 ; 
   reg __428035_428035;
   reg _428036_428036 ; 
   reg __428036_428036;
   reg _428037_428037 ; 
   reg __428037_428037;
   reg _428038_428038 ; 
   reg __428038_428038;
   reg _428039_428039 ; 
   reg __428039_428039;
   reg _428040_428040 ; 
   reg __428040_428040;
   reg _428041_428041 ; 
   reg __428041_428041;
   reg _428042_428042 ; 
   reg __428042_428042;
   reg _428043_428043 ; 
   reg __428043_428043;
   reg _428044_428044 ; 
   reg __428044_428044;
   reg _428045_428045 ; 
   reg __428045_428045;
   reg _428046_428046 ; 
   reg __428046_428046;
   reg _428047_428047 ; 
   reg __428047_428047;
   reg _428048_428048 ; 
   reg __428048_428048;
   reg _428049_428049 ; 
   reg __428049_428049;
   reg _428050_428050 ; 
   reg __428050_428050;
   reg _428051_428051 ; 
   reg __428051_428051;
   reg _428052_428052 ; 
   reg __428052_428052;
   reg _428053_428053 ; 
   reg __428053_428053;
   reg _428054_428054 ; 
   reg __428054_428054;
   reg _428055_428055 ; 
   reg __428055_428055;
   reg _428056_428056 ; 
   reg __428056_428056;
   reg _428057_428057 ; 
   reg __428057_428057;
   reg _428058_428058 ; 
   reg __428058_428058;
   reg _428059_428059 ; 
   reg __428059_428059;
   reg _428060_428060 ; 
   reg __428060_428060;
   reg _428061_428061 ; 
   reg __428061_428061;
   reg _428062_428062 ; 
   reg __428062_428062;
   reg _428063_428063 ; 
   reg __428063_428063;
   reg _428064_428064 ; 
   reg __428064_428064;
   reg _428065_428065 ; 
   reg __428065_428065;
   reg _428066_428066 ; 
   reg __428066_428066;
   reg _428067_428067 ; 
   reg __428067_428067;
   reg _428068_428068 ; 
   reg __428068_428068;
   reg _428069_428069 ; 
   reg __428069_428069;
   reg _428070_428070 ; 
   reg __428070_428070;
   reg _428071_428071 ; 
   reg __428071_428071;
   reg _428072_428072 ; 
   reg __428072_428072;
   reg _428073_428073 ; 
   reg __428073_428073;
   reg _428074_428074 ; 
   reg __428074_428074;
   reg _428075_428075 ; 
   reg __428075_428075;
   reg _428076_428076 ; 
   reg __428076_428076;
   reg _428077_428077 ; 
   reg __428077_428077;
   reg _428078_428078 ; 
   reg __428078_428078;
   reg _428079_428079 ; 
   reg __428079_428079;
   reg _428080_428080 ; 
   reg __428080_428080;
   reg _428081_428081 ; 
   reg __428081_428081;
   reg _428082_428082 ; 
   reg __428082_428082;
   reg _428083_428083 ; 
   reg __428083_428083;
   reg _428084_428084 ; 
   reg __428084_428084;
   reg _428085_428085 ; 
   reg __428085_428085;
   reg _428086_428086 ; 
   reg __428086_428086;
   reg _428087_428087 ; 
   reg __428087_428087;
   reg _428088_428088 ; 
   reg __428088_428088;
   reg _428089_428089 ; 
   reg __428089_428089;
   reg _428090_428090 ; 
   reg __428090_428090;
   reg _428091_428091 ; 
   reg __428091_428091;
   reg _428092_428092 ; 
   reg __428092_428092;
   reg _428093_428093 ; 
   reg __428093_428093;
   reg _428094_428094 ; 
   reg __428094_428094;
   reg _428095_428095 ; 
   reg __428095_428095;
   reg _428096_428096 ; 
   reg __428096_428096;
   reg _428097_428097 ; 
   reg __428097_428097;
   reg _428098_428098 ; 
   reg __428098_428098;
   reg _428099_428099 ; 
   reg __428099_428099;
   reg _428100_428100 ; 
   reg __428100_428100;
   reg _428101_428101 ; 
   reg __428101_428101;
   reg _428102_428102 ; 
   reg __428102_428102;
   reg _428103_428103 ; 
   reg __428103_428103;
   reg _428104_428104 ; 
   reg __428104_428104;
   reg _428105_428105 ; 
   reg __428105_428105;
   reg _428106_428106 ; 
   reg __428106_428106;
   reg _428107_428107 ; 
   reg __428107_428107;
   reg _428108_428108 ; 
   reg __428108_428108;
   reg _428109_428109 ; 
   reg __428109_428109;
   reg _428110_428110 ; 
   reg __428110_428110;
   reg _428111_428111 ; 
   reg __428111_428111;
   reg _428112_428112 ; 
   reg __428112_428112;
   reg _428113_428113 ; 
   reg __428113_428113;
   reg _428114_428114 ; 
   reg __428114_428114;
   reg _428115_428115 ; 
   reg __428115_428115;
   reg _428116_428116 ; 
   reg __428116_428116;
   reg _428117_428117 ; 
   reg __428117_428117;
   reg _428118_428118 ; 
   reg __428118_428118;
   reg _428119_428119 ; 
   reg __428119_428119;
   reg _428120_428120 ; 
   reg __428120_428120;
   reg _428121_428121 ; 
   reg __428121_428121;
   reg _428122_428122 ; 
   reg __428122_428122;
   reg _428123_428123 ; 
   reg __428123_428123;
   reg _428124_428124 ; 
   reg __428124_428124;
   reg _428125_428125 ; 
   reg __428125_428125;
   reg _428126_428126 ; 
   reg __428126_428126;
   reg _428127_428127 ; 
   reg __428127_428127;
   reg _428128_428128 ; 
   reg __428128_428128;
   reg _428129_428129 ; 
   reg __428129_428129;
   reg _428130_428130 ; 
   reg __428130_428130;
   reg _428131_428131 ; 
   reg __428131_428131;
   reg _428132_428132 ; 
   reg __428132_428132;
   reg _428133_428133 ; 
   reg __428133_428133;
   reg _428134_428134 ; 
   reg __428134_428134;
   reg _428135_428135 ; 
   reg __428135_428135;
   reg _428136_428136 ; 
   reg __428136_428136;
   reg _428137_428137 ; 
   reg __428137_428137;
   reg _428138_428138 ; 
   reg __428138_428138;
   reg _428139_428139 ; 
   reg __428139_428139;
   reg _428140_428140 ; 
   reg __428140_428140;
   reg _428141_428141 ; 
   reg __428141_428141;
   reg _428142_428142 ; 
   reg __428142_428142;
   reg _428143_428143 ; 
   reg __428143_428143;
   reg _428144_428144 ; 
   reg __428144_428144;
   reg _428145_428145 ; 
   reg __428145_428145;
   reg _428146_428146 ; 
   reg __428146_428146;
   reg _428147_428147 ; 
   reg __428147_428147;
   reg _428148_428148 ; 
   reg __428148_428148;
   reg _428149_428149 ; 
   reg __428149_428149;
   reg _428150_428150 ; 
   reg __428150_428150;
   reg _428151_428151 ; 
   reg __428151_428151;
   reg _428152_428152 ; 
   reg __428152_428152;
   reg _428153_428153 ; 
   reg __428153_428153;
   reg _428154_428154 ; 
   reg __428154_428154;
   reg _428155_428155 ; 
   reg __428155_428155;
   reg _428156_428156 ; 
   reg __428156_428156;
   reg _428157_428157 ; 
   reg __428157_428157;
   reg _428158_428158 ; 
   reg __428158_428158;
   reg _428159_428159 ; 
   reg __428159_428159;
   reg _428160_428160 ; 
   reg __428160_428160;
   reg _428161_428161 ; 
   reg __428161_428161;
   reg _428162_428162 ; 
   reg __428162_428162;
   reg _428163_428163 ; 
   reg __428163_428163;
   reg _428164_428164 ; 
   reg __428164_428164;
   reg _428165_428165 ; 
   reg __428165_428165;
   reg _428166_428166 ; 
   reg __428166_428166;
   reg _428167_428167 ; 
   reg __428167_428167;
   reg _428168_428168 ; 
   reg __428168_428168;
   reg _428169_428169 ; 
   reg __428169_428169;
   reg _428170_428170 ; 
   reg __428170_428170;
   reg _428171_428171 ; 
   reg __428171_428171;
   reg _428172_428172 ; 
   reg __428172_428172;
   reg _428173_428173 ; 
   reg __428173_428173;
   reg _428174_428174 ; 
   reg __428174_428174;
   reg _428175_428175 ; 
   reg __428175_428175;
   reg _428176_428176 ; 
   reg __428176_428176;
   reg _428177_428177 ; 
   reg __428177_428177;
   reg _428178_428178 ; 
   reg __428178_428178;
   reg _428179_428179 ; 
   reg __428179_428179;
   reg _428180_428180 ; 
   reg __428180_428180;
   reg _428181_428181 ; 
   reg __428181_428181;
   reg _428182_428182 ; 
   reg __428182_428182;
   reg _428183_428183 ; 
   reg __428183_428183;
   reg _428184_428184 ; 
   reg __428184_428184;
   reg _428185_428185 ; 
   reg __428185_428185;
   reg _428186_428186 ; 
   reg __428186_428186;
   reg _428187_428187 ; 
   reg __428187_428187;
   reg _428188_428188 ; 
   reg __428188_428188;
   reg _428189_428189 ; 
   reg __428189_428189;
   reg _428190_428190 ; 
   reg __428190_428190;
   reg _428191_428191 ; 
   reg __428191_428191;
   reg _428192_428192 ; 
   reg __428192_428192;
   reg _428193_428193 ; 
   reg __428193_428193;
   reg _428194_428194 ; 
   reg __428194_428194;
   reg _428195_428195 ; 
   reg __428195_428195;
   reg _428196_428196 ; 
   reg __428196_428196;
   reg _428197_428197 ; 
   reg __428197_428197;
   reg _428198_428198 ; 
   reg __428198_428198;
   reg _428199_428199 ; 
   reg __428199_428199;
   reg _428200_428200 ; 
   reg __428200_428200;
   reg _428201_428201 ; 
   reg __428201_428201;
   reg _428202_428202 ; 
   reg __428202_428202;
   reg _428203_428203 ; 
   reg __428203_428203;
   reg _428204_428204 ; 
   reg __428204_428204;
   reg _428205_428205 ; 
   reg __428205_428205;
   reg _428206_428206 ; 
   reg __428206_428206;
   reg _428207_428207 ; 
   reg __428207_428207;
   reg _428208_428208 ; 
   reg __428208_428208;
   reg _428209_428209 ; 
   reg __428209_428209;
   reg _428210_428210 ; 
   reg __428210_428210;
   reg _428211_428211 ; 
   reg __428211_428211;
   reg _428212_428212 ; 
   reg __428212_428212;
   reg _428213_428213 ; 
   reg __428213_428213;
   reg _428214_428214 ; 
   reg __428214_428214;
   reg _428215_428215 ; 
   reg __428215_428215;
   reg _428216_428216 ; 
   reg __428216_428216;
   reg _428217_428217 ; 
   reg __428217_428217;
   reg _428218_428218 ; 
   reg __428218_428218;
   reg _428219_428219 ; 
   reg __428219_428219;
   reg _428220_428220 ; 
   reg __428220_428220;
   reg _428221_428221 ; 
   reg __428221_428221;
   reg _428222_428222 ; 
   reg __428222_428222;
   reg _428223_428223 ; 
   reg __428223_428223;
   reg _428224_428224 ; 
   reg __428224_428224;
   reg _428225_428225 ; 
   reg __428225_428225;
   reg _428226_428226 ; 
   reg __428226_428226;
   reg _428227_428227 ; 
   reg __428227_428227;
   reg _428228_428228 ; 
   reg __428228_428228;
   reg _428229_428229 ; 
   reg __428229_428229;
   reg _428230_428230 ; 
   reg __428230_428230;
   reg _428231_428231 ; 
   reg __428231_428231;
   reg _428232_428232 ; 
   reg __428232_428232;
   reg _428233_428233 ; 
   reg __428233_428233;
   reg _428234_428234 ; 
   reg __428234_428234;
   reg _428235_428235 ; 
   reg __428235_428235;
   reg _428236_428236 ; 
   reg __428236_428236;
   reg _428237_428237 ; 
   reg __428237_428237;
   reg _428238_428238 ; 
   reg __428238_428238;
   reg _428239_428239 ; 
   reg __428239_428239;
   reg _428240_428240 ; 
   reg __428240_428240;
   reg _428241_428241 ; 
   reg __428241_428241;
   reg _428242_428242 ; 
   reg __428242_428242;
   reg _428243_428243 ; 
   reg __428243_428243;
   reg _428244_428244 ; 
   reg __428244_428244;
   reg _428245_428245 ; 
   reg __428245_428245;
   reg _428246_428246 ; 
   reg __428246_428246;
   reg _428247_428247 ; 
   reg __428247_428247;
   reg _428248_428248 ; 
   reg __428248_428248;
   reg _428249_428249 ; 
   reg __428249_428249;
   reg _428250_428250 ; 
   reg __428250_428250;
   reg _428251_428251 ; 
   reg __428251_428251;
   reg _428252_428252 ; 
   reg __428252_428252;
   reg _428253_428253 ; 
   reg __428253_428253;
   reg _428254_428254 ; 
   reg __428254_428254;
   reg _428255_428255 ; 
   reg __428255_428255;
   reg _428256_428256 ; 
   reg __428256_428256;
   reg _428257_428257 ; 
   reg __428257_428257;
   reg _428258_428258 ; 
   reg __428258_428258;
   reg _428259_428259 ; 
   reg __428259_428259;
   reg _428260_428260 ; 
   reg __428260_428260;
   reg _428261_428261 ; 
   reg __428261_428261;
   reg _428262_428262 ; 
   reg __428262_428262;
   reg _428263_428263 ; 
   reg __428263_428263;
   reg _428264_428264 ; 
   reg __428264_428264;
   reg _428265_428265 ; 
   reg __428265_428265;
   reg _428266_428266 ; 
   reg __428266_428266;
   reg _428267_428267 ; 
   reg __428267_428267;
   reg _428268_428268 ; 
   reg __428268_428268;
   reg _428269_428269 ; 
   reg __428269_428269;
   reg _428270_428270 ; 
   reg __428270_428270;
   reg _428271_428271 ; 
   reg __428271_428271;
   reg _428272_428272 ; 
   reg __428272_428272;
   reg _428273_428273 ; 
   reg __428273_428273;
   reg _428274_428274 ; 
   reg __428274_428274;
   reg _428275_428275 ; 
   reg __428275_428275;
   reg _428276_428276 ; 
   reg __428276_428276;
   reg _428277_428277 ; 
   reg __428277_428277;
   reg _428278_428278 ; 
   reg __428278_428278;
   reg _428279_428279 ; 
   reg __428279_428279;
   reg _428280_428280 ; 
   reg __428280_428280;
   reg _428281_428281 ; 
   reg __428281_428281;
   reg _428282_428282 ; 
   reg __428282_428282;
   reg _428283_428283 ; 
   reg __428283_428283;
   reg _428284_428284 ; 
   reg __428284_428284;
   reg _428285_428285 ; 
   reg __428285_428285;
   reg _428286_428286 ; 
   reg __428286_428286;
   reg _428287_428287 ; 
   reg __428287_428287;
   reg _428288_428288 ; 
   reg __428288_428288;
   reg _428289_428289 ; 
   reg __428289_428289;
   reg _428290_428290 ; 
   reg __428290_428290;
   reg _428291_428291 ; 
   reg __428291_428291;
   reg _428292_428292 ; 
   reg __428292_428292;
   reg _428293_428293 ; 
   reg __428293_428293;
   reg _428294_428294 ; 
   reg __428294_428294;
   reg _428295_428295 ; 
   reg __428295_428295;
   reg _428296_428296 ; 
   reg __428296_428296;
   reg _428297_428297 ; 
   reg __428297_428297;
   reg _428298_428298 ; 
   reg __428298_428298;
   reg _428299_428299 ; 
   reg __428299_428299;
   reg _428300_428300 ; 
   reg __428300_428300;
   reg _428301_428301 ; 
   reg __428301_428301;
   reg _428302_428302 ; 
   reg __428302_428302;
   reg _428303_428303 ; 
   reg __428303_428303;
   reg _428304_428304 ; 
   reg __428304_428304;
   reg _428305_428305 ; 
   reg __428305_428305;
   reg _428306_428306 ; 
   reg __428306_428306;
   reg _428307_428307 ; 
   reg __428307_428307;
   reg _428308_428308 ; 
   reg __428308_428308;
   reg _428309_428309 ; 
   reg __428309_428309;
   reg _428310_428310 ; 
   reg __428310_428310;
   reg _428311_428311 ; 
   reg __428311_428311;
   reg _428312_428312 ; 
   reg __428312_428312;
   reg _428313_428313 ; 
   reg __428313_428313;
   reg _428314_428314 ; 
   reg __428314_428314;
   reg _428315_428315 ; 
   reg __428315_428315;
   reg _428316_428316 ; 
   reg __428316_428316;
   reg _428317_428317 ; 
   reg __428317_428317;
   reg _428318_428318 ; 
   reg __428318_428318;
   reg _428319_428319 ; 
   reg __428319_428319;
   reg _428320_428320 ; 
   reg __428320_428320;
   reg _428321_428321 ; 
   reg __428321_428321;
   reg _428322_428322 ; 
   reg __428322_428322;
   reg _428323_428323 ; 
   reg __428323_428323;
   reg _428324_428324 ; 
   reg __428324_428324;
   reg _428325_428325 ; 
   reg __428325_428325;
   reg _428326_428326 ; 
   reg __428326_428326;
   reg _428327_428327 ; 
   reg __428327_428327;
   reg _428328_428328 ; 
   reg __428328_428328;
   reg _428329_428329 ; 
   reg __428329_428329;
   reg _428330_428330 ; 
   reg __428330_428330;
   reg _428331_428331 ; 
   reg __428331_428331;
   reg _428332_428332 ; 
   reg __428332_428332;
   reg _428333_428333 ; 
   reg __428333_428333;
   reg _428334_428334 ; 
   reg __428334_428334;
   reg _428335_428335 ; 
   reg __428335_428335;
   reg _428336_428336 ; 
   reg __428336_428336;
   reg _428337_428337 ; 
   reg __428337_428337;
   reg _428338_428338 ; 
   reg __428338_428338;
   reg _428339_428339 ; 
   reg __428339_428339;
   reg _428340_428340 ; 
   reg __428340_428340;
   reg _428341_428341 ; 
   reg __428341_428341;
   reg _428342_428342 ; 
   reg __428342_428342;
   reg _428343_428343 ; 
   reg __428343_428343;
   reg _428344_428344 ; 
   reg __428344_428344;
   reg _428345_428345 ; 
   reg __428345_428345;
   reg _428346_428346 ; 
   reg __428346_428346;
   reg _428347_428347 ; 
   reg __428347_428347;
   reg _428348_428348 ; 
   reg __428348_428348;
   reg _428349_428349 ; 
   reg __428349_428349;
   reg _428350_428350 ; 
   reg __428350_428350;
   reg _428351_428351 ; 
   reg __428351_428351;
   reg _428352_428352 ; 
   reg __428352_428352;
   reg _428353_428353 ; 
   reg __428353_428353;
   reg _428354_428354 ; 
   reg __428354_428354;
   reg _428355_428355 ; 
   reg __428355_428355;
   reg _428356_428356 ; 
   reg __428356_428356;
   reg _428357_428357 ; 
   reg __428357_428357;
   reg _428358_428358 ; 
   reg __428358_428358;
   reg _428359_428359 ; 
   reg __428359_428359;
   reg _428360_428360 ; 
   reg __428360_428360;
   reg _428361_428361 ; 
   reg __428361_428361;
   reg _428362_428362 ; 
   reg __428362_428362;
   reg _428363_428363 ; 
   reg __428363_428363;
   reg _428364_428364 ; 
   reg __428364_428364;
   reg _428365_428365 ; 
   reg __428365_428365;
   reg _428366_428366 ; 
   reg __428366_428366;
   reg _428367_428367 ; 
   reg __428367_428367;
   reg _428368_428368 ; 
   reg __428368_428368;
   reg _428369_428369 ; 
   reg __428369_428369;
   reg _428370_428370 ; 
   reg __428370_428370;
   reg _428371_428371 ; 
   reg __428371_428371;
   reg _428372_428372 ; 
   reg __428372_428372;
   reg _428373_428373 ; 
   reg __428373_428373;
   reg _428374_428374 ; 
   reg __428374_428374;
   reg _428375_428375 ; 
   reg __428375_428375;
   reg _428376_428376 ; 
   reg __428376_428376;
   reg _428377_428377 ; 
   reg __428377_428377;
   reg _428378_428378 ; 
   reg __428378_428378;
   reg _428379_428379 ; 
   reg __428379_428379;
   reg _428380_428380 ; 
   reg __428380_428380;
   reg _428381_428381 ; 
   reg __428381_428381;
   reg _428382_428382 ; 
   reg __428382_428382;
   reg _428383_428383 ; 
   reg __428383_428383;
   reg _428384_428384 ; 
   reg __428384_428384;
   reg _428385_428385 ; 
   reg __428385_428385;
   reg _428386_428386 ; 
   reg __428386_428386;
   reg _428387_428387 ; 
   reg __428387_428387;
   reg _428388_428388 ; 
   reg __428388_428388;
   reg _428389_428389 ; 
   reg __428389_428389;
   reg _428390_428390 ; 
   reg __428390_428390;
   reg _428391_428391 ; 
   reg __428391_428391;
   reg _428392_428392 ; 
   reg __428392_428392;
   reg _428393_428393 ; 
   reg __428393_428393;
   reg _428394_428394 ; 
   reg __428394_428394;
   reg _428395_428395 ; 
   reg __428395_428395;
   reg _428396_428396 ; 
   reg __428396_428396;
   reg _428397_428397 ; 
   reg __428397_428397;
   reg _428398_428398 ; 
   reg __428398_428398;
   reg _428399_428399 ; 
   reg __428399_428399;
   reg _428400_428400 ; 
   reg __428400_428400;
   reg _428401_428401 ; 
   reg __428401_428401;
   reg _428402_428402 ; 
   reg __428402_428402;
   reg _428403_428403 ; 
   reg __428403_428403;
   reg _428404_428404 ; 
   reg __428404_428404;
   reg _428405_428405 ; 
   reg __428405_428405;
   reg _428406_428406 ; 
   reg __428406_428406;
   reg _428407_428407 ; 
   reg __428407_428407;
   reg _428408_428408 ; 
   reg __428408_428408;
   reg _428409_428409 ; 
   reg __428409_428409;
   reg _428410_428410 ; 
   reg __428410_428410;
   reg _428411_428411 ; 
   reg __428411_428411;
   reg _428412_428412 ; 
   reg __428412_428412;
   reg _428413_428413 ; 
   reg __428413_428413;
   reg _428414_428414 ; 
   reg __428414_428414;
   reg _428415_428415 ; 
   reg __428415_428415;
   reg _428416_428416 ; 
   reg __428416_428416;
   reg _428417_428417 ; 
   reg __428417_428417;
   reg _428418_428418 ; 
   reg __428418_428418;
   reg _428419_428419 ; 
   reg __428419_428419;
   reg _428420_428420 ; 
   reg __428420_428420;
   reg _428421_428421 ; 
   reg __428421_428421;
   reg _428422_428422 ; 
   reg __428422_428422;
   reg _428423_428423 ; 
   reg __428423_428423;
   reg _428424_428424 ; 
   reg __428424_428424;
   reg _428425_428425 ; 
   reg __428425_428425;
   reg _428426_428426 ; 
   reg __428426_428426;
   reg _428427_428427 ; 
   reg __428427_428427;
   reg _428428_428428 ; 
   reg __428428_428428;
   reg _428429_428429 ; 
   reg __428429_428429;
   reg _428430_428430 ; 
   reg __428430_428430;
   reg _428431_428431 ; 
   reg __428431_428431;
   reg _428432_428432 ; 
   reg __428432_428432;
   reg _428433_428433 ; 
   reg __428433_428433;
   reg _428434_428434 ; 
   reg __428434_428434;
   reg _428435_428435 ; 
   reg __428435_428435;
   reg _428436_428436 ; 
   reg __428436_428436;
   reg _428437_428437 ; 
   reg __428437_428437;
   reg _428438_428438 ; 
   reg __428438_428438;
   reg _428439_428439 ; 
   reg __428439_428439;
   reg _428440_428440 ; 
   reg __428440_428440;
   reg _428441_428441 ; 
   reg __428441_428441;
   reg _428442_428442 ; 
   reg __428442_428442;
   reg _428443_428443 ; 
   reg __428443_428443;
   reg _428444_428444 ; 
   reg __428444_428444;
   reg _428445_428445 ; 
   reg __428445_428445;
   reg _428446_428446 ; 
   reg __428446_428446;
   reg _428447_428447 ; 
   reg __428447_428447;
   reg _428448_428448 ; 
   reg __428448_428448;
   reg _428449_428449 ; 
   reg __428449_428449;
   reg _428450_428450 ; 
   reg __428450_428450;
   reg _428451_428451 ; 
   reg __428451_428451;
   reg _428452_428452 ; 
   reg __428452_428452;
   reg _428453_428453 ; 
   reg __428453_428453;
   reg _428454_428454 ; 
   reg __428454_428454;
   reg _428455_428455 ; 
   reg __428455_428455;
   reg _428456_428456 ; 
   reg __428456_428456;
   reg _428457_428457 ; 
   reg __428457_428457;
   reg _428458_428458 ; 
   reg __428458_428458;
   reg _428459_428459 ; 
   reg __428459_428459;
   reg _428460_428460 ; 
   reg __428460_428460;
   reg _428461_428461 ; 
   reg __428461_428461;
   reg _428462_428462 ; 
   reg __428462_428462;
   reg _428463_428463 ; 
   reg __428463_428463;
   reg _428464_428464 ; 
   reg __428464_428464;
   reg _428465_428465 ; 
   reg __428465_428465;
   reg _428466_428466 ; 
   reg __428466_428466;
   reg _428467_428467 ; 
   reg __428467_428467;
   reg _428468_428468 ; 
   reg __428468_428468;
   reg _428469_428469 ; 
   reg __428469_428469;
   reg _428470_428470 ; 
   reg __428470_428470;
   reg _428471_428471 ; 
   reg __428471_428471;
   reg _428472_428472 ; 
   reg __428472_428472;
   reg _428473_428473 ; 
   reg __428473_428473;
   reg _428474_428474 ; 
   reg __428474_428474;
   reg _428475_428475 ; 
   reg __428475_428475;
   reg _428476_428476 ; 
   reg __428476_428476;
   reg _428477_428477 ; 
   reg __428477_428477;
   reg _428478_428478 ; 
   reg __428478_428478;
   reg _428479_428479 ; 
   reg __428479_428479;
   reg _428480_428480 ; 
   reg __428480_428480;
   reg _428481_428481 ; 
   reg __428481_428481;
   reg _428482_428482 ; 
   reg __428482_428482;
   reg _428483_428483 ; 
   reg __428483_428483;
   reg _428484_428484 ; 
   reg __428484_428484;
   reg _428485_428485 ; 
   reg __428485_428485;
   reg _428486_428486 ; 
   reg __428486_428486;
   reg _428487_428487 ; 
   reg __428487_428487;
   reg _428488_428488 ; 
   reg __428488_428488;
   reg _428489_428489 ; 
   reg __428489_428489;
   reg _428490_428490 ; 
   reg __428490_428490;
   reg _428491_428491 ; 
   reg __428491_428491;
   reg _428492_428492 ; 
   reg __428492_428492;
   reg _428493_428493 ; 
   reg __428493_428493;
   reg _428494_428494 ; 
   reg __428494_428494;
   reg _428495_428495 ; 
   reg __428495_428495;
   reg _428496_428496 ; 
   reg __428496_428496;
   reg _428497_428497 ; 
   reg __428497_428497;
   reg _428498_428498 ; 
   reg __428498_428498;
   reg _428499_428499 ; 
   reg __428499_428499;
   reg _428500_428500 ; 
   reg __428500_428500;
   reg _428501_428501 ; 
   reg __428501_428501;
   reg _428502_428502 ; 
   reg __428502_428502;
   reg _428503_428503 ; 
   reg __428503_428503;
   reg _428504_428504 ; 
   reg __428504_428504;
   reg _428505_428505 ; 
   reg __428505_428505;
   reg _428506_428506 ; 
   reg __428506_428506;
   reg _428507_428507 ; 
   reg __428507_428507;
   reg _428508_428508 ; 
   reg __428508_428508;
   reg _428509_428509 ; 
   reg __428509_428509;
   reg _428510_428510 ; 
   reg __428510_428510;
   reg _428511_428511 ; 
   reg __428511_428511;
   reg _428512_428512 ; 
   reg __428512_428512;
   reg _428513_428513 ; 
   reg __428513_428513;
   reg _428514_428514 ; 
   reg __428514_428514;
   reg _428515_428515 ; 
   reg __428515_428515;
   reg _428516_428516 ; 
   reg __428516_428516;
   reg _428517_428517 ; 
   reg __428517_428517;
   reg _428518_428518 ; 
   reg __428518_428518;
   reg _428519_428519 ; 
   reg __428519_428519;
   reg _428520_428520 ; 
   reg __428520_428520;
   reg _428521_428521 ; 
   reg __428521_428521;
   reg _428522_428522 ; 
   reg __428522_428522;
   reg _428523_428523 ; 
   reg __428523_428523;
   reg _428524_428524 ; 
   reg __428524_428524;
   reg _428525_428525 ; 
   reg __428525_428525;
   reg _428526_428526 ; 
   reg __428526_428526;
   reg _428527_428527 ; 
   reg __428527_428527;
   reg _428528_428528 ; 
   reg __428528_428528;
   reg _428529_428529 ; 
   reg __428529_428529;
   reg _428530_428530 ; 
   reg __428530_428530;
   reg _428531_428531 ; 
   reg __428531_428531;
   reg _428532_428532 ; 
   reg __428532_428532;
   reg _428533_428533 ; 
   reg __428533_428533;
   reg _428534_428534 ; 
   reg __428534_428534;
   reg _428535_428535 ; 
   reg __428535_428535;
   reg _428536_428536 ; 
   reg __428536_428536;
   reg _428537_428537 ; 
   reg __428537_428537;
   reg _428538_428538 ; 
   reg __428538_428538;
   reg _428539_428539 ; 
   reg __428539_428539;
   reg _428540_428540 ; 
   reg __428540_428540;
   reg _428541_428541 ; 
   reg __428541_428541;
   reg _428542_428542 ; 
   reg __428542_428542;
   reg _428543_428543 ; 
   reg __428543_428543;
   reg _428544_428544 ; 
   reg __428544_428544;
   reg _428545_428545 ; 
   reg __428545_428545;
   reg _428546_428546 ; 
   reg __428546_428546;
   reg _428547_428547 ; 
   reg __428547_428547;
   reg _428548_428548 ; 
   reg __428548_428548;
   reg _428549_428549 ; 
   reg __428549_428549;
   reg _428550_428550 ; 
   reg __428550_428550;
   reg _428551_428551 ; 
   reg __428551_428551;
   reg _428552_428552 ; 
   reg __428552_428552;
   reg _428553_428553 ; 
   reg __428553_428553;
   reg _428554_428554 ; 
   reg __428554_428554;
   reg _428555_428555 ; 
   reg __428555_428555;
   reg _428556_428556 ; 
   reg __428556_428556;
   reg _428557_428557 ; 
   reg __428557_428557;
   reg _428558_428558 ; 
   reg __428558_428558;
   reg _428559_428559 ; 
   reg __428559_428559;
   reg _428560_428560 ; 
   reg __428560_428560;
   reg _428561_428561 ; 
   reg __428561_428561;
   reg _428562_428562 ; 
   reg __428562_428562;
   reg _428563_428563 ; 
   reg __428563_428563;
   reg _428564_428564 ; 
   reg __428564_428564;
   reg _428565_428565 ; 
   reg __428565_428565;
   reg _428566_428566 ; 
   reg __428566_428566;
   reg _428567_428567 ; 
   reg __428567_428567;
   reg _428568_428568 ; 
   reg __428568_428568;
   reg _428569_428569 ; 
   reg __428569_428569;
   reg _428570_428570 ; 
   reg __428570_428570;
   reg _428571_428571 ; 
   reg __428571_428571;
   reg _428572_428572 ; 
   reg __428572_428572;
   reg _428573_428573 ; 
   reg __428573_428573;
   reg _428574_428574 ; 
   reg __428574_428574;
   reg _428575_428575 ; 
   reg __428575_428575;
   reg _428576_428576 ; 
   reg __428576_428576;
   reg _428577_428577 ; 
   reg __428577_428577;
   reg _428578_428578 ; 
   reg __428578_428578;
   reg _428579_428579 ; 
   reg __428579_428579;
   reg _428580_428580 ; 
   reg __428580_428580;
   reg _428581_428581 ; 
   reg __428581_428581;
   reg _428582_428582 ; 
   reg __428582_428582;
   reg _428583_428583 ; 
   reg __428583_428583;
   reg _428584_428584 ; 
   reg __428584_428584;
   reg _428585_428585 ; 
   reg __428585_428585;
   reg _428586_428586 ; 
   reg __428586_428586;
   reg _428587_428587 ; 
   reg __428587_428587;
   reg _428588_428588 ; 
   reg __428588_428588;
   reg _428589_428589 ; 
   reg __428589_428589;
   reg _428590_428590 ; 
   reg __428590_428590;
   reg _428591_428591 ; 
   reg __428591_428591;
   reg _428592_428592 ; 
   reg __428592_428592;
   reg _428593_428593 ; 
   reg __428593_428593;
   reg _428594_428594 ; 
   reg __428594_428594;
   reg _428595_428595 ; 
   reg __428595_428595;
   reg _428596_428596 ; 
   reg __428596_428596;
   reg _428597_428597 ; 
   reg __428597_428597;
   reg _428598_428598 ; 
   reg __428598_428598;
   reg _428599_428599 ; 
   reg __428599_428599;
   reg _428600_428600 ; 
   reg __428600_428600;
   reg _428601_428601 ; 
   reg __428601_428601;
   reg _428602_428602 ; 
   reg __428602_428602;
   reg _428603_428603 ; 
   reg __428603_428603;
   reg _428604_428604 ; 
   reg __428604_428604;
   reg _428605_428605 ; 
   reg __428605_428605;
   reg _428606_428606 ; 
   reg __428606_428606;
   reg _428607_428607 ; 
   reg __428607_428607;
   reg _428608_428608 ; 
   reg __428608_428608;
   reg _428609_428609 ; 
   reg __428609_428609;
   reg _428610_428610 ; 
   reg __428610_428610;
   reg _428611_428611 ; 
   reg __428611_428611;
   reg _428612_428612 ; 
   reg __428612_428612;
   reg _428613_428613 ; 
   reg __428613_428613;
   reg _428614_428614 ; 
   reg __428614_428614;
   reg _428615_428615 ; 
   reg __428615_428615;
   reg _428616_428616 ; 
   reg __428616_428616;
   reg _428617_428617 ; 
   reg __428617_428617;
   reg _428618_428618 ; 
   reg __428618_428618;
   reg _428619_428619 ; 
   reg __428619_428619;
   reg _428620_428620 ; 
   reg __428620_428620;
   reg _428621_428621 ; 
   reg __428621_428621;
   reg _428622_428622 ; 
   reg __428622_428622;
   reg _428623_428623 ; 
   reg __428623_428623;
   reg _428624_428624 ; 
   reg __428624_428624;
   reg _428625_428625 ; 
   reg __428625_428625;
   reg _428626_428626 ; 
   reg __428626_428626;
   reg _428627_428627 ; 
   reg __428627_428627;
   reg _428628_428628 ; 
   reg __428628_428628;
   reg _428629_428629 ; 
   reg __428629_428629;
   reg _428630_428630 ; 
   reg __428630_428630;
   reg _428631_428631 ; 
   reg __428631_428631;
   reg _428632_428632 ; 
   reg __428632_428632;
   reg _428633_428633 ; 
   reg __428633_428633;
   reg _428634_428634 ; 
   reg __428634_428634;
   reg _428635_428635 ; 
   reg __428635_428635;
   reg _428636_428636 ; 
   reg __428636_428636;
   reg _428637_428637 ; 
   reg __428637_428637;
   reg _428638_428638 ; 
   reg __428638_428638;
   reg _428639_428639 ; 
   reg __428639_428639;
   reg _428640_428640 ; 
   reg __428640_428640;
   reg _428641_428641 ; 
   reg __428641_428641;
   reg _428642_428642 ; 
   reg __428642_428642;
   reg _428643_428643 ; 
   reg __428643_428643;
   reg _428644_428644 ; 
   reg __428644_428644;
   reg _428645_428645 ; 
   reg __428645_428645;
   reg _428646_428646 ; 
   reg __428646_428646;
   reg _428647_428647 ; 
   reg __428647_428647;
   reg _428648_428648 ; 
   reg __428648_428648;
   reg _428649_428649 ; 
   reg __428649_428649;
   reg _428650_428650 ; 
   reg __428650_428650;
   reg _428651_428651 ; 
   reg __428651_428651;
   reg _428652_428652 ; 
   reg __428652_428652;
   reg _428653_428653 ; 
   reg __428653_428653;
   reg _428654_428654 ; 
   reg __428654_428654;
   reg _428655_428655 ; 
   reg __428655_428655;
   reg _428656_428656 ; 
   reg __428656_428656;
   reg _428657_428657 ; 
   reg __428657_428657;
   reg _428658_428658 ; 
   reg __428658_428658;
   reg _428659_428659 ; 
   reg __428659_428659;
   reg _428660_428660 ; 
   reg __428660_428660;
   reg _428661_428661 ; 
   reg __428661_428661;
   reg _428662_428662 ; 
   reg __428662_428662;
   reg _428663_428663 ; 
   reg __428663_428663;
   reg _428664_428664 ; 
   reg __428664_428664;
   reg _428665_428665 ; 
   reg __428665_428665;
   reg _428666_428666 ; 
   reg __428666_428666;
   reg _428667_428667 ; 
   reg __428667_428667;
   reg _428668_428668 ; 
   reg __428668_428668;
   reg _428669_428669 ; 
   reg __428669_428669;
   reg _428670_428670 ; 
   reg __428670_428670;
   reg _428671_428671 ; 
   reg __428671_428671;
   reg _428672_428672 ; 
   reg __428672_428672;
   reg _428673_428673 ; 
   reg __428673_428673;
   reg _428674_428674 ; 
   reg __428674_428674;
   reg _428675_428675 ; 
   reg __428675_428675;
   reg _428676_428676 ; 
   reg __428676_428676;
   reg _428677_428677 ; 
   reg __428677_428677;
   reg _428678_428678 ; 
   reg __428678_428678;
   reg _428679_428679 ; 
   reg __428679_428679;
   reg _428680_428680 ; 
   reg __428680_428680;
   reg _428681_428681 ; 
   reg __428681_428681;
   reg _428682_428682 ; 
   reg __428682_428682;
   reg _428683_428683 ; 
   reg __428683_428683;
   reg _428684_428684 ; 
   reg __428684_428684;
   reg _428685_428685 ; 
   reg __428685_428685;
   reg _428686_428686 ; 
   reg __428686_428686;
   reg _428687_428687 ; 
   reg __428687_428687;
   reg _428688_428688 ; 
   reg __428688_428688;
   reg _428689_428689 ; 
   reg __428689_428689;
   reg _428690_428690 ; 
   reg __428690_428690;
   reg _428691_428691 ; 
   reg __428691_428691;
   reg _428692_428692 ; 
   reg __428692_428692;
   reg _428693_428693 ; 
   reg __428693_428693;
   reg _428694_428694 ; 
   reg __428694_428694;
   reg _428695_428695 ; 
   reg __428695_428695;
   reg _428696_428696 ; 
   reg __428696_428696;
   reg _428697_428697 ; 
   reg __428697_428697;
   reg _428698_428698 ; 
   reg __428698_428698;
   reg _428699_428699 ; 
   reg __428699_428699;
   reg _428700_428700 ; 
   reg __428700_428700;
   reg _428701_428701 ; 
   reg __428701_428701;
   reg _428702_428702 ; 
   reg __428702_428702;
   reg _428703_428703 ; 
   reg __428703_428703;
   reg _428704_428704 ; 
   reg __428704_428704;
   reg _428705_428705 ; 
   reg __428705_428705;
   reg _428706_428706 ; 
   reg __428706_428706;
   reg _428707_428707 ; 
   reg __428707_428707;
   reg _428708_428708 ; 
   reg __428708_428708;
   reg _428709_428709 ; 
   reg __428709_428709;
   reg _428710_428710 ; 
   reg __428710_428710;
   reg _428711_428711 ; 
   reg __428711_428711;
   reg _428712_428712 ; 
   reg __428712_428712;
   reg _428713_428713 ; 
   reg __428713_428713;
   reg _428714_428714 ; 
   reg __428714_428714;
   reg _428715_428715 ; 
   reg __428715_428715;
   reg _428716_428716 ; 
   reg __428716_428716;
   reg _428717_428717 ; 
   reg __428717_428717;
   reg _428718_428718 ; 
   reg __428718_428718;
   reg _428719_428719 ; 
   reg __428719_428719;
   reg _428720_428720 ; 
   reg __428720_428720;
   reg _428721_428721 ; 
   reg __428721_428721;
   reg _428722_428722 ; 
   reg __428722_428722;
   reg _428723_428723 ; 
   reg __428723_428723;
   reg _428724_428724 ; 
   reg __428724_428724;
   reg _428725_428725 ; 
   reg __428725_428725;
   reg _428726_428726 ; 
   reg __428726_428726;
   reg _428727_428727 ; 
   reg __428727_428727;
   reg _428728_428728 ; 
   reg __428728_428728;
   reg _428729_428729 ; 
   reg __428729_428729;
   reg _428730_428730 ; 
   reg __428730_428730;
   reg _428731_428731 ; 
   reg __428731_428731;
   reg _428732_428732 ; 
   reg __428732_428732;
   reg _428733_428733 ; 
   reg __428733_428733;
   reg _428734_428734 ; 
   reg __428734_428734;
   reg _428735_428735 ; 
   reg __428735_428735;
   reg _428736_428736 ; 
   reg __428736_428736;
   reg _428737_428737 ; 
   reg __428737_428737;
   reg _428738_428738 ; 
   reg __428738_428738;
   reg _428739_428739 ; 
   reg __428739_428739;
   reg _428740_428740 ; 
   reg __428740_428740;
   reg _428741_428741 ; 
   reg __428741_428741;
   reg _428742_428742 ; 
   reg __428742_428742;
   reg _428743_428743 ; 
   reg __428743_428743;
   reg _428744_428744 ; 
   reg __428744_428744;
   reg _428745_428745 ; 
   reg __428745_428745;
   reg _428746_428746 ; 
   reg __428746_428746;
   reg _428747_428747 ; 
   reg __428747_428747;
   reg _428748_428748 ; 
   reg __428748_428748;
   reg _428749_428749 ; 
   reg __428749_428749;
   reg _428750_428750 ; 
   reg __428750_428750;
   reg _428751_428751 ; 
   reg __428751_428751;
   reg _428752_428752 ; 
   reg __428752_428752;
   reg _428753_428753 ; 
   reg __428753_428753;
   reg _428754_428754 ; 
   reg __428754_428754;
   reg _428755_428755 ; 
   reg __428755_428755;
   reg _428756_428756 ; 
   reg __428756_428756;
   reg _428757_428757 ; 
   reg __428757_428757;
   reg _428758_428758 ; 
   reg __428758_428758;
   reg _428759_428759 ; 
   reg __428759_428759;
   reg _428760_428760 ; 
   reg __428760_428760;
   reg _428761_428761 ; 
   reg __428761_428761;
   reg _428762_428762 ; 
   reg __428762_428762;
   reg _428763_428763 ; 
   reg __428763_428763;
   reg _428764_428764 ; 
   reg __428764_428764;
   reg _428765_428765 ; 
   reg __428765_428765;
   reg _428766_428766 ; 
   reg __428766_428766;
   reg _428767_428767 ; 
   reg __428767_428767;
   reg _428768_428768 ; 
   reg __428768_428768;
   reg _428769_428769 ; 
   reg __428769_428769;
   reg _428770_428770 ; 
   reg __428770_428770;
   reg _428771_428771 ; 
   reg __428771_428771;
   reg _428772_428772 ; 
   reg __428772_428772;
   reg _428773_428773 ; 
   reg __428773_428773;
   reg _428774_428774 ; 
   reg __428774_428774;
   reg _428775_428775 ; 
   reg __428775_428775;
   reg _428776_428776 ; 
   reg __428776_428776;
   reg _428777_428777 ; 
   reg __428777_428777;
   reg _428778_428778 ; 
   reg __428778_428778;
   reg _428779_428779 ; 
   reg __428779_428779;
   reg _428780_428780 ; 
   reg __428780_428780;
   reg _428781_428781 ; 
   reg __428781_428781;
   reg _428782_428782 ; 
   reg __428782_428782;
   reg _428783_428783 ; 
   reg __428783_428783;
   reg _428784_428784 ; 
   reg __428784_428784;
   reg _428785_428785 ; 
   reg __428785_428785;
   reg _428786_428786 ; 
   reg __428786_428786;
   reg _428787_428787 ; 
   reg __428787_428787;
   reg _428788_428788 ; 
   reg __428788_428788;
   reg _428789_428789 ; 
   reg __428789_428789;
   reg _428790_428790 ; 
   reg __428790_428790;
   reg _428791_428791 ; 
   reg __428791_428791;
   reg _428792_428792 ; 
   reg __428792_428792;
   reg _428793_428793 ; 
   reg __428793_428793;
   reg _428794_428794 ; 
   reg __428794_428794;
   reg _428795_428795 ; 
   reg __428795_428795;
   reg _428796_428796 ; 
   reg __428796_428796;
   reg _428797_428797 ; 
   reg __428797_428797;
   reg _428798_428798 ; 
   reg __428798_428798;
   reg _428799_428799 ; 
   reg __428799_428799;
   reg _428800_428800 ; 
   reg __428800_428800;
   reg _428801_428801 ; 
   reg __428801_428801;
   reg _428802_428802 ; 
   reg __428802_428802;
   reg _428803_428803 ; 
   reg __428803_428803;
   reg _428804_428804 ; 
   reg __428804_428804;
   reg _428805_428805 ; 
   reg __428805_428805;
   reg _428806_428806 ; 
   reg __428806_428806;
   reg _428807_428807 ; 
   reg __428807_428807;
   reg _428808_428808 ; 
   reg __428808_428808;
   reg _428809_428809 ; 
   reg __428809_428809;
   reg _428810_428810 ; 
   reg __428810_428810;
   reg _428811_428811 ; 
   reg __428811_428811;
   reg _428812_428812 ; 
   reg __428812_428812;
   reg _428813_428813 ; 
   reg __428813_428813;
   reg _428814_428814 ; 
   reg __428814_428814;
   reg _428815_428815 ; 
   reg __428815_428815;
   reg _428816_428816 ; 
   reg __428816_428816;
   reg _428817_428817 ; 
   reg __428817_428817;
   reg _428818_428818 ; 
   reg __428818_428818;
   reg _428819_428819 ; 
   reg __428819_428819;
   reg _428820_428820 ; 
   reg __428820_428820;
   reg _428821_428821 ; 
   reg __428821_428821;
   reg _428822_428822 ; 
   reg __428822_428822;
   reg _428823_428823 ; 
   reg __428823_428823;
   reg _428824_428824 ; 
   reg __428824_428824;
   reg _428825_428825 ; 
   reg __428825_428825;
   reg _428826_428826 ; 
   reg __428826_428826;
   reg _428827_428827 ; 
   reg __428827_428827;
   reg _428828_428828 ; 
   reg __428828_428828;
   reg _428829_428829 ; 
   reg __428829_428829;
   reg _428830_428830 ; 
   reg __428830_428830;
   reg _428831_428831 ; 
   reg __428831_428831;
   reg _428832_428832 ; 
   reg __428832_428832;
   reg _428833_428833 ; 
   reg __428833_428833;
   reg _428834_428834 ; 
   reg __428834_428834;
   reg _428835_428835 ; 
   reg __428835_428835;
   reg _428836_428836 ; 
   reg __428836_428836;
   reg _428837_428837 ; 
   reg __428837_428837;
   reg _428838_428838 ; 
   reg __428838_428838;
   reg _428839_428839 ; 
   reg __428839_428839;
   reg _428840_428840 ; 
   reg __428840_428840;
   reg _428841_428841 ; 
   reg __428841_428841;
   reg _428842_428842 ; 
   reg __428842_428842;
   reg _428843_428843 ; 
   reg __428843_428843;
   reg _428844_428844 ; 
   reg __428844_428844;
   reg _428845_428845 ; 
   reg __428845_428845;
   reg _428846_428846 ; 
   reg __428846_428846;
   reg _428847_428847 ; 
   reg __428847_428847;
   reg _428848_428848 ; 
   reg __428848_428848;
   reg _428849_428849 ; 
   reg __428849_428849;
   reg _428850_428850 ; 
   reg __428850_428850;
   reg _428851_428851 ; 
   reg __428851_428851;
   reg _428852_428852 ; 
   reg __428852_428852;
   reg _428853_428853 ; 
   reg __428853_428853;
   reg _428854_428854 ; 
   reg __428854_428854;
   reg _428855_428855 ; 
   reg __428855_428855;
   reg _428856_428856 ; 
   reg __428856_428856;
   reg _428857_428857 ; 
   reg __428857_428857;
   reg _428858_428858 ; 
   reg __428858_428858;
   reg _428859_428859 ; 
   reg __428859_428859;
   reg _428860_428860 ; 
   reg __428860_428860;
   reg _428861_428861 ; 
   reg __428861_428861;
   reg _428862_428862 ; 
   reg __428862_428862;
   reg _428863_428863 ; 
   reg __428863_428863;
   reg _428864_428864 ; 
   reg __428864_428864;
   reg _428865_428865 ; 
   reg __428865_428865;
   reg _428866_428866 ; 
   reg __428866_428866;
   reg _428867_428867 ; 
   reg __428867_428867;
   reg _428868_428868 ; 
   reg __428868_428868;
   reg _428869_428869 ; 
   reg __428869_428869;
   reg _428870_428870 ; 
   reg __428870_428870;
   reg _428871_428871 ; 
   reg __428871_428871;
   reg _428872_428872 ; 
   reg __428872_428872;
   reg _428873_428873 ; 
   reg __428873_428873;
   reg _428874_428874 ; 
   reg __428874_428874;
   reg _428875_428875 ; 
   reg __428875_428875;
   reg _428876_428876 ; 
   reg __428876_428876;
   reg _428877_428877 ; 
   reg __428877_428877;
   reg _428878_428878 ; 
   reg __428878_428878;
   reg _428879_428879 ; 
   reg __428879_428879;
   reg _428880_428880 ; 
   reg __428880_428880;
   reg _428881_428881 ; 
   reg __428881_428881;
   reg _428882_428882 ; 
   reg __428882_428882;
   reg _428883_428883 ; 
   reg __428883_428883;
   reg _428884_428884 ; 
   reg __428884_428884;
   reg _428885_428885 ; 
   reg __428885_428885;
   reg _428886_428886 ; 
   reg __428886_428886;
   reg _428887_428887 ; 
   reg __428887_428887;
   reg _428888_428888 ; 
   reg __428888_428888;
   reg _428889_428889 ; 
   reg __428889_428889;
   reg _428890_428890 ; 
   reg __428890_428890;
   reg _428891_428891 ; 
   reg __428891_428891;
   reg _428892_428892 ; 
   reg __428892_428892;
   reg _428893_428893 ; 
   reg __428893_428893;
   reg _428894_428894 ; 
   reg __428894_428894;
   reg _428895_428895 ; 
   reg __428895_428895;
   reg _428896_428896 ; 
   reg __428896_428896;
   reg _428897_428897 ; 
   reg __428897_428897;
   reg _428898_428898 ; 
   reg __428898_428898;
   reg _428899_428899 ; 
   reg __428899_428899;
   reg _428900_428900 ; 
   reg __428900_428900;
   reg _428901_428901 ; 
   reg __428901_428901;
   reg _428902_428902 ; 
   reg __428902_428902;
   reg _428903_428903 ; 
   reg __428903_428903;
   reg _428904_428904 ; 
   reg __428904_428904;
   reg _428905_428905 ; 
   reg __428905_428905;
   reg _428906_428906 ; 
   reg __428906_428906;
   reg _428907_428907 ; 
   reg __428907_428907;
   reg _428908_428908 ; 
   reg __428908_428908;
   reg _428909_428909 ; 
   reg __428909_428909;
   reg _428910_428910 ; 
   reg __428910_428910;
   reg _428911_428911 ; 
   reg __428911_428911;
   reg _428912_428912 ; 
   reg __428912_428912;
   reg _428913_428913 ; 
   reg __428913_428913;
   reg _428914_428914 ; 
   reg __428914_428914;
   reg _428915_428915 ; 
   reg __428915_428915;
   reg _428916_428916 ; 
   reg __428916_428916;
   reg _428917_428917 ; 
   reg __428917_428917;
   reg _428918_428918 ; 
   reg __428918_428918;
   reg _428919_428919 ; 
   reg __428919_428919;
   reg _428920_428920 ; 
   reg __428920_428920;
   reg _428921_428921 ; 
   reg __428921_428921;
   reg _428922_428922 ; 
   reg __428922_428922;
   reg _428923_428923 ; 
   reg __428923_428923;
   reg _428924_428924 ; 
   reg __428924_428924;
   reg _428925_428925 ; 
   reg __428925_428925;
   reg _428926_428926 ; 
   reg __428926_428926;
   reg _428927_428927 ; 
   reg __428927_428927;
   reg _428928_428928 ; 
   reg __428928_428928;
   reg _428929_428929 ; 
   reg __428929_428929;
   reg _428930_428930 ; 
   reg __428930_428930;
   reg _428931_428931 ; 
   reg __428931_428931;
   reg _428932_428932 ; 
   reg __428932_428932;
   reg _428933_428933 ; 
   reg __428933_428933;
   reg _428934_428934 ; 
   reg __428934_428934;
   reg _428935_428935 ; 
   reg __428935_428935;
   reg _428936_428936 ; 
   reg __428936_428936;
   reg _428937_428937 ; 
   reg __428937_428937;
   reg _428938_428938 ; 
   reg __428938_428938;
   reg _428939_428939 ; 
   reg __428939_428939;
   reg _428940_428940 ; 
   reg __428940_428940;
   reg _428941_428941 ; 
   reg __428941_428941;
   reg _428942_428942 ; 
   reg __428942_428942;
   reg _428943_428943 ; 
   reg __428943_428943;
   reg _428944_428944 ; 
   reg __428944_428944;
   reg _428945_428945 ; 
   reg __428945_428945;
   reg _428946_428946 ; 
   reg __428946_428946;
   reg _428947_428947 ; 
   reg __428947_428947;
   reg _428948_428948 ; 
   reg __428948_428948;
   reg _428949_428949 ; 
   reg __428949_428949;
   reg _428950_428950 ; 
   reg __428950_428950;
   reg _428951_428951 ; 
   reg __428951_428951;
   reg _428952_428952 ; 
   reg __428952_428952;
   reg _428953_428953 ; 
   reg __428953_428953;
   reg _428954_428954 ; 
   reg __428954_428954;
   reg _428955_428955 ; 
   reg __428955_428955;
   reg _428956_428956 ; 
   reg __428956_428956;
   reg _428957_428957 ; 
   reg __428957_428957;
   reg _428958_428958 ; 
   reg __428958_428958;
   reg _428959_428959 ; 
   reg __428959_428959;
   reg _428960_428960 ; 
   reg __428960_428960;
   reg _428961_428961 ; 
   reg __428961_428961;
   reg _428962_428962 ; 
   reg __428962_428962;
   reg _428963_428963 ; 
   reg __428963_428963;
   reg _428964_428964 ; 
   reg __428964_428964;
   reg _428965_428965 ; 
   reg __428965_428965;
   reg _428966_428966 ; 
   reg __428966_428966;
   reg _428967_428967 ; 
   reg __428967_428967;
   reg _428968_428968 ; 
   reg __428968_428968;
   reg _428969_428969 ; 
   reg __428969_428969;
   reg _428970_428970 ; 
   reg __428970_428970;
   reg _428971_428971 ; 
   reg __428971_428971;
   reg _428972_428972 ; 
   reg __428972_428972;
   reg _428973_428973 ; 
   reg __428973_428973;
   reg _428974_428974 ; 
   reg __428974_428974;
   reg _428975_428975 ; 
   reg __428975_428975;
   reg _428976_428976 ; 
   reg __428976_428976;
   reg _428977_428977 ; 
   reg __428977_428977;
   reg _428978_428978 ; 
   reg __428978_428978;
   reg _428979_428979 ; 
   reg __428979_428979;
   reg _428980_428980 ; 
   reg __428980_428980;
   reg _428981_428981 ; 
   reg __428981_428981;
   reg _428982_428982 ; 
   reg __428982_428982;
   reg _428983_428983 ; 
   reg __428983_428983;
   reg _428984_428984 ; 
   reg __428984_428984;
   reg _428985_428985 ; 
   reg __428985_428985;
   reg _428986_428986 ; 
   reg __428986_428986;
   reg _428987_428987 ; 
   reg __428987_428987;
   reg _428988_428988 ; 
   reg __428988_428988;
   reg _428989_428989 ; 
   reg __428989_428989;
   reg _428990_428990 ; 
   reg __428990_428990;
   reg _428991_428991 ; 
   reg __428991_428991;
   reg _428992_428992 ; 
   reg __428992_428992;
   reg _428993_428993 ; 
   reg __428993_428993;
   reg _428994_428994 ; 
   reg __428994_428994;
   reg _428995_428995 ; 
   reg __428995_428995;
   reg _428996_428996 ; 
   reg __428996_428996;
   reg _428997_428997 ; 
   reg __428997_428997;
   reg _428998_428998 ; 
   reg __428998_428998;
   reg _428999_428999 ; 
   reg __428999_428999;
   reg _429000_429000 ; 
   reg __429000_429000;
   reg _429001_429001 ; 
   reg __429001_429001;
   reg _429002_429002 ; 
   reg __429002_429002;
   reg _429003_429003 ; 
   reg __429003_429003;
   reg _429004_429004 ; 
   reg __429004_429004;
   reg _429005_429005 ; 
   reg __429005_429005;
   reg _429006_429006 ; 
   reg __429006_429006;
   reg _429007_429007 ; 
   reg __429007_429007;
   reg _429008_429008 ; 
   reg __429008_429008;
   reg _429009_429009 ; 
   reg __429009_429009;
   reg _429010_429010 ; 
   reg __429010_429010;
   reg _429011_429011 ; 
   reg __429011_429011;
   reg _429012_429012 ; 
   reg __429012_429012;
   reg _429013_429013 ; 
   reg __429013_429013;
   reg _429014_429014 ; 
   reg __429014_429014;
   reg _429015_429015 ; 
   reg __429015_429015;
   reg _429016_429016 ; 
   reg __429016_429016;
   reg _429017_429017 ; 
   reg __429017_429017;
   reg _429018_429018 ; 
   reg __429018_429018;
   reg _429019_429019 ; 
   reg __429019_429019;
   reg _429020_429020 ; 
   reg __429020_429020;
   reg _429021_429021 ; 
   reg __429021_429021;
   reg _429022_429022 ; 
   reg __429022_429022;
   reg _429023_429023 ; 
   reg __429023_429023;
   reg _429024_429024 ; 
   reg __429024_429024;
   reg _429025_429025 ; 
   reg __429025_429025;
   reg _429026_429026 ; 
   reg __429026_429026;
   reg _429027_429027 ; 
   reg __429027_429027;
   reg _429028_429028 ; 
   reg __429028_429028;
   reg _429029_429029 ; 
   reg __429029_429029;
   reg _429030_429030 ; 
   reg __429030_429030;
   reg _429031_429031 ; 
   reg __429031_429031;
   reg _429032_429032 ; 
   reg __429032_429032;
   reg _429033_429033 ; 
   reg __429033_429033;
   reg _429034_429034 ; 
   reg __429034_429034;
   reg _429035_429035 ; 
   reg __429035_429035;
   reg _429036_429036 ; 
   reg __429036_429036;
   reg _429037_429037 ; 
   reg __429037_429037;
   reg _429038_429038 ; 
   reg __429038_429038;
   reg _429039_429039 ; 
   reg __429039_429039;
   reg _429040_429040 ; 
   reg __429040_429040;
   reg _429041_429041 ; 
   reg __429041_429041;
   reg _429042_429042 ; 
   reg __429042_429042;
   reg _429043_429043 ; 
   reg __429043_429043;
   reg _429044_429044 ; 
   reg __429044_429044;
   reg _429045_429045 ; 
   reg __429045_429045;
   reg _429046_429046 ; 
   reg __429046_429046;
   reg _429047_429047 ; 
   reg __429047_429047;
   reg _429048_429048 ; 
   reg __429048_429048;
   reg _429049_429049 ; 
   reg __429049_429049;
   reg _429050_429050 ; 
   reg __429050_429050;
   reg _429051_429051 ; 
   reg __429051_429051;
   reg _429052_429052 ; 
   reg __429052_429052;
   reg _429053_429053 ; 
   reg __429053_429053;
   reg _429054_429054 ; 
   reg __429054_429054;
   reg _429055_429055 ; 
   reg __429055_429055;
   reg _429056_429056 ; 
   reg __429056_429056;
   reg _429057_429057 ; 
   reg __429057_429057;
   reg _429058_429058 ; 
   reg __429058_429058;
   reg _429059_429059 ; 
   reg __429059_429059;
   reg _429060_429060 ; 
   reg __429060_429060;
   reg _429061_429061 ; 
   reg __429061_429061;
   reg _429062_429062 ; 
   reg __429062_429062;
   reg _429063_429063 ; 
   reg __429063_429063;
   reg _429064_429064 ; 
   reg __429064_429064;
   reg _429065_429065 ; 
   reg __429065_429065;
   reg _429066_429066 ; 
   reg __429066_429066;
   reg _429067_429067 ; 
   reg __429067_429067;
   reg _429068_429068 ; 
   reg __429068_429068;
   reg _429069_429069 ; 
   reg __429069_429069;
   reg _429070_429070 ; 
   reg __429070_429070;
   reg _429071_429071 ; 
   reg __429071_429071;
   reg _429072_429072 ; 
   reg __429072_429072;
   reg _429073_429073 ; 
   reg __429073_429073;
   reg _429074_429074 ; 
   reg __429074_429074;
   reg _429075_429075 ; 
   reg __429075_429075;
   reg _429076_429076 ; 
   reg __429076_429076;
   reg _429077_429077 ; 
   reg __429077_429077;
   reg _429078_429078 ; 
   reg __429078_429078;
   reg _429079_429079 ; 
   reg __429079_429079;
   reg _429080_429080 ; 
   reg __429080_429080;
   reg _429081_429081 ; 
   reg __429081_429081;
   reg _429082_429082 ; 
   reg __429082_429082;
   reg _429083_429083 ; 
   reg __429083_429083;
   reg _429084_429084 ; 
   reg __429084_429084;
   reg _429085_429085 ; 
   reg __429085_429085;
   reg _429086_429086 ; 
   reg __429086_429086;
   reg _429087_429087 ; 
   reg __429087_429087;
   reg _429088_429088 ; 
   reg __429088_429088;
   reg _429089_429089 ; 
   reg __429089_429089;
   reg _429090_429090 ; 
   reg __429090_429090;
   reg _429091_429091 ; 
   reg __429091_429091;
   reg _429092_429092 ; 
   reg __429092_429092;
   reg _429093_429093 ; 
   reg __429093_429093;
   reg _429094_429094 ; 
   reg __429094_429094;
   reg _429095_429095 ; 
   reg __429095_429095;
   reg _429096_429096 ; 
   reg __429096_429096;
   reg _429097_429097 ; 
   reg __429097_429097;
   reg _429098_429098 ; 
   reg __429098_429098;
   reg _429099_429099 ; 
   reg __429099_429099;
   reg _429100_429100 ; 
   reg __429100_429100;
   reg _429101_429101 ; 
   reg __429101_429101;
   reg _429102_429102 ; 
   reg __429102_429102;
   reg _429103_429103 ; 
   reg __429103_429103;
   reg _429104_429104 ; 
   reg __429104_429104;
   reg _429105_429105 ; 
   reg __429105_429105;
   reg _429106_429106 ; 
   reg __429106_429106;
   reg _429107_429107 ; 
   reg __429107_429107;
   reg _429108_429108 ; 
   reg __429108_429108;
   reg _429109_429109 ; 
   reg __429109_429109;
   reg _429110_429110 ; 
   reg __429110_429110;
   reg _429111_429111 ; 
   reg __429111_429111;
   reg _429112_429112 ; 
   reg __429112_429112;
   reg _429113_429113 ; 
   reg __429113_429113;
   reg _429114_429114 ; 
   reg __429114_429114;
   reg _429115_429115 ; 
   reg __429115_429115;
   reg _429116_429116 ; 
   reg __429116_429116;
   reg _429117_429117 ; 
   reg __429117_429117;
   reg _429118_429118 ; 
   reg __429118_429118;
   reg _429119_429119 ; 
   reg __429119_429119;
   reg _429120_429120 ; 
   reg __429120_429120;
   reg _429121_429121 ; 
   reg __429121_429121;
   reg _429122_429122 ; 
   reg __429122_429122;
   reg _429123_429123 ; 
   reg __429123_429123;
   reg _429124_429124 ; 
   reg __429124_429124;
   reg _429125_429125 ; 
   reg __429125_429125;
   reg _429126_429126 ; 
   reg __429126_429126;
   reg _429127_429127 ; 
   reg __429127_429127;
   reg _429128_429128 ; 
   reg __429128_429128;
   reg _429129_429129 ; 
   reg __429129_429129;
   reg _429130_429130 ; 
   reg __429130_429130;
   reg _429131_429131 ; 
   reg __429131_429131;
   reg _429132_429132 ; 
   reg __429132_429132;
   reg _429133_429133 ; 
   reg __429133_429133;
   reg _429134_429134 ; 
   reg __429134_429134;
   reg _429135_429135 ; 
   reg __429135_429135;
   reg _429136_429136 ; 
   reg __429136_429136;
   reg _429137_429137 ; 
   reg __429137_429137;
   reg _429138_429138 ; 
   reg __429138_429138;
   reg _429139_429139 ; 
   reg __429139_429139;
   reg _429140_429140 ; 
   reg __429140_429140;
   reg _429141_429141 ; 
   reg __429141_429141;
   reg _429142_429142 ; 
   reg __429142_429142;
   reg _429143_429143 ; 
   reg __429143_429143;
   reg _429144_429144 ; 
   reg __429144_429144;
   reg _429145_429145 ; 
   reg __429145_429145;
   reg _429146_429146 ; 
   reg __429146_429146;
   reg _429147_429147 ; 
   reg __429147_429147;
   reg _429148_429148 ; 
   reg __429148_429148;
   reg _429149_429149 ; 
   reg __429149_429149;
   reg _429150_429150 ; 
   reg __429150_429150;
   reg _429151_429151 ; 
   reg __429151_429151;
   reg _429152_429152 ; 
   reg __429152_429152;
   reg _429153_429153 ; 
   reg __429153_429153;
   reg _429154_429154 ; 
   reg __429154_429154;
   reg _429155_429155 ; 
   reg __429155_429155;
   reg _429156_429156 ; 
   reg __429156_429156;
   reg _429157_429157 ; 
   reg __429157_429157;
   reg _429158_429158 ; 
   reg __429158_429158;
   reg _429159_429159 ; 
   reg __429159_429159;
   reg _429160_429160 ; 
   reg __429160_429160;
   reg _429161_429161 ; 
   reg __429161_429161;
   reg _429162_429162 ; 
   reg __429162_429162;
   reg _429163_429163 ; 
   reg __429163_429163;
   reg _429164_429164 ; 
   reg __429164_429164;
   reg _429165_429165 ; 
   reg __429165_429165;
   reg _429166_429166 ; 
   reg __429166_429166;
   reg _429167_429167 ; 
   reg __429167_429167;
   reg _429168_429168 ; 
   reg __429168_429168;
   reg _429169_429169 ; 
   reg __429169_429169;
   reg _429170_429170 ; 
   reg __429170_429170;
   reg _429171_429171 ; 
   reg __429171_429171;
   reg _429172_429172 ; 
   reg __429172_429172;
   reg _429173_429173 ; 
   reg __429173_429173;
   reg _429174_429174 ; 
   reg __429174_429174;
   reg _429175_429175 ; 
   reg __429175_429175;
   reg _429176_429176 ; 
   reg __429176_429176;
   reg _429177_429177 ; 
   reg __429177_429177;
   reg _429178_429178 ; 
   reg __429178_429178;
   reg _429179_429179 ; 
   reg __429179_429179;
   reg _429180_429180 ; 
   reg __429180_429180;
   reg _429181_429181 ; 
   reg __429181_429181;
   reg _429182_429182 ; 
   reg __429182_429182;
   reg _429183_429183 ; 
   reg __429183_429183;
   reg _429184_429184 ; 
   reg __429184_429184;
   reg _429185_429185 ; 
   reg __429185_429185;
   reg _429186_429186 ; 
   reg __429186_429186;
   reg _429187_429187 ; 
   reg __429187_429187;
   reg _429188_429188 ; 
   reg __429188_429188;
   reg _429189_429189 ; 
   reg __429189_429189;
   reg _429190_429190 ; 
   reg __429190_429190;
   reg _429191_429191 ; 
   reg __429191_429191;
   reg _429192_429192 ; 
   reg __429192_429192;
   reg _429193_429193 ; 
   reg __429193_429193;
   reg _429194_429194 ; 
   reg __429194_429194;
   reg _429195_429195 ; 
   reg __429195_429195;
   reg _429196_429196 ; 
   reg __429196_429196;
   reg _429197_429197 ; 
   reg __429197_429197;
   reg _429198_429198 ; 
   reg __429198_429198;
   reg _429199_429199 ; 
   reg __429199_429199;
   reg _429200_429200 ; 
   reg __429200_429200;
   reg _429201_429201 ; 
   reg __429201_429201;
   reg _429202_429202 ; 
   reg __429202_429202;
   reg _429203_429203 ; 
   reg __429203_429203;
   reg _429204_429204 ; 
   reg __429204_429204;
   reg _429205_429205 ; 
   reg __429205_429205;
   reg _429206_429206 ; 
   reg __429206_429206;
   reg _429207_429207 ; 
   reg __429207_429207;
   reg _429208_429208 ; 
   reg __429208_429208;
   reg _429209_429209 ; 
   reg __429209_429209;
   reg _429210_429210 ; 
   reg __429210_429210;
   reg _429211_429211 ; 
   reg __429211_429211;
   reg _429212_429212 ; 
   reg __429212_429212;
   reg _429213_429213 ; 
   reg __429213_429213;
   reg _429214_429214 ; 
   reg __429214_429214;
   reg _429215_429215 ; 
   reg __429215_429215;
   reg _429216_429216 ; 
   reg __429216_429216;
   reg _429217_429217 ; 
   reg __429217_429217;
   reg _429218_429218 ; 
   reg __429218_429218;
   reg _429219_429219 ; 
   reg __429219_429219;
   reg _429220_429220 ; 
   reg __429220_429220;
   reg _429221_429221 ; 
   reg __429221_429221;
   reg _429222_429222 ; 
   reg __429222_429222;
   reg _429223_429223 ; 
   reg __429223_429223;
   reg _429224_429224 ; 
   reg __429224_429224;
   reg _429225_429225 ; 
   reg __429225_429225;
   reg _429226_429226 ; 
   reg __429226_429226;
   reg _429227_429227 ; 
   reg __429227_429227;
   reg _429228_429228 ; 
   reg __429228_429228;
   reg _429229_429229 ; 
   reg __429229_429229;
   reg _429230_429230 ; 
   reg __429230_429230;
   reg _429231_429231 ; 
   reg __429231_429231;
   reg _429232_429232 ; 
   reg __429232_429232;
   reg _429233_429233 ; 
   reg __429233_429233;
   reg _429234_429234 ; 
   reg __429234_429234;
   reg _429235_429235 ; 
   reg __429235_429235;
   reg _429236_429236 ; 
   reg __429236_429236;
   reg _429237_429237 ; 
   reg __429237_429237;
   reg _429238_429238 ; 
   reg __429238_429238;
   reg _429239_429239 ; 
   reg __429239_429239;
   reg _429240_429240 ; 
   reg __429240_429240;
   reg _429241_429241 ; 
   reg __429241_429241;
   reg _429242_429242 ; 
   reg __429242_429242;
   reg _429243_429243 ; 
   reg __429243_429243;
   reg _429244_429244 ; 
   reg __429244_429244;
   reg _429245_429245 ; 
   reg __429245_429245;
   reg _429246_429246 ; 
   reg __429246_429246;
   reg _429247_429247 ; 
   reg __429247_429247;
   reg _429248_429248 ; 
   reg __429248_429248;
   reg _429249_429249 ; 
   reg __429249_429249;
   reg _429250_429250 ; 
   reg __429250_429250;
   reg _429251_429251 ; 
   reg __429251_429251;
   reg _429252_429252 ; 
   reg __429252_429252;
   reg _429253_429253 ; 
   reg __429253_429253;
   reg _429254_429254 ; 
   reg __429254_429254;
   reg _429255_429255 ; 
   reg __429255_429255;
   reg _429256_429256 ; 
   reg __429256_429256;
   reg _429257_429257 ; 
   reg __429257_429257;
   reg _429258_429258 ; 
   reg __429258_429258;
   reg _429259_429259 ; 
   reg __429259_429259;
   reg _429260_429260 ; 
   reg __429260_429260;
   reg _429261_429261 ; 
   reg __429261_429261;
   reg _429262_429262 ; 
   reg __429262_429262;
   reg _429263_429263 ; 
   reg __429263_429263;
   reg _429264_429264 ; 
   reg __429264_429264;
   reg _429265_429265 ; 
   reg __429265_429265;
   reg _429266_429266 ; 
   reg __429266_429266;
   reg _429267_429267 ; 
   reg __429267_429267;
   reg _429268_429268 ; 
   reg __429268_429268;
   reg _429269_429269 ; 
   reg __429269_429269;
   reg _429270_429270 ; 
   reg __429270_429270;
   reg _429271_429271 ; 
   reg __429271_429271;
   reg _429272_429272 ; 
   reg __429272_429272;
   reg _429273_429273 ; 
   reg __429273_429273;
   reg _429274_429274 ; 
   reg __429274_429274;
   reg _429275_429275 ; 
   reg __429275_429275;
   reg _429276_429276 ; 
   reg __429276_429276;
   reg _429277_429277 ; 
   reg __429277_429277;
   reg _429278_429278 ; 
   reg __429278_429278;
   reg _429279_429279 ; 
   reg __429279_429279;
   reg _429280_429280 ; 
   reg __429280_429280;
   reg _429281_429281 ; 
   reg __429281_429281;
   reg _429282_429282 ; 
   reg __429282_429282;
   reg _429283_429283 ; 
   reg __429283_429283;
   reg _429284_429284 ; 
   reg __429284_429284;
   reg _429285_429285 ; 
   reg __429285_429285;
   reg _429286_429286 ; 
   reg __429286_429286;
   reg _429287_429287 ; 
   reg __429287_429287;
   reg _429288_429288 ; 
   reg __429288_429288;
   reg _429289_429289 ; 
   reg __429289_429289;
   reg _429290_429290 ; 
   reg __429290_429290;
   reg _429291_429291 ; 
   reg __429291_429291;
   reg _429292_429292 ; 
   reg __429292_429292;
   reg _429293_429293 ; 
   reg __429293_429293;
   reg _429294_429294 ; 
   reg __429294_429294;
   reg _429295_429295 ; 
   reg __429295_429295;
   reg _429296_429296 ; 
   reg __429296_429296;
   reg _429297_429297 ; 
   reg __429297_429297;
   reg _429298_429298 ; 
   reg __429298_429298;
   reg _429299_429299 ; 
   reg __429299_429299;
   reg _429300_429300 ; 
   reg __429300_429300;
   reg _429301_429301 ; 
   reg __429301_429301;
   reg _429302_429302 ; 
   reg __429302_429302;
   reg _429303_429303 ; 
   reg __429303_429303;
   reg _429304_429304 ; 
   reg __429304_429304;
   reg _429305_429305 ; 
   reg __429305_429305;
   reg _429306_429306 ; 
   reg __429306_429306;
   reg _429307_429307 ; 
   reg __429307_429307;
   reg _429308_429308 ; 
   reg __429308_429308;
   reg _429309_429309 ; 
   reg __429309_429309;
   reg _429310_429310 ; 
   reg __429310_429310;
   reg _429311_429311 ; 
   reg __429311_429311;
   reg _429312_429312 ; 
   reg __429312_429312;
   reg _429313_429313 ; 
   reg __429313_429313;
   reg _429314_429314 ; 
   reg __429314_429314;
   reg _429315_429315 ; 
   reg __429315_429315;
   reg _429316_429316 ; 
   reg __429316_429316;
   reg _429317_429317 ; 
   reg __429317_429317;
   reg _429318_429318 ; 
   reg __429318_429318;
   reg _429319_429319 ; 
   reg __429319_429319;
   reg _429320_429320 ; 
   reg __429320_429320;
   reg _429321_429321 ; 
   reg __429321_429321;
   reg _429322_429322 ; 
   reg __429322_429322;
   reg _429323_429323 ; 
   reg __429323_429323;
   reg _429324_429324 ; 
   reg __429324_429324;
   reg _429325_429325 ; 
   reg __429325_429325;
   reg _429326_429326 ; 
   reg __429326_429326;
   reg _429327_429327 ; 
   reg __429327_429327;
   reg _429328_429328 ; 
   reg __429328_429328;
   reg _429329_429329 ; 
   reg __429329_429329;
   reg _429330_429330 ; 
   reg __429330_429330;
   reg _429331_429331 ; 
   reg __429331_429331;
   reg _429332_429332 ; 
   reg __429332_429332;
   reg _429333_429333 ; 
   reg __429333_429333;
   reg _429334_429334 ; 
   reg __429334_429334;
   reg _429335_429335 ; 
   reg __429335_429335;
   reg _429336_429336 ; 
   reg __429336_429336;
   reg _429337_429337 ; 
   reg __429337_429337;
   reg _429338_429338 ; 
   reg __429338_429338;
   reg _429339_429339 ; 
   reg __429339_429339;
   reg _429340_429340 ; 
   reg __429340_429340;
   reg _429341_429341 ; 
   reg __429341_429341;
   reg _429342_429342 ; 
   reg __429342_429342;
   reg _429343_429343 ; 
   reg __429343_429343;
   reg _429344_429344 ; 
   reg __429344_429344;
   reg _429345_429345 ; 
   reg __429345_429345;
   reg _429346_429346 ; 
   reg __429346_429346;
   reg _429347_429347 ; 
   reg __429347_429347;
   reg _429348_429348 ; 
   reg __429348_429348;
   reg _429349_429349 ; 
   reg __429349_429349;
   reg _429350_429350 ; 
   reg __429350_429350;
   reg _429351_429351 ; 
   reg __429351_429351;
   reg _429352_429352 ; 
   reg __429352_429352;
   reg _429353_429353 ; 
   reg __429353_429353;
   reg _429354_429354 ; 
   reg __429354_429354;
   reg _429355_429355 ; 
   reg __429355_429355;
   reg _429356_429356 ; 
   reg __429356_429356;
   reg _429357_429357 ; 
   reg __429357_429357;
   reg _429358_429358 ; 
   reg __429358_429358;
   reg _429359_429359 ; 
   reg __429359_429359;
   reg _429360_429360 ; 
   reg __429360_429360;
   reg _429361_429361 ; 
   reg __429361_429361;
   reg _429362_429362 ; 
   reg __429362_429362;
   reg _429363_429363 ; 
   reg __429363_429363;
   reg _429364_429364 ; 
   reg __429364_429364;
   reg _429365_429365 ; 
   reg __429365_429365;
   reg _429366_429366 ; 
   reg __429366_429366;
   reg _429367_429367 ; 
   reg __429367_429367;
   reg _429368_429368 ; 
   reg __429368_429368;
   reg _429369_429369 ; 
   reg __429369_429369;
   reg _429370_429370 ; 
   reg __429370_429370;
   reg _429371_429371 ; 
   reg __429371_429371;
   reg _429372_429372 ; 
   reg __429372_429372;
   reg _429373_429373 ; 
   reg __429373_429373;
   reg _429374_429374 ; 
   reg __429374_429374;
   reg _429375_429375 ; 
   reg __429375_429375;
   reg _429376_429376 ; 
   reg __429376_429376;
   reg _429377_429377 ; 
   reg __429377_429377;
   reg _429378_429378 ; 
   reg __429378_429378;
   reg _429379_429379 ; 
   reg __429379_429379;
   reg _429380_429380 ; 
   reg __429380_429380;
   reg _429381_429381 ; 
   reg __429381_429381;
   reg _429382_429382 ; 
   reg __429382_429382;
   reg _429383_429383 ; 
   reg __429383_429383;
   reg _429384_429384 ; 
   reg __429384_429384;
   reg _429385_429385 ; 
   reg __429385_429385;
   reg _429386_429386 ; 
   reg __429386_429386;
   reg _429387_429387 ; 
   reg __429387_429387;
   reg _429388_429388 ; 
   reg __429388_429388;
   reg _429389_429389 ; 
   reg __429389_429389;
   reg _429390_429390 ; 
   reg __429390_429390;
   reg _429391_429391 ; 
   reg __429391_429391;
   reg _429392_429392 ; 
   reg __429392_429392;
   reg _429393_429393 ; 
   reg __429393_429393;
   reg _429394_429394 ; 
   reg __429394_429394;
   reg _429395_429395 ; 
   reg __429395_429395;
   reg _429396_429396 ; 
   reg __429396_429396;
   reg _429397_429397 ; 
   reg __429397_429397;
   reg _429398_429398 ; 
   reg __429398_429398;
   reg _429399_429399 ; 
   reg __429399_429399;
   reg _429400_429400 ; 
   reg __429400_429400;
   reg _429401_429401 ; 
   reg __429401_429401;
   reg _429402_429402 ; 
   reg __429402_429402;
   reg _429403_429403 ; 
   reg __429403_429403;
   reg _429404_429404 ; 
   reg __429404_429404;
   reg _429405_429405 ; 
   reg __429405_429405;
   reg _429406_429406 ; 
   reg __429406_429406;
   reg _429407_429407 ; 
   reg __429407_429407;
   reg _429408_429408 ; 
   reg __429408_429408;
   reg _429409_429409 ; 
   reg __429409_429409;
   reg _429410_429410 ; 
   reg __429410_429410;
   reg _429411_429411 ; 
   reg __429411_429411;
   reg _429412_429412 ; 
   reg __429412_429412;
   reg _429413_429413 ; 
   reg __429413_429413;
   reg _429414_429414 ; 
   reg __429414_429414;
   reg _429415_429415 ; 
   reg __429415_429415;
   reg _429416_429416 ; 
   reg __429416_429416;
   reg _429417_429417 ; 
   reg __429417_429417;
   reg _429418_429418 ; 
   reg __429418_429418;
   reg _429419_429419 ; 
   reg __429419_429419;
   reg _429420_429420 ; 
   reg __429420_429420;
   reg _429421_429421 ; 
   reg __429421_429421;
   reg _429422_429422 ; 
   reg __429422_429422;
   reg _429423_429423 ; 
   reg __429423_429423;
   reg _429424_429424 ; 
   reg __429424_429424;
   reg _429425_429425 ; 
   reg __429425_429425;
   reg _429426_429426 ; 
   reg __429426_429426;
   reg _429427_429427 ; 
   reg __429427_429427;
   reg _429428_429428 ; 
   reg __429428_429428;
   reg _429429_429429 ; 
   reg __429429_429429;
   reg _429430_429430 ; 
   reg __429430_429430;
   reg _429431_429431 ; 
   reg __429431_429431;
   reg _429432_429432 ; 
   reg __429432_429432;
   reg _429433_429433 ; 
   reg __429433_429433;
   reg _429434_429434 ; 
   reg __429434_429434;
   reg _429435_429435 ; 
   reg __429435_429435;
   reg _429436_429436 ; 
   reg __429436_429436;
   reg _429437_429437 ; 
   reg __429437_429437;
   reg _429438_429438 ; 
   reg __429438_429438;
   reg _429439_429439 ; 
   reg __429439_429439;
   reg _429440_429440 ; 
   reg __429440_429440;
   reg _429441_429441 ; 
   reg __429441_429441;
   reg _429442_429442 ; 
   reg __429442_429442;
   reg _429443_429443 ; 
   reg __429443_429443;
   reg _429444_429444 ; 
   reg __429444_429444;
   reg _429445_429445 ; 
   reg __429445_429445;
   reg _429446_429446 ; 
   reg __429446_429446;
   reg _429447_429447 ; 
   reg __429447_429447;
   reg _429448_429448 ; 
   reg __429448_429448;
   reg _429449_429449 ; 
   reg __429449_429449;
   reg _429450_429450 ; 
   reg __429450_429450;
   reg _429451_429451 ; 
   reg __429451_429451;
   reg _429452_429452 ; 
   reg __429452_429452;
   reg _429453_429453 ; 
   reg __429453_429453;
   reg _429454_429454 ; 
   reg __429454_429454;
   reg _429455_429455 ; 
   reg __429455_429455;
   reg _429456_429456 ; 
   reg __429456_429456;
   reg _429457_429457 ; 
   reg __429457_429457;
   reg _429458_429458 ; 
   reg __429458_429458;
   reg _429459_429459 ; 
   reg __429459_429459;
   reg _429460_429460 ; 
   reg __429460_429460;
   reg _429461_429461 ; 
   reg __429461_429461;
   reg _429462_429462 ; 
   reg __429462_429462;
   reg _429463_429463 ; 
   reg __429463_429463;
   reg _429464_429464 ; 
   reg __429464_429464;
   reg _429465_429465 ; 
   reg __429465_429465;
   reg _429466_429466 ; 
   reg __429466_429466;
   reg _429467_429467 ; 
   reg __429467_429467;
   reg _429468_429468 ; 
   reg __429468_429468;
   reg _429469_429469 ; 
   reg __429469_429469;
   reg _429470_429470 ; 
   reg __429470_429470;
   reg _429471_429471 ; 
   reg __429471_429471;
   reg _429472_429472 ; 
   reg __429472_429472;
   reg _429473_429473 ; 
   reg __429473_429473;
   reg _429474_429474 ; 
   reg __429474_429474;
   reg _429475_429475 ; 
   reg __429475_429475;
   reg _429476_429476 ; 
   reg __429476_429476;
   reg _429477_429477 ; 
   reg __429477_429477;
   reg _429478_429478 ; 
   reg __429478_429478;
   reg _429479_429479 ; 
   reg __429479_429479;
   reg _429480_429480 ; 
   reg __429480_429480;
   reg _429481_429481 ; 
   reg __429481_429481;
   reg _429482_429482 ; 
   reg __429482_429482;
   reg _429483_429483 ; 
   reg __429483_429483;
   reg _429484_429484 ; 
   reg __429484_429484;
   reg _429485_429485 ; 
   reg __429485_429485;
   reg _429486_429486 ; 
   reg __429486_429486;
   reg _429487_429487 ; 
   reg __429487_429487;
   reg _429488_429488 ; 
   reg __429488_429488;
   reg _429489_429489 ; 
   reg __429489_429489;
   reg _429490_429490 ; 
   reg __429490_429490;
   reg _429491_429491 ; 
   reg __429491_429491;
   reg _429492_429492 ; 
   reg __429492_429492;
   reg _429493_429493 ; 
   reg __429493_429493;
   reg _429494_429494 ; 
   reg __429494_429494;
   reg _429495_429495 ; 
   reg __429495_429495;
   reg _429496_429496 ; 
endmodule
