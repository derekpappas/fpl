`include "defines.v"

module t1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 298
  output [1 - 1:0] ar_sa0_s10;
  s1 s10(.ar_sa0_s10(ar_sa0_s10));
  `include "t1.logic.vh"
endmodule

