// Test type: Continuous assignment - wk1, sup0 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous436;
wire a;
assign (weak1, supply0) a=1'b1;
endmodule
