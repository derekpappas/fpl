//cp.vh