// Test type: Binary Numbers - No size specified lower case base
// Vparser rule name: Numbers
// Author: andreib
module binary_num;
wire a;
assign a='b1011;
endmodule
