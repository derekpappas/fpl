-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./chip_cslc_generated/code/vhdl/mecluster.vhd
-- FILE GENERATED ON : Wed Feb 18 21:22:52 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \mecluster\ is
begin
end entity;

architecture \mecluster_logic\ of \mecluster\ is

  component \me\ is
  end component;
begin
  \me0\ : \me\;
  \me1\ : \me\;
  \me2\ : \me\;
  \me3\ : \me\;
end architecture;

