//test type : specify_block_declaration 
//author : Dramba Doru-Gabriel
module recrem_specify_block0(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" ); endspecify
endmodule
module recrem_specify_block1(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , ); endspecify
endmodule
module recrem_specify_block2(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , ); endspecify
endmodule
module recrem_specify_block3(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , ); endspecify
endmodule
module recrem_specify_block4(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , ); endspecify
endmodule
module recrem_specify_block5(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , , ); endspecify
endmodule
module recrem_specify_block6(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block7(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block8(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block9(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier , ); endspecify
endmodule
module recrem_specify_block10(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block11(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block12(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier[3:3:3] ); endspecify
endmodule
module recrem_specify_block13(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier[3:3:3] , ); endspecify
endmodule
module recrem_specify_block14(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block15(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block16(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 ); endspecify
endmodule
module recrem_specify_block17(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , ); endspecify
endmodule
module recrem_specify_block18(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , , ); endspecify
endmodule
module recrem_specify_block19(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block20(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block21(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block22(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier , ); endspecify
endmodule
module recrem_specify_block23(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block24(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block25(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier[3:3:3] ); endspecify
endmodule
module recrem_specify_block26(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier[3:3:3] , ); endspecify
endmodule
module recrem_specify_block27(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block28(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block29(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 ); endspecify
endmodule
module recrem_specify_block30(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , ); endspecify
endmodule
module recrem_specify_block31(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , ); endspecify
endmodule
module recrem_specify_block32(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , , ); endspecify
endmodule
module recrem_specify_block33(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block34(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block35(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block36(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier , ); endspecify
endmodule
module recrem_specify_block37(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block38(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block39(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier[3:3:3] ); endspecify
endmodule
module recrem_specify_block40(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier[3:3:3] , ); endspecify
endmodule
module recrem_specify_block41(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block42(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block43(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 ); endspecify
endmodule
module recrem_specify_block44(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , ); endspecify
endmodule
module recrem_specify_block45(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , , ); endspecify
endmodule
module recrem_specify_block46(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block47(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block48(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block49(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier , ); endspecify
endmodule
module recrem_specify_block50(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block51(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block52(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] ); endspecify
endmodule
module recrem_specify_block53(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] , ); endspecify
endmodule
module recrem_specify_block54(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block55(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block56(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block57(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , ); endspecify
endmodule
module recrem_specify_block58(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , ); endspecify
endmodule
module recrem_specify_block59(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , ); endspecify
endmodule
module recrem_specify_block60(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , , ); endspecify
endmodule
module recrem_specify_block61(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block62(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block63(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block64(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier , ); endspecify
endmodule
module recrem_specify_block65(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block66(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block67(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier[3:3:3] ); endspecify
endmodule
module recrem_specify_block68(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier[3:3:3] , ); endspecify
endmodule
module recrem_specify_block69(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block70(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block71(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 ); endspecify
endmodule
module recrem_specify_block72(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , ); endspecify
endmodule
module recrem_specify_block73(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , , ); endspecify
endmodule
module recrem_specify_block74(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block75(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block76(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block77(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier , ); endspecify
endmodule
module recrem_specify_block78(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block79(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block80(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier[3:3:3] ); endspecify
endmodule
module recrem_specify_block81(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier[3:3:3] , ); endspecify
endmodule
module recrem_specify_block82(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block83(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block84(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 ); endspecify
endmodule
module recrem_specify_block85(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , ); endspecify
endmodule
module recrem_specify_block86(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , ); endspecify
endmodule
module recrem_specify_block87(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , , ); endspecify
endmodule
module recrem_specify_block88(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block89(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block90(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block91(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier , ); endspecify
endmodule
module recrem_specify_block92(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block93(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block94(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier[3:3:3] ); endspecify
endmodule
module recrem_specify_block95(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier[3:3:3] , ); endspecify
endmodule
module recrem_specify_block96(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block97(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block98(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 ); endspecify
endmodule
module recrem_specify_block99(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , ); endspecify
endmodule
module recrem_specify_block100(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , , ); endspecify
endmodule
module recrem_specify_block101(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block102(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block103(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block104(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier , ); endspecify
endmodule
module recrem_specify_block105(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block106(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
module recrem_specify_block107(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] ); endspecify
endmodule
module recrem_specify_block108(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] , ); endspecify
endmodule
module recrem_specify_block109(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier ); endspecify
endmodule
module recrem_specify_block110(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $recrem( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] ); endspecify
endmodule
