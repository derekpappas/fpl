//this is a celldefine legal test
`celldefine/*dsdsdsd*/
module mymodule;
endmodule

