//this is a celldefine legal test
`celldefine//
module mod;
wire x;
/**//***//**/`celldefine/***///sa
module mymodule;
endmodule
/****/`endcelldefine//haha
/*hihi*/endmodule
`endcelldefine
hihi
`endcelldefine
