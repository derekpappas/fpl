// Test type: Continuous assignment - pl1, wk0 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous421;
wire a;
assign (pull1, weak0) a=1'b1;
endmodule
