// Test type: loop statement - while
// Vparser rule name:
// Author: andreib
module loop_statement3;
reg a,b;
initial while (a==4'b0111) b=4'b1000;
endmodule
