//this is an illegal celldefine test
`celldefine
module x;
endmodule
hihihaha`endcelldefine
//
