//test type : block_item_declaration ::= integer list_of_block_variable_identifiers;
//vparser rule name : 
//author : Codrin
module test_0500;
  (* ints, realx = 0 *)
  integer a, b, c;
endmodule
