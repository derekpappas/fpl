// Test type: net_assignment - unary operator, 1 attribute instance
// Vparser rule name:
// Author: andreib
module netasign3;
wire a, b;
assign a=!(*b*)2;
endmodule
