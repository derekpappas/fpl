// Test type: Octal Numbers - space between base and octal value
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a=9'o 453;
endmodule
