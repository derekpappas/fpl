//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : reg.v
//FILE GENERATED ON : Wed Jul  9 20:26:20 2008

`include "defines.v"

module reg(dwdata,
           dwwr);
// Location of source csl unit: file name = generated/mitch.csl line number = 30
  input [31:0] dwdata;
  output dwwr;
  `include "reg.logic.v"
endmodule

