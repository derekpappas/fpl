//gate_instantiation = pullup ...;
//tests by Gabrield
module gate_instantiation_pullup0;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( output_terminal ) ;
endmodule
module gate_instantiation_pullup1;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup2;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup3;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup4;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup5;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup6;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup7;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup8;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup9;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup10;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup11;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup12;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup13;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup14;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup15;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup16;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup17;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup18;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup19;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup20;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup21;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup22;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup23;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup24;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup25;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup26;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup27;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup28;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup29;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup30;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup31;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup32;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup33;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup34;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup35;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup36;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup37;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup38;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup39;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup40;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup41;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup42;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup43;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup44;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup45;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup46;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup47;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup48;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup49;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup50;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup51;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup52;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup53;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup54;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup55;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup56;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup57;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup58;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup59;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup60;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup61;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup62;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup63;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup64;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup65;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup66;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup67;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup68;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup69;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup70;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup71;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup72;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup73;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup74;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup75;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup76;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup77;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup78;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup79;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup80;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup81;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup82;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup83;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup84;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup85;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup86;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup87;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup88;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup89;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup90;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup91;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup92;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup93;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup94;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup95;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup96;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup97;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup98;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup99;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup100;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup101;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup102;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup103;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup104;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup105;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup106;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup107;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup108;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup109;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup110;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup111;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup112;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup113;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup114;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup115;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup116;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup117;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup118;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup119;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup120;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup121;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup122;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup123;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup124;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup125;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup126;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup127;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup128;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup129;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup130;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup131;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup132;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup133;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup134;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup135;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup136;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup137;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup138;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup139;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup140;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup141;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup142;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup143;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup144;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup145;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup146;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup147;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup148;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup149;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup150;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup151;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup152;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup153;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup154;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup155;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup156;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup157;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup158;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup159;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup160;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup161;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup162;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup163;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup164;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup165;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup166;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup167;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup168;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup169;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup170;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup171;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup172;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup173;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup174;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup175;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup176;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup177;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup178;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup179;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup180;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup181;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup182;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup183;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup184;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup185;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup186;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup187;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup188;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup189;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup190;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup191;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup192;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup193;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup194;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup195;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup196;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup197;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup198;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup199;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup200;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup201;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup202;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup203;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup204;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup205;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup206;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup207;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup208;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup209;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup210;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup211;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup212;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup213;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup214;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup215;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup216;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup217;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup218;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup219;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup220;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup221;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup222;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup223;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup224;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup225;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup226;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup227;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup228;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup229;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup230;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup231;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup232;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup233;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup234;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup235;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup236;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup237;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup238;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup239;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup240;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup241;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup242;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup243;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup244;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup245;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup246;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup247;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup248;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup249;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup250;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup251;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup252;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup253;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup254;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup255;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup256;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup257;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup258;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup259;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup260;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup261;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup262;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup263;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup264;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup265;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup266;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup267;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup268;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup269;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup270;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup271;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup272;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup273;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup274;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup275;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup276;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup277;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup278;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup279;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , supply1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup280;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup281;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup282;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup283;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup284;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup285;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup286;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup287;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup288;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup289;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup290;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup291;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup292;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup293;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup294;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup295;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup296;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup297;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup298;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup299;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , strong1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup300;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup301;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup302;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup303;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup304;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup305;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup306;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup307;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup308;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup309;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup310;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup311;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup312;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup313;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup314;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup315;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup316;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup317;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup318;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup319;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , pull1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup320;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup321;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup322;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup323;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup324;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup325;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup326;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup327;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup328;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup329;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup330;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup331;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup332;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup333;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup334;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup335;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup336;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup337;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup338;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup339;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak0 , weak1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup340;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup341;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup342;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup343;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup344;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup345;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup346;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup347;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup348;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup349;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup350;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup351;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup352;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup353;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup354;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup355;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup356;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup357;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup358;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup359;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup360;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup361;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup362;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup363;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup364;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup365;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup366;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup367;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup368;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup369;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup370;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup371;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup372;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup373;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup374;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup375;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup376;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup377;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup378;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup379;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup380;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup381;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup382;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup383;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup384;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup385;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup386;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup387;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup388;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup389;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup390;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup391;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup392;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup393;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup394;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup395;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup396;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup397;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup398;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup399;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup400;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup401;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup402;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup403;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup404;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup405;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup406;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup407;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup408;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup409;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup410;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup411;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup412;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup413;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup414;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup415;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup416;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup417;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup418;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup419;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup420;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup421;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup422;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup423;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup424;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup425;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup426;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup427;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup428;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup429;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup430;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup431;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup432;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup433;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup434;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup435;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup436;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup437;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup438;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup439;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup440;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup441;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup442;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup443;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup444;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup445;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup446;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup447;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup448;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup449;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup450;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup451;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup452;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup453;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup454;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup455;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup456;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup457;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup458;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup459;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup460;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup461;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup462;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup463;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup464;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup465;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup466;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup467;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup468;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup469;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup470;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup471;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup472;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup473;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup474;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup475;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup476;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup477;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup478;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup479;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup480;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup481;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup482;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup483;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup484;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup485;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup486;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup487;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup488;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup489;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup490;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup491;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup492;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup493;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup494;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup495;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup496;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup497;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup498;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup499;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup500;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup501;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup502;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup503;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup504;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup505;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup506;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup507;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup508;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup509;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup510;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup511;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup512;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup513;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup514;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup515;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup516;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup517;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup518;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup519;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup520;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup521;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup522;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup523;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup524;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup525;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup526;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup527;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup528;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup529;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup530;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup531;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup532;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup533;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup534;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup535;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup536;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup537;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup538;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup539;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup540;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup541;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup542;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup543;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup544;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup545;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup546;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup547;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup548;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup549;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup550;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup551;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup552;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup553;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup554;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup555;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup556;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup557;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup558;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup559;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup560;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup561;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup562;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup563;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup564;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup565;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup566;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup567;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup568;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup569;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup570;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup571;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup572;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup573;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup574;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup575;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup576;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup577;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup578;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup579;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup580;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup581;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup582;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup583;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup584;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup585;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup586;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup587;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup588;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup589;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup590;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup591;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup592;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup593;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup594;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup595;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup596;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup597;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup598;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup599;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , supply0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup600;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup601;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup602;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup603;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup604;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup605;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup606;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup607;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup608;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup609;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup610;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup611;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup612;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup613;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup614;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup615;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup616;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup617;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup618;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup619;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , strong0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup620;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup621;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup622;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup623;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup624;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup625;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup626;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup627;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup628;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup629;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup630;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup631;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup632;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup633;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup634;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup635;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup636;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup637;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup638;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup639;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , pull0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup640;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup641;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup642;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup643;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup644;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup645;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup646;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup647;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup648;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup649;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup650;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup651;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup652;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup653;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup654;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup655;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup656;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup657;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup658;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup659;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 , weak0 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup660;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup661;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup662;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup663;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup664;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup665;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup666;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup667;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup668;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup669;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup670;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup671;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup672;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup673;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup674;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup675;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup676;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup677;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup678;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup679;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( supply1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup680;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup681;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup682;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup683;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup684;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup685;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup686;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup687;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup688;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup689;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup690;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup691;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup692;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup693;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup694;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup695;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup696;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup697;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup698;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup699;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( strong1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup700;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup701;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup702;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup703;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup704;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup705;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup706;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup707;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup708;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup709;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup710;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup711;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup712;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup713;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup714;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup715;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup716;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup717;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup718;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup719;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( pull1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup720;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pullup721;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup722;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup723;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup724;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup725;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup726;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup727;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup728;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup729;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup730;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) name1 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup731;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) name1 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup732;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) name1 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup733;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) name1 ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup734;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) name1 ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup735;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) name1 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup736;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) name1 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pullup737;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) name1 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pullup738;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pullup739;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pullup ( weak1 ) name1 ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
